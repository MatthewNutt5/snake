magic
tech scmos
timestamp 1745462530
<< m2contact >>
rect -2 -2 2 2
<< end >>
