../Synthesis/logic.vh