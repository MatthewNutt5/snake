../Synthesis/top.vh