//======================================
// Snake Game Logic Datapath - logic.v
//======================================
module logic (clka, clkb, restart, from_controller, direction_state, prng_done,
  random_num, to_controller, led_array_flat, request_rand);

/*
 *  This datapath module handles all of the game logic for Snake.
 *  On each game tick,
 *    1) Based on the direction the snake is currently moving, the head position
 *       is updated.
 *    2) After updating the head, the new head position is loaded onto a shift
 *       register holding the locations of each body piece.
 *    3) The new head position is checked for collisions with any body piece.
 *       If a collision is detected, then the game ends.
 *    4) The new head position is checked for a collision with the current apple
 *       location. If a collision is detected, then the snake grows one segment
 *       longer, and a new apple position must be generated by the PRNG module.
 *    5) After all updates are complete, the LED array representing the game
 *       board/display must be updated with each body piece and the apple.
 */

/*
 *  NOTE: To make development easier, we should probably try to keep things
 *        simple for now. It isn't ideal if the PRNG module returns an apple
 *        location that coincides with a current body location, but that would
 *        be another collision check, necessitate a repeat, etc.
 */



//========== Setup ==========

//---------- Input Ports ----------

/*
 *  Various single-wire inputs.
 *  - clka and clkb are provided by oscillator
 *  - restart could come from a button
 */
input wire clka, clkb, restart;

/*
 *  Signal array from controller FSM. Each index represents a different signal.
 *  - to_logic[LOGIC_TICK] tells the logic datapath when to intake a new
 *    direction input and update the game board.
 *  - to_logic[NO_UPDATE], when enabled during the tick, will blink the LED that
 *    represents the head position, instead of taking input and updating. Used
 *    after the game has ended.
 */
input wire [1:0] from_controller;
parameter LOGIC_TICK = 0, NO_UPDATE = 1;

/*
 *  Represents the direction the snake is moving.
 */
input wire [1:0] direction_state;
parameter UP_STATE = 0, DOWN_STATE = 1, LEFT_STATE = 2, RIGHT_STATE = 3;

/*
 *  Signal from PRNG module indicating when a new random number is ready.
 */
input wire prng_done;

/*
 *  6-bit random number generated by PRNG module.
 */
input wire [5:0] random_num;



//---------- Output Ports ----------

/*
 *  Signal array to controller FSM. Each index represents a different signal.
 */
output reg [1:0] to_controller;
parameter LOGIC_DONE = 0, GAME_END = 1;

/*
 *  Flattened version of a nested array denoting which LEDs should be lit.
 *  - led_array[r] is the r-th row, led_array[r][c] is the c-th column in the
 *    r-th row.
 *  - Indexes off the bottom-left corner of the display matrix.
 *  - Flattened version starts with 0-th row, then 1-st row, etc., unflattened
 *    by internal wire.
 */
output reg [63:0] led_array_flat;

/*
 *  Signal sent to PRNG datapath when a new random number is needed.
 */
output reg request_rand;



//---------- Internal Variables ----------

/*
 *  Unflattens output led_array_flat.
 *  NOTE: Is it necessary to unflatten led_array if we just end up having to 
 *  flatten it for output anyway?
 */
wire [7:0] led_array [7:0];
assign led_array[0] = led_array_flat[7:0];
assign led_array[1] = led_array_flat[15:8];
assign led_array[2] = led_array_flat[23:16];
assign led_array[3] = led_array_flat[31:24];
assign led_array[4] = led_array_flat[39:32];
assign led_array[5] = led_array_flat[47:40];
assign led_array[6] = led_array_flat[55:48];
assign led_array[7] = led_array_flat[63:56];


/*
 *  Various registers for holding the value of inputs at clka.
 */
reg restart_temp;
reg direction_state_temp;
reg [1:0] from_controller_temp;
reg prng_done_temp;
reg [5:0] random_num_temp;

/*
 *  Temp registers for holding the value of outputs at clka.
 */
reg [1:0] to_controller_temp;
reg request_rand_temp;

// May need counters here for iterating over multiple clock cycles
// Definitely put the shift register, next head location, apple location, and
// current snake length here

/*
*  64 6-bit registers. The n-th register keeps track of the position of the n-th
*  body part of the snake. snake_body[n][2:0] will be the x-position, and
*  snake_body[n][5:3] will be the y-position.
*/
reg [5:0] snake_body [63:0];

/*
*  Register to store the location of the next head, determined by the current
*  direction_state.
*/
reg [5:0] next_head;

/*
*  Register to store the location of the apple on the board. This is determined
*  by our PRNG module. 
*/
reg [5:0] apple_location;

/*
*  Register to keep track of the current snake length, for score keeping purposes
*  as well as boundary conditions.
*/
reg [5:0] snake_length;


/*
*  Logic to determine next_head based on direction_state. 
*  NOTE: Our direction FSM takes care of cases where we're moving up
*  and an up or down input is applied, so we don't need to worry about
*  those cases here. We do however, care about the grid boundaries.
*  Enter collision detection.
*/
always @(*) begin
  if (direction_state == UP_STATE)begin
    next_head[5:3] = snake_body[0][5:3] + 1'b1; 
  end else if (direction_state == DOWN_STATE) begin
    next_head[5:3] = snake_body[0][5:3] - 1'b1; 
  end else if (direction_state == RIGHT_STATE) begin
    next_head[2:0] = snake_body[0][2:0] + 1'b1; 
  end else if (direction_state == LEFT_STATE) begin
    next_head[2:0] = snake_body[0][2:0] - 1'b1; 
  end
end


//========== Code ==========

//---------- Sequential Logic ----------

/*
 *  Inputs should be evaluated/saved on clka to maintain timing discipline.
 *  Internal logic can also be updated in this section, but avoid updating
 *  any outputs until clkb; use temporary registers if necessary.
 */

always @(negedge clka) begin
  
  integer i = 0;
  integer j = 0;
  restart_temp = restart;
  direction_state_temp = direction_state;
  from_controller_temp = from_controller;

  if (restart) begin

    to_controller_temp = 2'b11;
    snake_body[0] = 100100; //"middle" of board for now
    for (i = 1; i < 64; i = i + 1)begin //reset all registers to 0
      snake_body[i] = 0;
    end
    for (j = 0; j < 64; j = j + 1)begin
      led_array_flat[j] = 0;
    end
    snake_length = 1; 
    led_array_flat[36] = 1; //turn on led at middle of board. could turn on at game_start instead

  end else begin
    for (i = 0; i < snake_length; i = i + 1)begin
      snake_body[i + 1] = snake_body[i];
      //turn on the led at (x_pos, y_pos) of i-th body piece
      //led_array[snake_body[i + 1][5:3]][snake_body[i + 1][2:0]] = 1;
      led_array_flat[(8*snake_body[i + 1][5:3]) + snake_body[i + 1][2:0]] = 1
    end
    snake_body[0] = next_head;
    led_array_flat[(8*snake_body[0][5:3]) + snake_body[0][2:0]] = 1;

  end

end



//---------- Output Logic ----------

/*
 *  Outputs should be updated on clkb to maintain timing discipline.
 */

always @(negedge clkb) begin

  if (restart_temp) begin
    led_array_flat <= 0;
  end

end



endmodule
