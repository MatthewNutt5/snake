../Synthesis/prng.vh