magic
tech scmos
magscale 1 2
timestamp 1744683001
<< nwell >>
rect -16 96 92 210
<< ntransistor >>
rect 14 12 18 52
rect 30 12 34 52
rect 46 12 50 52
rect 62 12 66 52
<< ptransistor >>
rect 14 108 18 188
rect 24 108 28 188
rect 52 108 56 188
rect 62 108 66 188
<< ndiffusion >>
rect 4 51 14 52
rect 12 13 14 51
rect 4 12 14 13
rect 18 42 30 52
rect 18 14 20 42
rect 28 14 30 42
rect 18 12 30 14
rect 34 51 46 52
rect 34 13 36 51
rect 44 13 46 51
rect 34 12 46 13
rect 50 24 52 52
rect 60 24 62 52
rect 50 12 62 24
rect 66 51 76 52
rect 66 13 68 51
rect 66 12 76 13
<< pdiffusion >>
rect 4 187 14 188
rect 12 109 14 187
rect 4 108 14 109
rect 18 108 24 188
rect 28 187 52 188
rect 28 109 31 187
rect 49 109 52 187
rect 28 108 52 109
rect 56 108 62 188
rect 66 187 76 188
rect 66 109 68 187
rect 66 108 76 109
<< ndcontact >>
rect 4 13 12 51
rect 20 14 28 42
rect 36 13 44 51
rect 52 24 60 52
rect 68 13 76 51
<< pdcontact >>
rect 4 109 12 187
rect 31 109 49 187
rect 68 109 76 187
<< psubstratepcontact >>
rect -4 -4 4 4
rect 28 -4 36 4
rect 60 -4 68 4
<< nsubstratencontact >>
rect -4 196 4 204
rect 28 196 36 204
rect 60 196 68 204
<< polysilicon >>
rect 14 188 18 192
rect 24 188 28 192
rect 52 188 56 192
rect 62 188 66 192
rect 14 98 18 108
rect 24 106 28 108
rect 52 106 56 108
rect 24 102 34 106
rect 8 94 18 98
rect 8 66 12 94
rect 30 86 34 102
rect 28 78 34 86
rect 14 52 18 62
rect 30 52 34 78
rect 50 102 56 106
rect 62 106 66 108
rect 62 102 74 106
rect 50 86 54 102
rect 50 78 52 86
rect 70 82 74 102
rect 50 62 54 78
rect 46 58 54 62
rect 70 60 74 74
rect 46 52 50 58
rect 62 56 74 60
rect 62 52 66 56
rect 14 8 18 12
rect 30 8 34 12
rect 46 8 50 12
rect 62 8 66 12
<< polycontact >>
rect 20 78 28 86
rect 12 62 20 70
rect 52 78 60 86
rect 68 74 76 82
<< metal1 >>
rect -4 204 84 206
rect 4 196 28 204
rect 36 196 60 204
rect 68 196 84 204
rect -4 194 84 196
rect 4 187 12 194
rect 4 108 12 109
rect 30 187 50 188
rect 30 109 31 187
rect 49 109 50 187
rect 30 108 50 109
rect 68 187 76 194
rect 68 108 76 109
rect 20 86 28 94
rect 36 74 42 108
rect 52 86 60 94
rect 4 72 12 74
rect 36 72 44 74
rect 4 70 20 72
rect 4 66 12 70
rect 36 66 60 72
rect 68 66 76 74
rect 6 52 42 56
rect 54 52 60 66
rect 4 51 44 52
rect 12 50 36 51
rect 4 12 12 13
rect 20 42 28 44
rect 20 6 28 14
rect 68 51 76 52
rect 44 13 68 18
rect 36 12 76 13
rect -4 4 84 6
rect 4 -4 28 4
rect 36 -4 60 4
rect 68 -4 84 4
rect -4 -6 84 -4
<< m1p >>
rect 20 86 28 94
rect 52 86 60 94
rect 4 66 12 74
rect 36 66 44 74
rect 68 66 76 74
<< labels >>
rlabel metal1 8 0 8 0 4 gnd
rlabel metal1 8 200 8 200 4 vdd
rlabel metal1 56 90 56 90 4 D
rlabel metal1 72 70 72 70 4 C
rlabel metal1 8 70 8 70 4 A
rlabel metal1 24 90 24 90 4 B
rlabel metal1 40 70 40 70 4 Y
<< end >>
