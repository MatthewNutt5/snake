magic
tech scmos
timestamp 1744683001
<< nwell >>
rect -8 48 104 105
<< ntransistor >>
rect 7 6 9 26
rect 15 6 17 16
rect 21 6 23 16
rect 29 6 31 16
rect 34 6 36 16
rect 43 6 45 16
rect 59 6 61 16
rect 64 6 66 16
rect 74 6 76 16
rect 79 6 81 16
rect 87 6 89 26
<< ptransistor >>
rect 7 54 9 94
rect 15 74 17 94
rect 21 74 23 94
rect 29 74 31 94
rect 35 74 37 94
rect 43 74 45 94
rect 59 74 61 94
rect 64 74 66 94
rect 74 84 76 94
rect 79 84 81 94
rect 87 54 89 94
<< ndiffusion >>
rect 2 25 7 26
rect 6 6 7 25
rect 9 25 14 26
rect 9 6 10 25
rect 82 25 87 26
rect 14 6 15 16
rect 17 6 21 16
rect 23 15 29 16
rect 23 6 24 15
rect 28 6 29 15
rect 31 6 34 16
rect 36 15 43 16
rect 36 6 37 15
rect 41 6 43 15
rect 45 15 50 16
rect 45 6 46 15
rect 54 15 59 16
rect 58 6 59 15
rect 61 6 64 16
rect 66 15 74 16
rect 66 6 68 15
rect 72 6 74 15
rect 76 6 79 16
rect 81 6 82 16
rect 86 6 87 25
rect 89 25 94 26
rect 89 6 90 25
<< pdiffusion >>
rect 2 93 7 94
rect 6 54 7 93
rect 9 55 10 94
rect 14 74 15 94
rect 17 74 21 94
rect 23 93 29 94
rect 23 74 24 93
rect 28 74 29 93
rect 31 74 35 94
rect 37 93 43 94
rect 37 74 38 93
rect 42 74 43 93
rect 45 93 50 94
rect 45 74 46 93
rect 54 93 59 94
rect 58 74 59 93
rect 61 74 64 94
rect 66 93 74 94
rect 66 74 68 93
rect 72 84 74 93
rect 76 84 79 94
rect 81 93 87 94
rect 81 84 82 93
rect 72 74 73 84
rect 9 54 14 55
rect 86 54 87 93
rect 89 93 94 94
rect 89 54 90 93
<< ndcontact >>
rect 2 6 6 25
rect 10 6 14 25
rect 24 6 28 15
rect 37 6 41 15
rect 46 6 50 15
rect 54 6 58 15
rect 68 6 72 15
rect 82 6 86 25
rect 90 6 94 25
<< pdcontact >>
rect 2 54 6 93
rect 10 55 14 94
rect 24 74 28 93
rect 38 74 42 93
rect 46 74 50 93
rect 54 74 58 93
rect 68 74 72 93
rect 82 54 86 93
rect 90 54 94 93
<< psubstratepcontact >>
rect -2 -2 2 2
rect 14 -2 18 2
rect 30 -2 34 2
rect 46 -2 50 2
rect 62 -2 66 2
rect 78 -2 82 2
<< nsubstratencontact >>
rect -2 98 2 102
rect 14 98 18 102
rect 30 98 34 102
rect 46 98 50 102
rect 62 98 66 102
rect 78 98 82 102
<< polysilicon >>
rect 7 94 9 96
rect 15 94 17 96
rect 21 94 23 96
rect 29 94 31 96
rect 35 94 37 96
rect 43 94 45 96
rect 59 94 61 96
rect 64 94 66 96
rect 74 94 76 96
rect 79 94 81 96
rect 87 94 89 96
rect 7 37 9 54
rect 15 46 17 74
rect 21 54 23 74
rect 29 71 31 74
rect 35 71 37 74
rect 25 50 31 52
rect 7 26 9 33
rect 15 16 17 42
rect 21 16 23 23
rect 29 16 31 50
rect 35 23 37 67
rect 43 61 45 74
rect 59 73 61 74
rect 50 71 61 73
rect 34 19 35 23
rect 34 16 36 19
rect 43 16 45 57
rect 64 67 66 74
rect 49 19 51 67
rect 63 65 66 67
rect 54 57 55 60
rect 54 24 56 57
rect 63 37 65 65
rect 74 61 76 84
rect 73 57 76 61
rect 79 53 81 84
rect 75 51 81 53
rect 64 33 65 37
rect 60 29 62 33
rect 74 31 76 47
rect 87 45 89 54
rect 85 41 89 45
rect 60 27 71 29
rect 74 27 75 31
rect 54 22 66 24
rect 49 17 61 19
rect 59 16 61 17
rect 64 16 66 22
rect 69 19 71 27
rect 69 17 76 19
rect 74 16 76 17
rect 79 16 81 31
rect 87 26 89 41
rect 7 4 9 6
rect 15 4 17 6
rect 21 4 23 6
rect 29 4 31 6
rect 34 4 36 6
rect 43 4 45 6
rect 59 4 61 6
rect 64 4 66 6
rect 74 4 76 6
rect 79 4 81 6
rect 87 4 89 6
<< polycontact >>
rect 27 67 31 71
rect 35 67 39 71
rect 21 50 25 54
rect 14 42 18 46
rect 6 33 10 37
rect 21 23 25 27
rect 41 57 45 61
rect 35 19 39 23
rect 49 67 53 71
rect 55 57 59 61
rect 69 57 73 61
rect 73 47 77 51
rect 60 33 64 37
rect 81 41 85 45
rect 75 27 79 31
<< metal1 >>
rect -2 102 98 103
rect 2 98 14 102
rect 18 98 30 102
rect 34 98 46 102
rect 50 98 62 102
rect 66 98 78 102
rect 82 98 98 102
rect -2 97 98 98
rect 10 94 14 97
rect 2 93 6 94
rect 24 93 28 94
rect 18 74 24 77
rect 38 93 42 97
rect 46 93 50 94
rect 54 93 58 97
rect 67 93 73 94
rect 67 74 68 93
rect 72 74 73 93
rect 82 93 86 97
rect 46 71 49 74
rect 39 68 49 71
rect 22 57 41 60
rect 54 57 55 61
rect 59 57 69 60
rect 54 54 57 57
rect 90 93 94 94
rect 6 50 21 52
rect 25 51 57 54
rect 90 51 94 54
rect 2 49 25 50
rect 77 48 94 51
rect 34 46 38 47
rect 18 43 38 46
rect 70 41 81 44
rect 10 34 26 37
rect 30 34 60 37
rect 10 33 14 34
rect 20 27 24 34
rect 90 31 94 48
rect 79 28 94 31
rect 2 25 6 26
rect 10 25 14 26
rect 90 25 94 28
rect 39 19 49 22
rect 46 16 49 19
rect 18 15 28 16
rect 18 13 24 15
rect 37 15 42 16
rect 41 6 42 15
rect 46 15 50 16
rect 54 15 58 16
rect 66 15 73 16
rect 66 13 68 15
rect 67 6 68 13
rect 72 6 73 15
rect 10 3 14 6
rect 37 3 42 6
rect 54 3 58 6
rect 82 3 86 6
rect -2 2 98 3
rect 2 -2 14 2
rect 18 -2 30 2
rect 34 -2 46 2
rect 50 -2 62 2
rect 66 -2 78 2
rect 82 -2 98 2
rect -2 -3 98 -2
<< m2contact >>
rect 18 70 22 74
rect 66 70 70 74
rect 26 63 30 67
rect 18 57 22 61
rect 2 50 6 54
rect 66 40 70 44
rect 26 34 30 38
rect 2 26 6 30
rect 18 16 22 20
rect 66 16 70 20
<< metal2 >>
rect 18 61 22 70
rect 18 54 22 57
rect 2 30 6 50
rect 18 50 21 54
rect 18 20 22 50
rect 26 38 30 63
rect 66 61 70 70
rect 66 57 69 61
rect 66 44 70 57
rect 66 20 70 40
<< m1p >>
rect 34 43 38 47
rect 90 43 94 47
rect 10 33 14 37
<< labels >>
rlabel metal1 12 35 12 35 4 CLK
rlabel metal1 4 100 4 100 4 vdd
rlabel metal1 36 45 36 45 4 D
rlabel metal1 4 0 4 0 4 gnd
rlabel metal1 92 45 92 45 4 Q
<< end >>
