//======================================
// Snake Game PRNG Datapath - prng.v
//======================================
module prng (clka, clkb, restart, request_rand, random_num);

/*
 *  This datapath module handles the random number generation for the game.
 *  It is based around a 6-bit LFSR.
 */

/*
 *  NOTE: To make development easier, we should probably try to keep things
 *        simple for now. We discussed different ways to seed the LFSR to make
 *        each game different from the last, but maybe this can wait until we
 *        get other parts working?
 */



//========== Setup ==========

//---------- Input Ports ----------

/*
 *  Various single-wire inputs.
 *  - clka and clkb are provided by oscillator
 *  - restart could come from a button
 */
input wire clka, clkb, restart;

/*
 *  Signal sent by the logic datapath when a new random number is needed.
 */
input wire request_rand;



//---------- Output Ports ----------

/*
 *  6-bit random number generated by PRNG module.
 */
output reg [5:0] random_num;



//---------- Internal Variables ----------

/*
 *  Hard-coded seed to initialize the LFSR with. In future versions, this may
 *  be replaced by some mechanism to randomize the seed.
 *  TODO: This is currently set to the initial position of the apple, since
 *        the logic datapath will always update the apple position with the
 *        current random number; besides the starting condition, this works
 *        since the datapath will only request a new random number when it's
 *        needed.
 */
parameter SEED = 6'b011101;

/*
 *  Temp registers to hold values of inputs at clka.
 */
reg restart_temp, request_rand_temp;





//========== Code ==========

//---------- Sequential Logic ----------

/*
 *  Inputs should be evaluated/saved on clka to maintain timing discipline.
 *  Internal logic can also be updated in this section, but avoid updating
 *  any outputs until clkb; use temporary registers if necessary.
 */

always @(negedge clka) begin

  restart_temp <= restart;
  request_rand_temp <= request_rand;

end



//---------- Output Logic ----------

/*
 *  Outputs should be updated on clkb to maintain timing discipline.
 */

always @(negedge clkb) begin

  if (restart_temp) 
    random_num <= SEED;
  else if (request_rand_temp) begin
    random_num <= (random_num >> 1) | ( (random_num[0] ^ random_num[1]) << 5);
  end

end



endmodule
