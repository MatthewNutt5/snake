//======================================
// Snake Game PRNG Datapath - prng.v
//======================================
module prng (clka, clkb, restart, request_rand, prng_done, random_num);

/*
 *  This datapath module handles the random number generation for the game.
 *  It is based around a 6-bit LFSR.
 */

/*
 *  NOTE: To make development easier, we should probably try to keep things
 *        simple for now. We discussed different ways to seed the LFSR to make
 *        each game different from the last, but maybe this can wait until we
 *        get other parts working?
 *  TODO: I forgot our LFSR research; is there a way to get a PRNG period longer
 *        than (2^6 - 1)?
 */



//========== Setup ==========

//---------- Input Ports ----------

/*
 *  Various single-wire inputs.
 *  - clka and clkb are provided by oscillator
 *  - restart could come from a button
 */
input wire clka, clkb, restart;

/*
 *  Signal sent by the logic datapath when a new random number is needed.
 */
input wire request_rand;



//---------- Output Ports ----------

/*
 *  Signal sent to the logic datapath when the next random number is ready.
 */
output reg prng_done;

/*
 *  6-bit random number generated by PRNG module.
 */
output reg [5:0] random_num;





//---------- Internal Variables ----------

/*
 *  Hard-coded seed to initialize the LFSR with. In future versions, this may
 *  be replaced by some mechanism to randomize the seed.
 */
parameter SEED = 6'b000000;

/*
 *  Temporary register for holding the next random number, in order to maintain
 *  timing discipline.
 */
reg [5:0] random_num_temp;





//========== Code ==========

//---------- Sequential Logic ----------

/*
 *  Inputs should be evaluated/saved on clka to maintain timing discipline.
 *  Internal logic can also be updated in this section, but avoid updating
 *  any outputs until clkb; use temporary registers if necessary.
 */

always @(negedge clka) begin

  if (restart) begin
    random_num_temp <= SEED;
  end

end



//---------- Output Logic ----------

/*
 *  Outputs should be updated on clkb to maintain timing discipline.
 */

always @(negedge clkb) begin

  random_num <= random_num_temp;

end



endmodule
