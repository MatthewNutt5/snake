magic
tech scmos
timestamp 1745960911
<< polysilicon >>
rect 1020 6540 5780 6800
rect 0 1020 260 5780
rect 1048 5569 5749 5772
rect 1048 1244 1204 5569
rect 1048 1241 1205 1244
rect 5636 1241 5749 5569
rect 1048 1047 5750 1241
rect 6540 1020 6800 5780
rect 1020 0 5780 260
<< metal1 >>
rect 0 6478 1015 6800
rect 1125 6494 1176 6531
rect 1420 6486 1480 6532
rect 1719 6492 1784 6531
rect 2016 6487 2081 6536
rect 2320 6496 2377 6530
rect 2625 6490 2682 6528
rect 2913 6484 2984 6531
rect 3215 6489 3285 6535
rect 3519 6485 3583 6535
rect 3817 6491 3882 6532
rect 4114 6495 4183 6536
rect 4420 6491 4481 6529
rect 4719 6485 4776 6529
rect 5327 6492 5376 6528
rect 5629 6493 5679 6526
rect 5785 6478 6800 6800
rect 0 5785 322 6478
rect 1619 5771 1632 5777
rect 2935 5771 2958 5807
rect 6478 5785 6800 6478
rect 1035 5757 1067 5771
rect 1088 5757 1095 5771
rect 1318 5758 1319 5771
rect 1333 5758 1917 5771
rect 1935 5759 2217 5771
rect 1935 5758 2154 5759
rect 2173 5758 2217 5759
rect 2236 5758 2519 5771
rect 2534 5758 3118 5771
rect 3134 5758 3417 5771
rect 3433 5758 3719 5771
rect 3733 5758 4018 5771
rect 4032 5758 4318 5771
rect 265 5619 310 5683
rect 1035 5532 1048 5757
rect 1204 5752 2838 5753
rect 267 5317 309 5384
rect 1035 5231 1048 5520
rect 266 5083 311 5085
rect 266 5018 314 5083
rect 266 5015 311 5018
rect 1035 4932 1048 5221
rect 272 4717 308 4782
rect 1035 4632 1048 4921
rect 1035 4280 1048 4620
rect 264 4111 306 4187
rect 265 4110 304 4111
rect 1035 3733 1048 4268
rect 1035 3432 1048 3721
rect 1035 3131 1048 3419
rect 271 2930 309 2979
rect 1035 2831 1048 3122
rect 279 2630 304 2666
rect 1035 2660 1048 2820
rect 1053 5569 2838 5752
rect 2935 5713 2958 5758
rect 4333 5758 4620 5771
rect 4633 5758 5220 5771
rect 5234 5758 5520 5771
rect 5534 5758 5771 5771
rect 2843 5693 2958 5713
rect 1053 2665 1204 5569
rect 2843 5543 2863 5693
rect 2963 5577 5749 5754
rect 5646 5484 5749 5577
rect 998 2647 1234 2660
rect 998 2640 1011 2647
rect 1030 2481 1043 2647
rect 1030 1934 1043 2468
rect 1030 1634 1043 1918
rect 1030 1331 1043 1619
rect 1030 1042 1043 1318
rect 1048 1244 1204 2641
rect 2335 1249 2358 1268
rect 1048 1241 1205 1244
rect 5636 1241 5749 5484
rect 5755 5532 5768 5758
rect 6494 5627 6532 5674
rect 5755 5231 5768 5517
rect 6496 5331 6523 5372
rect 5755 4931 5768 5221
rect 6480 5012 6540 5088
rect 5755 4900 5768 4919
rect 5755 4632 5768 4661
rect 5755 4331 5768 4617
rect 5755 4159 5768 4319
rect 5755 4140 5791 4159
rect 5755 3731 5768 4140
rect 5755 3430 5768 3719
rect 5755 3133 5768 3418
rect 5755 2834 5768 3121
rect 5755 2532 5768 2822
rect 5755 1932 5768 2519
rect 5755 1633 5768 1918
rect 5755 1332 5768 1621
rect 1048 1047 5750 1241
rect 5755 1042 5768 1321
rect 1035 1029 1317 1042
rect 1332 1029 1620 1042
rect 1632 1029 1919 1042
rect 1934 1029 2520 1042
rect 2533 1029 2820 1042
rect 2832 1029 3120 1042
rect 3133 1029 3420 1042
rect 3433 1029 3721 1042
rect 3734 1029 4322 1042
rect 4333 1029 4621 1042
rect 4632 1029 4921 1042
rect 4933 1029 5221 1042
rect 5233 1029 5521 1042
rect 5535 1040 5768 1042
rect 5535 1029 5758 1040
rect 0 322 322 1015
rect 6478 322 6800 1015
rect 0 0 1015 322
rect 5785 0 6800 322
<< m2contact >>
rect 1619 5777 1632 5784
rect 1067 5757 1088 5771
rect 1319 5758 1333 5771
rect 1917 5757 1935 5771
rect 2217 5758 2236 5771
rect 2519 5758 2534 5771
rect 3118 5758 3134 5771
rect 3417 5758 3433 5771
rect 3719 5758 3733 5771
rect 4018 5758 4032 5771
rect 1035 5520 1048 5532
rect 1035 5221 1048 5231
rect 1035 4921 1048 4932
rect 1035 4620 1048 4632
rect 1035 4268 1048 4280
rect 1035 3721 1048 3733
rect 1035 3419 1048 3432
rect 1035 3122 1048 3131
rect 1035 2820 1048 2831
rect 4318 5757 4333 5771
rect 4620 5758 4633 5771
rect 5220 5758 5234 5771
rect 5520 5758 5534 5771
rect 1234 2642 1254 2662
rect 1030 2468 1043 2481
rect 1030 1918 1043 1934
rect 1030 1619 1043 1634
rect 1030 1318 1043 1331
rect 5755 5517 5768 5532
rect 5755 5221 5768 5231
rect 5755 4919 5768 4931
rect 5755 4617 5768 4632
rect 5755 4319 5768 4331
rect 5755 3719 5768 3731
rect 5755 3418 5768 3430
rect 5755 3121 5768 3133
rect 5755 2822 5768 2834
rect 5755 2519 5768 2532
rect 5755 1918 5768 1932
rect 5755 1621 5768 1633
rect 5755 1321 5768 1332
rect 1024 1029 1035 1042
rect 1317 1029 1332 1042
rect 1620 1029 1632 1042
rect 1919 1029 1934 1042
rect 2520 1029 2533 1042
rect 2820 1029 2832 1042
rect 3120 1029 3133 1042
rect 3420 1029 3433 1042
rect 3721 1029 3734 1042
rect 4322 1029 4333 1042
rect 4621 1029 4632 1042
rect 4921 1029 4933 1042
rect 5221 1029 5233 1042
rect 5521 1029 5535 1042
rect 5758 1029 5768 1040
<< metal2 >>
rect 1023 5778 1029 5787
rect 1023 5774 1083 5778
rect 1071 5771 1083 5774
rect 1007 5757 1039 5766
rect 1030 5734 1039 5757
rect 1030 5725 1170 5734
rect 1019 5523 1035 5529
rect 1008 5457 1150 5466
rect 1141 5358 1150 5457
rect 1161 5378 1170 5725
rect 1257 5585 1266 5793
rect 1323 5771 1329 5781
rect 1344 5612 1353 5790
rect 1557 5784 1566 5790
rect 1644 5750 1653 5791
rect 1857 5786 1866 5790
rect 1923 5771 1929 5789
rect 1643 5748 1653 5750
rect 1643 5641 1652 5748
rect 1944 5741 1953 5790
rect 2157 5784 2166 5791
rect 2223 5771 2229 5781
rect 1943 5734 1953 5741
rect 1643 5632 1695 5641
rect 1344 5596 1352 5612
rect 1686 5608 1695 5632
rect 1943 5635 1952 5734
rect 2244 5650 2253 5791
rect 2457 5787 2466 5790
rect 2523 5771 2529 5781
rect 2544 5738 2553 5791
rect 3747 5790 3750 5792
rect 2757 5789 2766 5790
rect 3123 5771 3129 5781
rect 3144 5752 3153 5790
rect 3423 5771 3429 5782
rect 2398 5735 2553 5738
rect 2565 5749 3153 5752
rect 2244 5647 2314 5650
rect 1943 5626 2253 5635
rect 2244 5614 2253 5626
rect 2244 5611 2297 5614
rect 1686 5607 1953 5608
rect 1686 5604 2217 5607
rect 1344 5593 2009 5596
rect 1257 5582 1785 5585
rect 1782 5569 1785 5582
rect 2006 5568 2009 5593
rect 2214 5572 2217 5604
rect 2294 5572 2297 5611
rect 2311 5589 2314 5647
rect 2311 5586 2385 5589
rect 2382 5572 2385 5586
rect 2398 5569 2401 5735
rect 2565 5729 2568 5749
rect 3444 5742 3453 5790
rect 3723 5771 3729 5781
rect 2478 5726 2568 5729
rect 2583 5739 3453 5742
rect 2478 5571 2481 5726
rect 2583 5718 2586 5739
rect 3744 5733 3753 5790
rect 4023 5771 4029 5782
rect 2494 5715 2586 5718
rect 2597 5730 3753 5733
rect 2494 5568 2497 5715
rect 2597 5705 2600 5730
rect 4044 5717 4053 5790
rect 4323 5771 4329 5782
rect 2534 5702 2600 5705
rect 2613 5714 4053 5717
rect 2534 5568 2537 5702
rect 2613 5687 2616 5714
rect 4344 5707 4353 5790
rect 4623 5771 4629 5782
rect 2582 5684 2616 5687
rect 2678 5704 4353 5707
rect 2582 5567 2585 5684
rect 2678 5571 2681 5704
rect 4644 5698 4653 5790
rect 5223 5771 5229 5781
rect 2830 5695 4653 5698
rect 2830 5570 2833 5695
rect 5244 5689 5253 5790
rect 5523 5771 5529 5783
rect 5544 5736 5553 5790
rect 2926 5686 5253 5689
rect 2926 5573 2929 5686
rect 5244 5685 5253 5686
rect 5454 5733 5553 5736
rect 5454 5573 5457 5733
rect 5673 5544 5790 5553
rect 5673 5457 5682 5544
rect 5768 5523 5781 5529
rect 5643 5448 5682 5457
rect 1161 5369 1184 5378
rect 1141 5349 1184 5358
rect 5652 5360 5740 5369
rect 1153 5324 1182 5333
rect 1019 5223 1035 5229
rect 1153 5166 1162 5324
rect 1008 5157 1162 5166
rect 1173 5287 1190 5296
rect 1173 5132 1182 5287
rect 5731 5253 5740 5360
rect 5652 5246 5716 5253
rect 5641 5244 5716 5246
rect 5731 5244 5790 5253
rect 1126 5123 1182 5132
rect 1019 4923 1035 4929
rect 1126 4866 1135 5123
rect 1007 4857 1135 4866
rect 1178 5053 1186 5066
rect 1019 4623 1035 4629
rect 1019 4271 1035 4277
rect 1178 4043 1187 5053
rect 5707 4953 5716 5244
rect 5768 5223 5782 5229
rect 5707 4944 5790 4953
rect 5768 4923 5782 4929
rect 5768 4623 5781 4629
rect 5768 4323 5781 4329
rect 1007 4034 1187 4043
rect 1019 3723 1035 3729
rect 5768 3723 5781 3729
rect 1019 3423 1035 3429
rect 1019 3123 1035 3129
rect 1183 3066 1192 3471
rect 5768 3423 5781 3429
rect 5768 3123 5782 3129
rect 1006 3057 1192 3066
rect 1019 2823 1035 2829
rect 5768 2823 5781 2829
rect 5768 2522 5782 2529
rect 1019 2471 1030 2477
rect 1019 1923 1030 1929
rect 5768 1923 5782 1929
rect 1019 1623 1030 1629
rect 5768 1623 5782 1629
rect 1019 1323 1030 1329
rect 5768 1323 5784 1329
rect 1013 1029 1024 1035
rect 5768 1030 5779 1036
rect 5773 1029 5779 1030
rect 1013 1023 1019 1029
rect 1027 1019 1033 1029
rect 1323 1019 1329 1029
rect 1623 1019 1629 1029
rect 1923 1019 1929 1029
rect 2523 1019 2529 1029
rect 2823 1019 2829 1029
rect 3123 1019 3129 1029
rect 3423 1019 3429 1029
rect 3723 1019 3729 1029
rect 4323 1019 4329 1029
rect 4623 1019 4629 1029
rect 4923 1019 4929 1029
rect 5223 1019 5229 1029
rect 5523 1019 5529 1029
rect 5773 1023 5787 1029
rect 1023 1013 1033 1019
<< m3contact >>
rect 5638 5448 5643 5457
rect 1184 5367 1198 5380
rect 1184 5344 1201 5359
rect 5638 5356 5652 5371
rect 1182 5320 1199 5335
rect 1190 5285 1201 5297
rect 5641 5246 5652 5256
rect 1186 5053 1200 5067
rect 1183 3471 1202 3488
<< metal3 >>
rect 5637 5457 5644 5458
rect 5637 5448 5638 5457
rect 5643 5448 5644 5457
rect 5637 5447 5644 5448
rect 1183 5380 1199 5381
rect 1183 5367 1184 5380
rect 1198 5367 1199 5380
rect 1183 5366 1199 5367
rect 5637 5371 5653 5372
rect 1183 5359 1202 5360
rect 1183 5344 1184 5359
rect 1201 5344 1202 5359
rect 5637 5356 5638 5371
rect 5652 5356 5653 5371
rect 5637 5355 5653 5356
rect 1183 5343 1202 5344
rect 1181 5335 1200 5336
rect 1181 5320 1182 5335
rect 1199 5320 1200 5335
rect 1181 5319 1200 5320
rect 1189 5297 1202 5298
rect 1189 5285 1190 5297
rect 1201 5285 1202 5297
rect 1189 5284 1202 5285
rect 5640 5256 5653 5257
rect 5640 5246 5641 5256
rect 5652 5246 5653 5256
rect 5640 5245 5653 5246
rect 1185 5067 1201 5068
rect 1185 5053 1186 5067
rect 1200 5053 1201 5067
rect 1185 5052 1201 5053
rect 1182 3488 1203 3489
rect 1182 3471 1183 3488
rect 1202 3471 1203 3488
rect 1182 3470 1203 3471
use PadFrame64  PadFrame64_0
timestamp 1745621596
transform 1 0 2500 0 1 2400
box -2500 -2400 4300 4400
use top  top_0
timestamp 1745462530
transform 1 0 1196 0 1 1236
box 0 13 4448 4340
<< labels >>
rlabel metal1 290 2648 290 2648 1 GND!
rlabel metal1 284 4147 284 4147 1 p_in_restart
rlabel metal1 288 2955 288 2955 1 p_in_clkb
rlabel metal1 285 5652 286 5652 1 p_in_direction2
rlabel metal1 286 5349 286 5349 1 p_in_direction3
rlabel metal1 286 5051 286 5051 1 p_in_direction1
rlabel metal1 289 4750 289 4750 1 p_in_direction0
rlabel metal1 1149 6513 1149 6513 1 p_in_clka
rlabel metal1 1448 6509 1448 6509 1 p_out_row_cathode7
rlabel metal1 1749 6512 1749 6512 1 p_out_row_cathode6
rlabel metal1 2045 6512 2045 6512 1 p_out_row_cathode3
rlabel metal1 2651 6510 2651 6510 1 p_out_row_cathode1
rlabel metal1 2347 6515 2347 6515 1 p_out_row_cathode5
rlabel metal1 3250 6514 3250 6514 1 p_out_row_cathode2
rlabel metal1 3549 6511 3549 6511 1 p_out_row_cathode4
rlabel metal1 3847 6512 3847 6512 1 p_out_row_cathode0
rlabel metal1 2948 6508 2948 6508 1 Vdd!
rlabel metal1 4147 6515 4147 6515 1 p_out_column_anode7
rlabel metal1 4450 6511 4450 6511 1 p_out_column_anode6
rlabel metal1 4746 6509 4746 6509 1 p_out_column_anode1
rlabel metal1 5351 6512 5351 6512 1 p_out_column_anode0
rlabel metal1 5653 6511 5653 6511 1 p_out_column_anode5
rlabel metal1 6512 5651 6512 5651 1 p_out_column_anode3
rlabel metal1 6509 5352 6509 5352 1 p_out_column_anode2
rlabel metal1 6480 5012 6540 5088 1 p_out_column_anode4
<< end >>
