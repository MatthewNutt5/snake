magic
tech scmos
timestamp 1745462530
<< metal1 >>
rect 1714 4334 4445 4336
rect 1706 4333 4445 4334
rect 1706 4331 1717 4333
rect 14 4307 4434 4327
rect 38 4283 4410 4303
rect 14 4267 4434 4273
rect 4442 4256 4445 4333
rect 4370 4253 4445 4256
rect 138 4216 141 4225
rect 212 4223 229 4226
rect 602 4216 605 4225
rect 66 4213 92 4216
rect 114 4213 132 4216
rect 138 4213 173 4216
rect 268 4213 293 4216
rect 324 4213 341 4216
rect 380 4213 405 4216
rect 436 4213 453 4216
rect 492 4213 517 4216
rect 548 4213 565 4216
rect 572 4213 581 4216
rect 602 4213 613 4216
rect 620 4213 629 4216
rect 756 4213 773 4216
rect 852 4213 877 4216
rect 948 4213 973 4216
rect 1044 4213 1069 4216
rect 1140 4213 1165 4216
rect 1332 4213 1357 4216
rect 1428 4213 1445 4216
rect 1580 4213 1589 4216
rect 1786 4213 1804 4216
rect 1818 4213 1836 4216
rect 1938 4213 1949 4216
rect 1994 4213 2004 4216
rect 2060 4213 2085 4216
rect 2236 4213 2261 4216
rect 2372 4213 2397 4216
rect 2468 4213 2493 4216
rect 2586 4213 2596 4216
rect 2748 4213 2757 4216
rect 2906 4213 2917 4216
rect 108 4203 117 4206
rect 138 4203 148 4206
rect 562 4205 565 4213
rect 1946 4206 1949 4213
rect 2914 4206 2917 4213
rect 2986 4213 2997 4216
rect 3468 4213 3477 4216
rect 3484 4213 3493 4216
rect 3660 4213 3685 4216
rect 3812 4213 3821 4216
rect 3858 4213 3868 4216
rect 4010 4213 4020 4216
rect 4034 4213 4052 4216
rect 4074 4213 4084 4216
rect 4098 4213 4109 4216
rect 4156 4213 4165 4216
rect 636 4203 668 4206
rect 682 4203 692 4206
rect 1490 4203 1500 4206
rect 1946 4203 1956 4206
rect 1980 4203 1996 4206
rect 2572 4203 2588 4206
rect 2628 4203 2644 4206
rect 2914 4203 2924 4206
rect 2948 4203 2964 4206
rect 2986 4205 2989 4213
rect 3474 4205 3477 4213
rect 3818 4205 3821 4213
rect 4106 4206 4109 4213
rect 4106 4203 4116 4206
rect 38 4167 4410 4173
rect 66 4133 84 4136
rect 90 4133 100 4136
rect 154 4133 164 4136
rect 170 4133 180 4136
rect 204 4133 221 4136
rect 66 4103 69 4133
rect 90 4125 93 4133
rect 586 4127 589 4134
rect 98 4123 108 4126
rect 188 4123 197 4126
rect 260 4123 285 4126
rect 322 4123 332 4126
rect 338 4123 348 4126
rect 388 4123 413 4126
rect 450 4123 460 4126
rect 524 4123 549 4126
rect 580 4124 589 4127
rect 596 4123 605 4126
rect 618 4125 621 4146
rect 682 4133 700 4136
rect 746 4133 756 4136
rect 876 4133 884 4136
rect 898 4126 901 4134
rect 962 4133 972 4136
rect 1018 4133 1036 4136
rect 1050 4126 1053 4145
rect 3978 4143 3988 4146
rect 1394 4133 1412 4136
rect 1418 4133 1428 4136
rect 1450 4126 1453 4134
rect 1522 4133 1532 4136
rect 1572 4133 1581 4136
rect 1706 4126 1709 4135
rect 2226 4133 2236 4136
rect 642 4123 652 4126
rect 778 4123 796 4126
rect 802 4123 820 4126
rect 826 4123 844 4126
rect 892 4123 901 4126
rect 994 4123 1012 4126
rect 1018 4123 1053 4126
rect 1138 4123 1156 4126
rect 1162 4123 1180 4126
rect 1212 4123 1221 4126
rect 1420 4123 1429 4126
rect 1450 4123 1461 4126
rect 1644 4123 1669 4126
rect 1700 4123 1709 4126
rect 1772 4123 1797 4126
rect 1866 4123 1876 4126
rect 1956 4123 1981 4126
rect 2012 4123 2021 4126
rect 2148 4123 2157 4126
rect 2164 4123 2173 4126
rect 2210 4123 2220 4126
rect 2322 4123 2332 4126
rect 2442 4123 2452 4126
rect 2458 4123 2476 4126
rect 2522 4123 2532 4126
rect 2580 4123 2605 4126
rect 2682 4123 2692 4126
rect 2698 4123 2715 4126
rect 2732 4123 2741 4126
rect 2778 4123 2788 4126
rect 2932 4123 2957 4126
rect 2988 4123 2997 4126
rect 3050 4123 3060 4126
rect 3226 4123 3236 4126
rect 3266 4123 3269 4134
rect 3282 4133 3292 4136
rect 3418 4133 3436 4136
rect 3548 4133 3557 4136
rect 3578 4133 3588 4136
rect 3932 4133 3948 4136
rect 3972 4133 3989 4136
rect 3996 4133 4005 4136
rect 4100 4133 4109 4136
rect 4140 4133 4149 4136
rect 4156 4133 4173 4136
rect 4204 4133 4213 4136
rect 4244 4133 4253 4136
rect 4260 4133 4269 4136
rect 3282 4123 3300 4126
rect 3306 4123 3316 4126
rect 3372 4123 3381 4126
rect 3418 4123 3428 4126
rect 3562 4123 3572 4126
rect 3578 4123 3596 4126
rect 3626 4123 3636 4126
rect 3746 4123 3756 4126
rect 3890 4123 3900 4126
rect 3946 4123 3956 4126
rect 4036 4123 4045 4126
rect 4170 4123 4188 4126
rect 4210 4123 4228 4126
rect 4372 4123 4381 4126
rect 602 4116 605 4123
rect 602 4113 612 4116
rect 716 4113 725 4116
rect 802 4115 805 4123
rect 994 4115 997 4123
rect 1020 4113 1029 4116
rect 1076 4113 1085 4116
rect 122 4103 140 4106
rect 1074 4103 1092 4106
rect 3418 4103 3421 4123
rect 3972 4113 3981 4116
rect 14 4067 4434 4073
rect 66 4033 100 4036
rect 210 4033 236 4036
rect 698 4033 708 4036
rect 1074 4033 1092 4036
rect 1106 4026 1109 4036
rect 292 4023 301 4026
rect 308 4023 317 4026
rect 364 4023 373 4026
rect 530 4016 533 4025
rect 676 4023 685 4026
rect 874 4016 877 4026
rect 1076 4023 1085 4026
rect 1100 4023 1109 4026
rect 3034 4016 3037 4036
rect 3980 4023 3989 4026
rect 4188 4023 4197 4026
rect 114 4013 124 4016
rect 202 4006 205 4014
rect 266 4013 276 4016
rect 148 4003 180 4006
rect 202 4003 213 4006
rect 250 4003 268 4006
rect 292 4003 301 4006
rect 314 4003 317 4014
rect 338 4013 348 4016
rect 418 4013 436 4016
rect 450 4013 468 4016
rect 530 4013 548 4016
rect 586 4013 604 4016
rect 644 4013 653 4016
rect 860 4013 892 4016
rect 1042 4013 1068 4016
rect 1154 4013 1172 4016
rect 1282 4013 1300 4016
rect 1322 4013 1356 4016
rect 1370 4013 1413 4016
rect 1524 4013 1549 4016
rect 1644 4013 1685 4016
rect 1730 4013 1748 4016
rect 1754 4013 1764 4016
rect 1780 4013 1805 4016
rect 1852 4013 1877 4016
rect 2004 4013 2021 4016
rect 2060 4013 2077 4016
rect 2194 4013 2237 4016
rect 2346 4013 2364 4016
rect 610 4003 636 4006
rect 650 4005 653 4013
rect 1730 4006 1733 4013
rect 2194 4006 2197 4013
rect 834 4003 852 4006
rect 916 4003 941 4006
rect 1178 4003 1204 4006
rect 1234 4003 1252 4006
rect 1282 4003 1292 4006
rect 1306 4003 1348 4006
rect 1362 4003 1372 4006
rect 1650 4003 1684 4006
rect 1716 4003 1733 4006
rect 2066 4003 2092 4006
rect 2122 4003 2164 4006
rect 2180 4003 2197 4006
rect 2234 4003 2237 4013
rect 2338 4003 2356 4006
rect 2410 4005 2413 4016
rect 2540 4013 2549 4016
rect 2554 4013 2572 4016
rect 2626 4013 2644 4016
rect 2706 4013 2724 4016
rect 2892 4013 2917 4016
rect 3034 4013 3044 4016
rect 3148 4013 3173 4016
rect 3204 4013 3213 4016
rect 3268 4013 3293 4016
rect 3484 4013 3501 4016
rect 3748 4013 3757 4016
rect 3794 4013 3812 4016
rect 3930 4013 3964 4016
rect 4002 4013 4020 4016
rect 4076 4013 4101 4016
rect 4116 4013 4125 4016
rect 2626 4006 2629 4013
rect 2620 4003 2629 4006
rect 2658 4003 2676 4006
rect 3026 4003 3052 4006
rect 3210 4003 3213 4013
rect 3450 4003 3460 4006
rect 3980 4003 4005 4006
rect 4036 4003 4052 4006
rect 4090 4003 4108 4006
rect 4138 4003 4163 4006
rect 4188 4003 4197 4006
rect 4228 4003 4237 4006
rect 4244 4003 4269 4006
rect 130 3993 140 3996
rect 210 3983 213 4003
rect 474 3993 484 3996
rect 1106 3993 1132 3996
rect 1282 3993 1285 4003
rect 4082 3993 4099 3996
rect 38 3967 4410 3973
rect 532 3943 548 3946
rect 762 3943 772 3946
rect 108 3933 124 3936
rect 138 3933 156 3936
rect 290 3933 308 3936
rect 498 3926 501 3936
rect 556 3933 581 3936
rect 612 3933 629 3936
rect 730 3933 756 3936
rect 1026 3933 1044 3936
rect 1482 3926 1485 3935
rect 1602 3926 1605 3935
rect 1698 3933 1708 3936
rect 1762 3933 1780 3936
rect 146 3923 164 3926
rect 228 3923 245 3926
rect 284 3923 301 3926
rect 306 3923 316 3926
rect 428 3923 469 3926
rect 476 3923 501 3926
rect 532 3923 549 3926
rect 570 3923 596 3926
rect 964 3923 989 3926
rect 1026 3923 1052 3926
rect 1058 3923 1076 3926
rect 1132 3923 1157 3926
rect 1188 3923 1197 3926
rect 1244 3923 1269 3926
rect 1300 3923 1317 3926
rect 1412 3923 1437 3926
rect 1468 3923 1485 3926
rect 1492 3923 1501 3926
rect 1540 3923 1565 3926
rect 1596 3923 1605 3926
rect 1682 3923 1692 3926
rect 1746 3923 1756 3926
rect 1818 3923 1828 3926
rect 1834 3923 1852 3926
rect 172 3913 189 3916
rect 1058 3915 1061 3923
rect 1914 3903 1917 3956
rect 3210 3936 3213 3956
rect 2204 3933 2212 3936
rect 2004 3923 2013 3926
rect 2060 3923 2069 3926
rect 2106 3923 2116 3926
rect 2178 3923 2188 3926
rect 2210 3923 2220 3926
rect 2250 3923 2253 3935
rect 2314 3933 2325 3936
rect 3060 3933 3077 3936
rect 3138 3933 3156 3936
rect 3210 3933 3228 3936
rect 3242 3933 3252 3936
rect 3274 3933 3292 3936
rect 3354 3933 3364 3936
rect 3418 3933 3444 3936
rect 3538 3933 3556 3936
rect 3572 3933 3589 3936
rect 2266 3923 2276 3926
rect 2298 3923 2308 3926
rect 2314 3915 2317 3933
rect 3658 3926 3661 3946
rect 3972 3933 3989 3936
rect 4020 3933 4036 3936
rect 4066 3933 4084 3936
rect 4090 3933 4108 3936
rect 4114 3933 4140 3936
rect 4188 3933 4197 3936
rect 4228 3933 4237 3936
rect 4244 3933 4269 3936
rect 2356 3923 2365 3926
rect 2418 3923 2428 3926
rect 2540 3923 2549 3926
rect 2604 3923 2629 3926
rect 2666 3923 2684 3926
rect 2714 3923 2724 3926
rect 2730 3923 2739 3926
rect 2802 3923 2819 3926
rect 2874 3923 2884 3926
rect 2898 3923 2907 3926
rect 3122 3923 3132 3926
rect 3194 3923 3204 3926
rect 3226 3923 3236 3926
rect 3282 3923 3300 3926
rect 3330 3923 3340 3926
rect 3402 3923 3412 3926
rect 3418 3923 3452 3926
rect 3586 3923 3604 3926
rect 3634 3923 3644 3926
rect 3658 3923 3676 3926
rect 3682 3923 3692 3926
rect 3722 3923 3740 3926
rect 4060 3923 4077 3926
rect 2666 3883 2669 3923
rect 2748 3913 2757 3916
rect 4020 3913 4037 3916
rect 4188 3913 4197 3916
rect 14 3867 4434 3873
rect 92 3813 101 3816
rect 132 3813 149 3816
rect 154 3806 157 3814
rect 180 3813 197 3816
rect 340 3813 365 3816
rect 466 3813 492 3816
rect 604 3813 637 3816
rect 732 3813 765 3816
rect 804 3813 853 3816
rect 892 3813 917 3816
rect 948 3813 965 3816
rect 1020 3813 1045 3816
rect 1076 3813 1109 3816
rect 1116 3813 1133 3816
rect 1188 3813 1205 3816
rect 1220 3813 1229 3816
rect 1244 3813 1277 3816
rect 1284 3813 1293 3816
rect 1308 3813 1333 3816
rect 1372 3813 1397 3816
rect 1484 3813 1509 3816
rect 1572 3813 1589 3816
rect 1626 3813 1636 3816
rect 1698 3813 1708 3816
rect 138 3803 157 3806
rect 178 3803 196 3806
rect 220 3803 245 3806
rect 474 3803 484 3806
rect 762 3805 765 3813
rect 1106 3805 1109 3813
rect 1122 3803 1132 3806
rect 1162 3803 1180 3806
rect 1274 3805 1277 3813
rect 1714 3806 1717 3836
rect 2706 3833 2724 3836
rect 2058 3823 2069 3826
rect 2186 3823 2196 3826
rect 2220 3823 2229 3826
rect 2292 3823 2301 3826
rect 2306 3823 2316 3826
rect 2340 3823 2349 3826
rect 2380 3823 2397 3826
rect 1770 3813 1780 3816
rect 1932 3813 1949 3816
rect 1989 3813 2005 3816
rect 2052 3813 2061 3816
rect 1546 3803 1564 3806
rect 1578 3803 1588 3806
rect 1642 3803 1660 3806
rect 1714 3803 1732 3806
rect 1804 3803 1821 3806
rect 1852 3803 1861 3806
rect 2002 3805 2005 3813
rect 2018 3803 2028 3806
rect 2066 3805 2069 3823
rect 2076 3813 2108 3816
rect 2234 3813 2244 3816
rect 2298 3813 2301 3823
rect 2346 3816 2349 3823
rect 2306 3813 2324 3816
rect 2346 3813 2364 3816
rect 2474 3813 2483 3816
rect 2306 3806 2309 3813
rect 2506 3806 2509 3826
rect 2524 3823 2533 3826
rect 2604 3823 2613 3826
rect 2692 3823 2701 3826
rect 2708 3823 2717 3826
rect 3460 3823 3469 3826
rect 3572 3823 3581 3826
rect 2516 3813 2525 3816
rect 2530 3813 2540 3816
rect 2572 3813 2589 3816
rect 2596 3813 2613 3816
rect 2658 3813 2674 3816
rect 2698 3813 2716 3816
rect 2874 3813 2891 3816
rect 3044 3813 3069 3816
rect 3154 3813 3164 3816
rect 3276 3813 3301 3816
rect 3338 3813 3356 3816
rect 3386 3813 3396 3816
rect 3402 3813 3428 3816
rect 3620 3813 3629 3816
rect 3666 3813 3684 3816
rect 3690 3813 3700 3816
rect 3748 3813 3757 3816
rect 3860 3813 3869 3816
rect 3956 3813 3965 3816
rect 4132 3813 4157 3816
rect 4210 3813 4220 3816
rect 4250 3813 4260 3816
rect 2698 3806 2701 3813
rect 2124 3803 2133 3806
rect 2292 3803 2309 3806
rect 2434 3803 2444 3806
rect 2466 3803 2476 3806
rect 2522 3803 2548 3806
rect 2570 3803 2588 3806
rect 2644 3803 2661 3806
rect 2692 3803 2701 3806
rect 3210 3803 3219 3806
rect 3500 3803 3509 3806
rect 3514 3803 3532 3806
rect 3548 3803 3565 3806
rect 3922 3803 3948 3806
rect 4018 3803 4028 3806
rect 4066 3803 4076 3806
rect 4114 3803 4124 3806
rect 4130 3803 4155 3806
rect 180 3793 189 3796
rect 3178 3793 3188 3796
rect 4066 3783 4069 3803
rect 38 3767 4410 3773
rect 1858 3743 1884 3746
rect 2042 3736 2045 3746
rect 2346 3736 2349 3756
rect 2498 3743 2508 3746
rect 2698 3743 2707 3746
rect 650 3733 668 3736
rect 682 3726 685 3735
rect 1306 3733 1332 3736
rect 1458 3733 1484 3736
rect 1490 3733 1500 3736
rect 1690 3733 1708 3736
rect 1730 3733 1740 3736
rect 1754 3733 1772 3736
rect 1796 3733 1813 3736
rect 580 3723 605 3726
rect 676 3723 685 3726
rect 692 3723 701 3726
rect 764 3723 789 3726
rect 820 3723 837 3726
rect 876 3723 901 3726
rect 932 3723 941 3726
rect 964 3723 980 3726
rect 1060 3723 1085 3726
rect 1122 3723 1140 3726
rect 1188 3723 1213 3726
rect 1300 3723 1309 3726
rect 1314 3723 1340 3726
rect 1426 3723 1436 3726
rect 1458 3716 1461 3733
rect 1866 3726 1869 3736
rect 1892 3733 1901 3736
rect 1922 3727 1925 3735
rect 2018 3733 2028 3736
rect 2042 3733 2060 3736
rect 1498 3723 1508 3726
rect 1532 3723 1557 3726
rect 1594 3723 1604 3726
rect 1610 3723 1636 3726
rect 1452 3713 1461 3716
rect 1644 3713 1653 3716
rect 1666 3706 1669 3725
rect 1732 3723 1773 3726
rect 1780 3723 1789 3726
rect 1844 3723 1869 3726
rect 1916 3724 1925 3727
rect 1973 3723 1981 3726
rect 2090 3713 2093 3735
rect 2164 3733 2181 3736
rect 2196 3733 2205 3736
rect 2258 3733 2276 3736
rect 2300 3733 2325 3736
rect 2332 3733 2349 3736
rect 2380 3733 2405 3736
rect 2436 3733 2453 3736
rect 2484 3733 2509 3736
rect 2610 3733 2619 3736
rect 2650 3733 2659 3736
rect 2690 3733 2715 3736
rect 2722 3733 2739 3736
rect 2914 3733 2923 3736
rect 2949 3733 2957 3736
rect 2964 3733 2973 3736
rect 3012 3733 3021 3736
rect 3028 3733 3053 3736
rect 3082 3726 3085 3734
rect 3106 3733 3124 3736
rect 3180 3733 3189 3736
rect 3218 3726 3221 3734
rect 3250 3726 3253 3734
rect 2114 3723 2124 3726
rect 2204 3723 2221 3726
rect 2274 3723 2284 3726
rect 2402 3723 2419 3726
rect 2644 3723 2653 3726
rect 2684 3723 2693 3726
rect 2724 3723 2741 3726
rect 2890 3723 2900 3726
rect 3050 3723 3068 3726
rect 3082 3723 3093 3726
rect 3122 3723 3132 3726
rect 3154 3723 3163 3726
rect 3186 3723 3204 3726
rect 3218 3723 3229 3726
rect 3250 3723 3261 3726
rect 3282 3725 3285 3746
rect 3314 3743 3322 3746
rect 3378 3743 3388 3746
rect 3300 3733 3325 3736
rect 3332 3733 3341 3736
rect 3396 3733 3405 3736
rect 3684 3733 3693 3736
rect 3706 3733 3732 3736
rect 3756 3733 3765 3736
rect 3772 3733 3797 3736
rect 3994 3733 4020 3736
rect 4034 3733 4044 3736
rect 4204 3733 4213 3736
rect 4266 3734 4284 3736
rect 4266 3733 4285 3734
rect 4354 3733 4364 3736
rect 3404 3723 3413 3726
rect 3492 3723 3501 3726
rect 3540 3723 3549 3726
rect 3626 3723 3636 3726
rect 3722 3723 3740 3726
rect 3818 3723 3828 3726
rect 3858 3723 3884 3726
rect 4028 3723 4045 3726
rect 4082 3723 4108 3726
rect 4212 3723 4229 3726
rect 4282 3723 4285 3733
rect 4298 3723 4308 3726
rect 4338 3723 4372 3726
rect 2650 3716 2653 3723
rect 2108 3713 2117 3716
rect 2436 3713 2453 3716
rect 2650 3713 2661 3716
rect 3186 3713 3189 3723
rect 3258 3713 3261 3723
rect 3436 3713 3445 3716
rect 1658 3703 1669 3706
rect 3546 3706 3549 3723
rect 3546 3703 3565 3706
rect 14 3667 4434 3673
rect 1538 3636 1541 3646
rect 1538 3633 1564 3636
rect 1690 3633 1708 3636
rect 1802 3633 1836 3636
rect 308 3623 317 3626
rect 1626 3616 1629 3626
rect 1682 3623 1692 3626
rect 1716 3623 1725 3626
rect 1810 3623 1820 3626
rect 1844 3623 1853 3626
rect 2164 3623 2181 3626
rect 2356 3623 2365 3626
rect 2436 3623 2453 3626
rect 2578 3616 2581 3626
rect 2612 3623 2621 3626
rect 2733 3623 2741 3626
rect 210 3613 228 3616
rect 242 3613 252 3616
rect 314 3613 324 3616
rect 354 3613 364 3616
rect 596 3613 621 3616
rect 788 3613 813 3616
rect 844 3613 861 3616
rect 924 3613 949 3616
rect 980 3613 997 3616
rect 1018 3613 1029 3616
rect 1036 3613 1077 3616
rect 1106 3613 1140 3616
rect 1196 3613 1221 3616
rect 1252 3613 1277 3616
rect 1332 3613 1341 3616
rect 1356 3613 1373 3616
rect 234 3603 260 3606
rect 274 3603 284 3606
rect 322 3603 332 3606
rect 346 3603 356 3606
rect 858 3605 861 3613
rect 986 3603 996 3606
rect 1026 3605 1029 3613
rect 1074 3605 1077 3613
rect 1314 3603 1324 3606
rect 1338 3595 1341 3613
rect 1458 3606 1461 3614
rect 1484 3613 1493 3616
rect 1626 3613 1636 3616
rect 1650 3613 1668 3616
rect 1796 3613 1805 3616
rect 1892 3613 1901 3616
rect 1940 3613 1965 3616
rect 2002 3613 2020 3616
rect 2050 3613 2060 3616
rect 2092 3613 2101 3616
rect 2116 3613 2141 3616
rect 2234 3613 2253 3616
rect 2402 3613 2419 3616
rect 2442 3613 2460 3616
rect 2506 3613 2516 3616
rect 2530 3613 2541 3616
rect 2578 3613 2596 3616
rect 2250 3606 2253 3613
rect 2530 3607 2533 3613
rect 2610 3607 2613 3616
rect 1348 3603 1365 3606
rect 1370 3603 1380 3606
rect 1404 3603 1413 3606
rect 1444 3603 1461 3606
rect 1490 3603 1499 3606
rect 1532 3603 1541 3606
rect 1642 3603 1660 3606
rect 2066 3603 2084 3606
rect 2108 3603 2133 3606
rect 2228 3603 2245 3606
rect 2276 3603 2285 3606
rect 2300 3603 2317 3606
rect 2322 3603 2332 3606
rect 2356 3603 2373 3606
rect 2498 3603 2508 3606
rect 2322 3596 2325 3603
rect 2282 3593 2292 3596
rect 2306 3593 2325 3596
rect 2362 3593 2380 3596
rect 2618 3593 2621 3623
rect 2818 3616 2821 3636
rect 3546 3626 3549 3646
rect 3540 3623 3549 3626
rect 3748 3623 3757 3626
rect 2692 3613 2709 3616
rect 2764 3613 2773 3616
rect 2818 3613 2829 3616
rect 2882 3613 2907 3616
rect 2970 3613 2980 3616
rect 3002 3613 3012 3616
rect 3074 3613 3085 3616
rect 3106 3613 3132 3616
rect 3146 3613 3157 3616
rect 3178 3613 3188 3616
rect 2826 3607 2829 3613
rect 2733 3603 2749 3606
rect 2762 3603 2770 3606
rect 2852 3603 2861 3606
rect 2868 3603 2893 3606
rect 2924 3603 2933 3606
rect 2940 3603 2957 3606
rect 3028 3603 3045 3606
rect 3074 3605 3077 3613
rect 3092 3603 3117 3606
rect 3146 3605 3149 3613
rect 3210 3606 3213 3616
rect 3340 3613 3349 3616
rect 3378 3613 3403 3616
rect 3426 3613 3436 3616
rect 3508 3613 3517 3616
rect 3722 3613 3732 3616
rect 3746 3613 3773 3616
rect 3802 3613 3812 3616
rect 3956 3613 3973 3616
rect 4042 3613 4052 3616
rect 4082 3613 4100 3616
rect 4226 3613 4236 3616
rect 4266 3613 4276 3616
rect 3154 3603 3163 3606
rect 3170 3603 3179 3606
rect 3210 3603 3219 3606
rect 3226 3603 3258 3606
rect 3318 3603 3325 3606
rect 3332 3603 3341 3606
rect 3378 3596 3381 3613
rect 3770 3606 3773 3613
rect 3386 3603 3396 3606
rect 3452 3603 3461 3606
rect 3468 3603 3493 3606
rect 3500 3603 3509 3606
rect 3546 3603 3564 3606
rect 3620 3603 3629 3606
rect 3636 3603 3653 3606
rect 3684 3603 3701 3606
rect 3762 3605 3773 3606
rect 3762 3603 3772 3605
rect 3828 3603 3853 3606
rect 3860 3603 3877 3606
rect 3884 3603 3901 3606
rect 4018 3603 4028 3606
rect 4202 3603 4212 3606
rect 2666 3593 2674 3596
rect 3378 3593 3389 3596
rect 3474 3593 3492 3596
rect 3842 3593 3852 3596
rect 38 3567 4410 3573
rect 204 3543 221 3546
rect 916 3543 925 3546
rect 1082 3543 1092 3546
rect 1402 3536 1405 3545
rect 106 3526 109 3534
rect 140 3533 164 3536
rect 92 3523 109 3526
rect 178 3525 181 3536
rect 202 3533 229 3536
rect 282 3533 292 3536
rect 204 3523 213 3526
rect 226 3525 229 3533
rect 794 3526 797 3534
rect 842 3533 852 3536
rect 914 3533 940 3536
rect 954 3533 972 3536
rect 1020 3533 1029 3536
rect 1100 3533 1109 3536
rect 1154 3533 1164 3536
rect 1178 3533 1196 3536
rect 1244 3533 1261 3536
rect 1396 3533 1405 3536
rect 1442 3533 1452 3536
rect 1484 3533 1493 3536
rect 1514 3533 1524 3536
rect 1538 3526 1541 3545
rect 1650 3543 1676 3546
rect 1548 3533 1557 3536
rect 1594 3533 1604 3536
rect 1570 3526 1573 3533
rect 252 3523 269 3526
rect 306 3523 332 3526
rect 346 3523 364 3526
rect 418 3523 428 3526
rect 660 3523 677 3526
rect 716 3523 741 3526
rect 772 3523 797 3526
rect 804 3523 820 3526
rect 874 3523 892 3526
rect 956 3523 965 3526
rect 996 3523 1029 3526
rect 1066 3523 1076 3526
rect 1108 3523 1117 3526
rect 1156 3523 1165 3526
rect 1172 3523 1197 3526
rect 1300 3523 1325 3526
rect 1362 3523 1380 3526
rect 1450 3523 1460 3526
rect 1532 3523 1541 3526
rect 1556 3523 1573 3526
rect 1644 3523 1677 3526
rect 1762 3525 1765 3546
rect 1802 3543 1820 3546
rect 2042 3543 2052 3546
rect 2730 3536 2733 3556
rect 3770 3553 3781 3556
rect 2826 3536 2829 3546
rect 3706 3543 3716 3546
rect 3778 3536 3781 3553
rect 1828 3533 1845 3536
rect 1932 3533 1949 3536
rect 1964 3533 1981 3536
rect 266 3513 269 3523
rect 348 3513 357 3516
rect 388 3513 397 3516
rect 836 3513 845 3516
rect 876 3513 885 3516
rect 1026 3506 1029 3523
rect 1036 3513 1045 3516
rect 1700 3513 1709 3516
rect 1724 3513 1733 3516
rect 1772 3513 1781 3516
rect 1796 3513 1813 3516
rect 1842 3506 1845 3533
rect 2018 3526 2021 3534
rect 2092 3533 2117 3536
rect 2162 3533 2180 3536
rect 2212 3533 2229 3536
rect 2260 3533 2269 3536
rect 2274 3533 2291 3536
rect 2412 3533 2421 3536
rect 2466 3533 2500 3536
rect 2530 3533 2556 3536
rect 2586 3533 2612 3536
rect 2634 3533 2645 3536
rect 2678 3533 2685 3536
rect 2716 3533 2733 3536
rect 2738 3533 2747 3536
rect 2818 3533 2829 3536
rect 2956 3533 2965 3536
rect 2988 3533 2997 3536
rect 1882 3523 1916 3526
rect 2018 3523 2053 3526
rect 1876 3513 1901 3516
rect 2114 3506 2117 3533
rect 2642 3526 2645 3533
rect 2730 3526 2733 3533
rect 2818 3527 2821 3533
rect 3002 3527 3005 3536
rect 3042 3533 3060 3536
rect 3082 3533 3093 3536
rect 3124 3533 3133 3536
rect 3210 3533 3219 3536
rect 3330 3533 3340 3536
rect 3362 3533 3388 3536
rect 3410 3533 3418 3536
rect 3444 3533 3461 3536
rect 3484 3533 3493 3536
rect 3572 3533 3589 3536
rect 3620 3533 3629 3536
rect 3660 3533 3669 3536
rect 3764 3533 3773 3536
rect 3778 3533 3788 3536
rect 3812 3533 3821 3536
rect 3828 3533 3853 3536
rect 3884 3533 3893 3536
rect 3906 3533 3940 3536
rect 3994 3533 4028 3536
rect 4042 3533 4068 3536
rect 4106 3533 4116 3536
rect 2154 3523 2188 3526
rect 2290 3523 2300 3526
rect 2314 3523 2340 3526
rect 2354 3523 2388 3526
rect 2420 3523 2429 3526
rect 2468 3523 2485 3526
rect 2524 3523 2541 3526
rect 2642 3523 2659 3526
rect 2730 3523 2749 3526
rect 2834 3523 2844 3526
rect 2866 3523 2875 3526
rect 2954 3523 2964 3526
rect 2148 3513 2173 3516
rect 2260 3513 2277 3516
rect 2316 3513 2325 3516
rect 2356 3513 2373 3516
rect 1026 3503 1052 3506
rect 1698 3503 1716 3506
rect 1770 3503 1788 3506
rect 1842 3503 1868 3506
rect 2114 3503 2140 3506
rect 2530 3503 2533 3523
rect 2678 3513 2685 3516
rect 2773 3513 2781 3516
rect 2860 3513 2869 3516
rect 2866 3493 2869 3513
rect 3090 3483 3093 3533
rect 3162 3523 3179 3526
rect 3218 3523 3226 3526
rect 3442 3523 3460 3526
rect 3538 3523 3548 3526
rect 3618 3523 3644 3526
rect 3658 3523 3684 3526
rect 3778 3523 3796 3526
rect 3850 3523 3868 3526
rect 3948 3523 3957 3526
rect 4036 3523 4061 3526
rect 4106 3523 4124 3526
rect 4140 3523 4149 3526
rect 3164 3513 3173 3516
rect 3765 3513 3773 3516
rect 14 3467 4434 3473
rect 1666 3433 1676 3436
rect 1722 3433 1748 3436
rect 1826 3433 1837 3436
rect 860 3423 877 3426
rect 1412 3423 1421 3426
rect 1452 3423 1469 3426
rect 1650 3423 1660 3426
rect 1684 3423 1693 3426
rect 116 3413 141 3416
rect 186 3413 196 3416
rect 210 3413 228 3416
rect 234 3413 252 3416
rect 266 3413 309 3416
rect 338 3413 357 3416
rect 580 3413 589 3416
rect 628 3413 653 3416
rect 684 3413 701 3416
rect 740 3413 765 3416
rect 796 3413 821 3416
rect 828 3413 844 3416
rect 1028 3413 1053 3416
rect 1204 3413 1229 3416
rect 1316 3413 1341 3416
rect 1458 3413 1484 3416
rect 1538 3413 1548 3416
rect 1586 3413 1596 3416
rect 178 3403 188 3406
rect 306 3405 309 3413
rect 354 3405 357 3413
rect 818 3405 821 3413
rect 1722 3406 1725 3433
rect 1786 3423 1796 3426
rect 1820 3423 1829 3426
rect 1834 3425 1837 3433
rect 2018 3426 2021 3436
rect 2122 3433 2157 3436
rect 1860 3423 1885 3426
rect 1916 3423 1925 3426
rect 2004 3423 2021 3426
rect 2138 3423 2148 3426
rect 1882 3416 1885 3423
rect 2138 3416 2141 3423
rect 1780 3413 1804 3416
rect 1882 3413 1900 3416
rect 1970 3413 1988 3416
rect 2010 3413 2029 3416
rect 2060 3413 2085 3416
rect 2092 3413 2101 3416
rect 2116 3413 2141 3416
rect 2154 3415 2157 3433
rect 2210 3433 2236 3436
rect 2258 3433 2284 3436
rect 2172 3423 2181 3426
rect 2026 3406 2029 3413
rect 2210 3406 2213 3433
rect 2220 3423 2229 3426
rect 2292 3423 2309 3426
rect 2461 3423 2477 3426
rect 2338 3416 2341 3423
rect 2418 3416 2421 3423
rect 2522 3416 2525 3426
rect 2708 3423 2717 3426
rect 2868 3423 2885 3426
rect 3652 3423 3661 3426
rect 2298 3413 2324 3416
rect 2338 3413 2357 3416
rect 2418 3413 2429 3416
rect 2516 3413 2525 3416
rect 2570 3413 2587 3416
rect 2762 3413 2787 3416
rect 2842 3413 2852 3416
rect 2866 3413 2885 3416
rect 2988 3413 2997 3416
rect 3074 3413 3083 3416
rect 3106 3413 3115 3416
rect 3234 3413 3244 3416
rect 3266 3413 3274 3416
rect 3314 3413 3322 3416
rect 3394 3413 3403 3416
rect 3690 3413 3701 3416
rect 3738 3413 3748 3416
rect 3788 3413 3805 3416
rect 3834 3413 3852 3416
rect 3962 3413 3972 3416
rect 4002 3413 4012 3416
rect 4068 3413 4077 3416
rect 4170 3413 4180 3416
rect 4210 3413 4220 3416
rect 4250 3413 4268 3416
rect 866 3403 892 3406
rect 906 3403 932 3406
rect 986 3403 1004 3406
rect 1098 3403 1108 3406
rect 1378 3403 1388 3406
rect 1524 3403 1541 3406
rect 1572 3403 1588 3406
rect 1610 3403 1620 3406
rect 1708 3403 1725 3406
rect 1882 3403 1892 3406
rect 1916 3403 1933 3406
rect 1940 3403 1965 3406
rect 2004 3403 2021 3406
rect 2026 3403 2036 3406
rect 2066 3403 2084 3406
rect 2108 3403 2141 3406
rect 2196 3403 2213 3406
rect 2380 3403 2389 3406
rect 2474 3403 2492 3406
rect 2508 3403 2525 3406
rect 1690 3393 1700 3396
rect 2018 3393 2028 3396
rect 2178 3393 2188 3396
rect 2570 3393 2573 3413
rect 2882 3406 2885 3413
rect 2618 3403 2644 3406
rect 2714 3403 2731 3406
rect 2750 3403 2773 3406
rect 2804 3403 2821 3406
rect 2834 3403 2844 3406
rect 2868 3403 2877 3406
rect 2882 3403 2900 3406
rect 2916 3403 2925 3406
rect 2962 3403 2980 3406
rect 2986 3403 2996 3406
rect 3034 3403 3044 3406
rect 3066 3403 3076 3406
rect 3114 3403 3124 3406
rect 3180 3403 3189 3406
rect 3226 3403 3236 3406
rect 3262 3403 3277 3406
rect 3302 3403 3309 3406
rect 3354 3403 3362 3406
rect 3474 3403 3484 3406
rect 3506 3403 3522 3406
rect 3690 3405 3693 3413
rect 3724 3403 3733 3406
rect 3765 3403 3773 3406
rect 3780 3403 3805 3406
rect 3868 3403 3901 3406
rect 3908 3403 3925 3406
rect 3938 3403 3948 3406
rect 4186 3403 4196 3406
rect 4244 3403 4253 3406
rect 2962 3393 2972 3396
rect 3874 3393 3900 3396
rect 38 3367 4410 3373
rect 1292 3343 1309 3346
rect 1484 3343 1493 3346
rect 2010 3343 2028 3346
rect 970 3333 980 3336
rect 1002 3333 1036 3336
rect 1114 3333 1124 3336
rect 1266 3333 1276 3336
rect 172 3323 197 3326
rect 292 3323 309 3326
rect 348 3323 365 3326
rect 404 3323 413 3326
rect 460 3323 477 3326
rect 580 3323 597 3326
rect 756 3323 781 3326
rect 876 3323 901 3326
rect 938 3323 964 3326
rect 1004 3323 1013 3326
rect 1060 3323 1093 3326
rect 1114 3315 1117 3333
rect 1306 3326 1309 3343
rect 1348 3333 1365 3336
rect 1394 3333 1412 3336
rect 1442 3333 1468 3336
rect 1570 3333 1580 3336
rect 1770 3333 1796 3336
rect 1820 3333 1829 3336
rect 1842 3333 1851 3336
rect 1876 3333 1901 3336
rect 1914 3333 1940 3336
rect 1946 3333 1980 3336
rect 2036 3333 2053 3336
rect 1196 3323 1221 3326
rect 1306 3323 1317 3326
rect 1394 3325 1397 3333
rect 1570 3323 1588 3326
rect 1604 3323 1621 3326
rect 1490 3313 1509 3316
rect 1524 3313 1533 3316
rect 1618 3313 1621 3323
rect 1628 3313 1637 3316
rect 1658 3313 1668 3316
rect 1674 3306 1677 3325
rect 1772 3323 1781 3326
rect 1948 3323 1973 3326
rect 1978 3323 1988 3326
rect 1698 3313 1708 3316
rect 1732 3313 1749 3316
rect 1820 3313 1845 3316
rect 1876 3313 1885 3316
rect 2050 3306 2053 3333
rect 2098 3323 2101 3346
rect 2106 3343 2124 3346
rect 2138 3343 2156 3346
rect 2132 3333 2157 3336
rect 2178 3333 2196 3336
rect 2362 3333 2388 3336
rect 2426 3333 2429 3356
rect 2474 3336 2477 3346
rect 2434 3333 2444 3336
rect 2474 3333 2508 3336
rect 2538 3333 2572 3336
rect 2602 3333 2628 3336
rect 2652 3333 2669 3336
rect 2682 3333 2707 3336
rect 2732 3333 2741 3336
rect 2746 3333 2763 3336
rect 2780 3333 2797 3336
rect 2850 3333 2876 3336
rect 2898 3333 2940 3336
rect 3108 3333 3117 3336
rect 2746 3326 2749 3333
rect 3122 3326 3125 3346
rect 3842 3343 3852 3346
rect 3866 3343 3876 3346
rect 3162 3333 3179 3336
rect 3218 3333 3228 3336
rect 3258 3333 3268 3336
rect 3294 3333 3301 3336
rect 3332 3333 3349 3336
rect 3468 3333 3477 3336
rect 3482 3333 3500 3336
rect 3518 3333 3525 3336
rect 3530 3333 3540 3336
rect 3564 3333 3573 3336
rect 3604 3333 3613 3336
rect 3618 3326 3621 3335
rect 3676 3333 3693 3336
rect 3762 3333 3772 3336
rect 3796 3333 3805 3336
rect 3836 3333 3853 3336
rect 3860 3333 3877 3336
rect 3884 3333 3893 3336
rect 2140 3323 2149 3326
rect 2172 3323 2204 3326
rect 2362 3323 2396 3326
rect 2532 3323 2557 3326
rect 2618 3323 2635 3326
rect 2698 3323 2715 3326
rect 2738 3323 2749 3326
rect 2858 3323 2868 3326
rect 2902 3323 2909 3326
rect 2914 3323 2932 3326
rect 2058 3313 2068 3316
rect 2092 3313 2117 3316
rect 2252 3313 2269 3316
rect 2314 3313 2332 3316
rect 2356 3313 2381 3316
rect 2412 3313 2429 3316
rect 2468 3313 2493 3316
rect 1490 3303 1516 3306
rect 1530 3303 1556 3306
rect 1666 3303 1677 3306
rect 1706 3303 1724 3306
rect 2050 3303 2084 3306
rect 2210 3303 2244 3306
rect 2258 3303 2292 3306
rect 2306 3303 2348 3306
rect 2698 3293 2701 3323
rect 2733 3313 2749 3316
rect 2844 3313 2861 3316
rect 3010 3313 3020 3316
rect 3026 3306 3029 3325
rect 3050 3323 3060 3326
rect 3082 3323 3092 3326
rect 3114 3323 3125 3326
rect 3162 3323 3172 3326
rect 3298 3323 3314 3326
rect 3386 3323 3396 3326
rect 3562 3323 3588 3326
rect 3602 3323 3621 3326
rect 3642 3323 3660 3326
rect 3730 3323 3740 3326
rect 3762 3323 3773 3326
rect 3810 3323 3820 3326
rect 3948 3323 3965 3326
rect 4010 3323 4020 3326
rect 4026 3323 4036 3326
rect 4082 3323 4100 3326
rect 4218 3323 4228 3326
rect 4258 3323 4276 3326
rect 3114 3316 3117 3323
rect 3762 3316 3765 3323
rect 3108 3313 3117 3316
rect 3122 3313 3132 3316
rect 3756 3313 3765 3316
rect 3002 3303 3029 3306
rect 3130 3303 3148 3306
rect 14 3267 4434 3273
rect 642 3216 645 3236
rect 940 3223 965 3226
rect 986 3216 989 3236
rect 1098 3233 1108 3236
rect 1634 3233 1668 3236
rect 1682 3233 1693 3236
rect 1698 3233 1708 3236
rect 1730 3233 1748 3236
rect 1762 3233 1788 3236
rect 2290 3233 2332 3236
rect 2858 3233 2869 3236
rect 2914 3233 2948 3236
rect 2986 3233 3012 3236
rect 3066 3233 3083 3236
rect 3098 3233 3115 3236
rect 3138 3233 3165 3236
rect 1052 3223 1061 3226
rect 1548 3223 1557 3226
rect 1628 3223 1645 3226
rect 1676 3223 1685 3226
rect 1690 3225 1693 3233
rect 1716 3223 1725 3226
rect 1732 3223 1741 3226
rect 1988 3223 1997 3226
rect 2156 3223 2165 3226
rect 2340 3223 2349 3226
rect 2388 3223 2413 3226
rect 2508 3223 2533 3226
rect 116 3213 141 3216
rect 186 3213 220 3216
rect 226 3213 236 3216
rect 306 3213 316 3216
rect 346 3206 349 3214
rect 410 3213 420 3216
rect 442 3206 445 3214
rect 524 3213 541 3216
rect 580 3213 589 3216
rect 612 3213 621 3216
rect 642 3213 660 3216
rect 674 3213 708 3216
rect 722 3213 740 3216
rect 788 3213 805 3216
rect 826 3213 868 3216
rect 892 3213 901 3216
rect 980 3213 989 3216
rect 1050 3213 1100 3216
rect 1172 3213 1197 3216
rect 1228 3213 1245 3216
rect 1274 3213 1292 3216
rect 1298 3213 1315 3216
rect 1340 3213 1357 3216
rect 1484 3213 1501 3216
rect 1498 3206 1501 3213
rect 1554 3206 1557 3223
rect 1562 3213 1572 3216
rect 1596 3213 1605 3216
rect 1620 3213 1629 3216
rect 1810 3213 1828 3216
rect 1884 3213 1917 3216
rect 1946 3213 1972 3216
rect 2108 3213 2125 3216
rect 2154 3213 2196 3216
rect 2258 3213 2268 3216
rect 1602 3206 1605 3213
rect 338 3203 349 3206
rect 434 3203 445 3206
rect 468 3203 493 3206
rect 516 3203 556 3206
rect 578 3203 604 3206
rect 676 3203 693 3206
rect 770 3203 780 3206
rect 794 3203 804 3206
rect 828 3203 837 3206
rect 874 3203 884 3206
rect 890 3203 916 3206
rect 946 3203 972 3206
rect 1018 3203 1028 3206
rect 1052 3203 1061 3206
rect 1298 3203 1324 3206
rect 1498 3203 1508 3206
rect 1554 3203 1564 3206
rect 1578 3203 1588 3206
rect 1602 3203 1612 3206
rect 1802 3203 1820 3206
rect 1882 3203 1916 3206
rect 1954 3203 1964 3206
rect 1988 3203 2021 3206
rect 2028 3203 2045 3206
rect 2106 3203 2132 3206
rect 2212 3203 2237 3206
rect 2244 3203 2261 3206
rect 2346 3203 2349 3223
rect 2578 3216 2581 3226
rect 2628 3223 2653 3226
rect 2684 3223 2701 3226
rect 2852 3223 2861 3226
rect 2866 3216 2869 3233
rect 2986 3216 2989 3233
rect 2996 3223 3005 3226
rect 3042 3223 3068 3226
rect 3102 3223 3109 3226
rect 3130 3223 3156 3226
rect 2410 3213 2420 3216
rect 2474 3213 2492 3216
rect 2506 3213 2540 3216
rect 2578 3213 2612 3216
rect 2658 3213 2668 3216
rect 2682 3213 2708 3216
rect 2746 3213 2763 3216
rect 2796 3213 2805 3216
rect 2810 3213 2836 3216
rect 2866 3213 2876 3216
rect 2962 3213 2989 3216
rect 3026 3213 3061 3216
rect 3162 3215 3165 3233
rect 3378 3216 3381 3236
rect 3420 3223 3429 3226
rect 3556 3223 3565 3226
rect 3668 3223 3685 3226
rect 3812 3223 3821 3226
rect 3198 3213 3213 3216
rect 3282 3206 3285 3216
rect 3330 3213 3340 3216
rect 3372 3213 3381 3216
rect 3418 3213 3444 3216
rect 3466 3213 3476 3216
rect 3554 3213 3580 3216
rect 3628 3213 3645 3216
rect 3708 3213 3717 3216
rect 3732 3213 3749 3216
rect 3810 3213 3836 3216
rect 3940 3213 3949 3216
rect 4066 3213 4084 3216
rect 4210 3213 4220 3216
rect 4250 3213 4268 3216
rect 2418 3203 2428 3206
rect 2458 3203 2483 3206
rect 2522 3203 2548 3206
rect 2634 3203 2659 3206
rect 2690 3203 2715 3206
rect 2733 3203 2765 3206
rect 2818 3203 2828 3206
rect 2902 3203 2925 3206
rect 3244 3203 3253 3206
rect 3266 3203 3298 3206
rect 3322 3203 3346 3206
rect 3420 3203 3429 3206
rect 3522 3203 3532 3206
rect 3596 3203 3613 3206
rect 3620 3203 3637 3206
rect 3700 3203 3709 3206
rect 3724 3203 3741 3206
rect 3772 3203 3781 3206
rect 3812 3203 3821 3206
rect 3884 3203 3901 3206
rect 3908 3203 3925 3206
rect 3986 3203 4012 3206
rect 4186 3203 4196 3206
rect 4244 3203 4253 3206
rect 338 3183 341 3203
rect 434 3183 437 3203
rect 490 3196 493 3203
rect 490 3193 508 3196
rect 3250 3195 3253 3203
rect 3426 3193 3429 3203
rect 3602 3193 3612 3196
rect 3674 3193 3692 3196
rect 3778 3183 3781 3203
rect 3858 3193 3876 3196
rect 3890 3193 3900 3196
rect 38 3167 4410 3173
rect 562 3143 572 3146
rect 778 3143 788 3146
rect 1130 3143 1140 3146
rect 282 3133 292 3136
rect 602 3133 612 3136
rect 778 3126 781 3143
rect 1298 3136 1301 3156
rect 1810 3143 1820 3146
rect 1866 3143 1892 3146
rect 1906 3143 1916 3146
rect 1970 3143 1980 3146
rect 2090 3136 2093 3156
rect 3738 3143 3764 3146
rect 4194 3136 4197 3156
rect 818 3133 828 3136
rect 932 3133 941 3136
rect 1020 3133 1029 3136
rect 1148 3133 1165 3136
rect 1266 3133 1276 3136
rect 1298 3133 1308 3136
rect 1444 3133 1453 3136
rect 1554 3133 1564 3136
rect 1596 3133 1605 3136
rect 1730 3133 1755 3136
rect 1900 3133 1917 3136
rect 1924 3133 1949 3136
rect 1964 3133 1981 3136
rect 1988 3133 2013 3136
rect 2084 3133 2093 3136
rect 2148 3133 2165 3136
rect 2180 3133 2197 3136
rect 2226 3133 2236 3136
rect 2314 3133 2340 3136
rect 2396 3133 2429 3136
rect 2452 3133 2469 3136
rect 2538 3133 2565 3136
rect 2650 3133 2660 3136
rect 2714 3133 2724 3136
rect 2868 3133 2901 3136
rect 3098 3133 3116 3136
rect 3130 3133 3140 3136
rect 3170 3133 3180 3136
rect 3194 3133 3219 3136
rect 3242 3133 3276 3136
rect 3298 3133 3322 3136
rect 3350 3133 3373 3136
rect 3418 3133 3436 3136
rect 3458 3133 3492 3136
rect 3522 3133 3540 3136
rect 3564 3133 3581 3136
rect 3612 3133 3637 3136
rect 3772 3133 3805 3136
rect 3972 3133 3997 3136
rect 4044 3133 4069 3136
rect 4170 3133 4180 3136
rect 4194 3133 4204 3136
rect 938 3126 941 3133
rect 2194 3126 2197 3133
rect 124 3123 149 3126
rect 186 3123 228 3126
rect 644 3123 677 3126
rect 716 3123 725 3126
rect 772 3123 781 3126
rect 812 3123 829 3126
rect 938 3123 948 3126
rect 970 3123 980 3126
rect 1204 3123 1229 3126
rect 1260 3123 1277 3126
rect 1284 3123 1309 3126
rect 1346 3123 1380 3126
rect 1404 3123 1421 3126
rect 1492 3123 1517 3126
rect 1562 3123 1572 3126
rect 1602 3123 1620 3126
rect 1650 3123 1668 3126
rect 1932 3123 1949 3126
rect 2002 3123 2020 3126
rect 2194 3123 2204 3126
rect 2234 3123 2244 3126
rect 2306 3123 2348 3126
rect 2370 3123 2380 3126
rect 2410 3123 2428 3126
rect 2498 3123 2508 3126
rect 2538 3125 2541 3133
rect 2642 3123 2668 3126
rect 2714 3116 2717 3133
rect 2754 3123 2780 3126
rect 2938 3123 2964 3126
rect 3138 3123 3147 3126
rect 3188 3123 3205 3126
rect 3244 3123 3261 3126
rect 3346 3123 3370 3126
rect 3410 3123 3428 3126
rect 3466 3123 3484 3126
rect 3530 3123 3548 3126
rect 3562 3123 3596 3126
rect 3676 3123 3685 3126
rect 3844 3123 3853 3126
rect 3906 3123 3932 3126
rect 2300 3113 2333 3116
rect 2700 3113 2717 3116
rect 2882 3113 2908 3116
rect 2970 3113 2980 3116
rect 3010 3113 3028 3116
rect 3052 3113 3061 3116
rect 3066 3106 3069 3115
rect 3092 3113 3109 3116
rect 3994 3113 3997 3133
rect 4188 3123 4197 3126
rect 4202 3123 4212 3126
rect 4242 3123 4252 3126
rect 2602 3103 2619 3106
rect 2682 3103 2692 3106
rect 2882 3103 2924 3106
rect 3018 3103 3044 3106
rect 3058 3103 3069 3106
rect 14 3067 4434 3073
rect 1178 3033 1195 3036
rect 180 3023 189 3026
rect 220 3023 237 3026
rect 1162 3023 1180 3026
rect 1300 3023 1309 3026
rect 1612 3023 1629 3026
rect 1700 3023 1709 3026
rect 1162 3016 1165 3023
rect 2154 3016 2157 3036
rect 2474 3033 2492 3036
rect 2562 3033 2587 3036
rect 2706 3033 2733 3036
rect 2754 3033 2772 3036
rect 2890 3033 2908 3036
rect 2994 3033 3020 3036
rect 2636 3023 2653 3026
rect 2706 3023 2724 3026
rect 108 3013 141 3016
rect 276 3013 293 3016
rect 396 3013 413 3016
rect 500 3013 525 3016
rect 604 3013 637 3016
rect 676 3013 693 3016
rect 1092 3013 1109 3016
rect 1132 3013 1165 3016
rect 1210 3013 1220 3016
rect 1250 3013 1268 3016
rect 1436 3013 1453 3016
rect 1546 3013 1580 3016
rect 1660 3013 1708 3016
rect 1764 3013 1797 3016
rect 1852 3013 1885 3016
rect 1890 3013 1900 3016
rect 2044 3013 2060 3016
rect 2098 3013 2116 3016
rect 2148 3013 2157 3016
rect 522 3006 525 3013
rect 2162 3006 2165 3014
rect 132 3003 149 3006
rect 226 3003 244 3006
rect 292 3003 317 3006
rect 346 3003 364 3006
rect 450 3003 468 3006
rect 522 3003 533 3006
rect 562 3003 572 3006
rect 1066 3003 1084 3006
rect 1098 3003 1108 3006
rect 1157 3003 1173 3006
rect 1242 3003 1260 3006
rect 1380 3003 1397 3006
rect 1554 3003 1572 3006
rect 1804 3003 1821 3006
rect 2002 3003 2020 3006
rect 2090 3003 2124 3006
rect 2146 3003 2165 3006
rect 2202 3013 2228 3016
rect 2394 3013 2402 3016
rect 2428 3013 2453 3016
rect 2602 3013 2620 3016
rect 2730 3015 2733 3033
rect 2836 3023 2845 3026
rect 2892 3023 2901 3026
rect 3060 3023 3069 3026
rect 2866 3013 2884 3016
rect 306 2993 316 2996
rect 522 2993 532 2996
rect 2202 2993 2205 3013
rect 2210 3003 2220 3006
rect 2244 3003 2253 3006
rect 2410 3003 2420 3006
rect 2532 3003 2541 3006
rect 2602 3003 2605 3013
rect 2668 3003 2685 3006
rect 2692 3003 2717 3006
rect 2794 3003 2812 3006
rect 2866 3003 2869 3013
rect 2426 2993 2452 2996
rect 2506 2993 2524 2996
rect 2674 2993 2684 2996
rect 2786 2993 2804 2996
rect 2898 2993 2901 3014
rect 2922 3013 2956 3016
rect 2962 3013 2972 3016
rect 3108 3013 3133 3016
rect 3164 3013 3181 3016
rect 3188 3013 3197 3016
rect 3596 3013 3621 3016
rect 3652 3013 3677 3016
rect 3684 3013 3693 3016
rect 3748 3013 3757 3016
rect 3828 3013 3837 3016
rect 3906 3013 3916 3016
rect 3946 3013 3964 3016
rect 4082 3013 4100 3016
rect 4130 3013 4140 3016
rect 4146 3013 4172 3016
rect 4202 3013 4212 3016
rect 2922 3003 2948 3006
rect 3178 3005 3181 3013
rect 3674 3005 3677 3013
rect 3946 3006 3949 3013
rect 3730 3003 3740 3006
rect 3940 3003 3949 3006
rect 4082 3003 4092 3006
rect 4146 3003 4164 3006
rect 38 2967 4410 2973
rect 290 2926 293 2935
rect 650 2933 676 2936
rect 780 2933 789 2936
rect 810 2933 828 2936
rect 938 2933 948 2936
rect 980 2933 989 2936
rect 1650 2933 1660 2936
rect 1676 2933 1693 2936
rect 1906 2933 1932 2936
rect 1978 2933 1988 2936
rect 786 2926 789 2933
rect 212 2923 237 2926
rect 268 2923 293 2926
rect 300 2923 309 2926
rect 356 2923 381 2926
rect 658 2923 684 2926
rect 714 2923 749 2926
rect 786 2923 804 2926
rect 866 2923 875 2926
rect 882 2923 908 2926
rect 1252 2923 1261 2926
rect 1308 2923 1317 2926
rect 1364 2923 1373 2926
rect 1572 2923 1597 2926
rect 1628 2923 1637 2926
rect 1642 2923 1652 2926
rect 1732 2923 1757 2926
rect 1957 2923 1965 2926
rect 1970 2923 1980 2926
rect 2012 2923 2021 2926
rect 2034 2925 2037 2936
rect 2060 2933 2085 2936
rect 2130 2933 2172 2936
rect 2594 2933 2604 2936
rect 2970 2933 2980 2936
rect 2970 2926 2973 2933
rect 3154 2926 3157 2935
rect 3210 2933 3220 2936
rect 2132 2923 2141 2926
rect 2146 2923 2164 2926
rect 2202 2923 2236 2926
rect 2420 2923 2445 2926
rect 2532 2923 2557 2926
rect 2612 2923 2621 2926
rect 2628 2923 2645 2926
rect 2684 2923 2701 2926
rect 2796 2923 2813 2926
rect 2908 2923 2933 2926
rect 2964 2923 2973 2926
rect 3084 2923 3109 2926
rect 3140 2923 3157 2926
rect 3164 2923 3173 2926
rect 3210 2923 3228 2926
rect 3258 2923 3268 2926
rect 3274 2923 3292 2926
rect 3322 2923 3332 2926
rect 3396 2923 3405 2926
rect 3498 2923 3508 2926
rect 3562 2923 3572 2926
rect 3690 2923 3708 2926
rect 3930 2923 3940 2926
rect 4050 2923 4060 2926
rect 4090 2923 4100 2926
rect 4196 2923 4205 2926
rect 4218 2923 4228 2926
rect 4258 2923 4268 2926
rect 14 2867 4434 2873
rect 2930 2853 2949 2856
rect 570 2816 573 2846
rect 1274 2817 1277 2826
rect 116 2813 141 2816
rect 172 2813 189 2816
rect 196 2813 205 2816
rect 250 2813 285 2816
rect 322 2813 348 2816
rect 484 2813 501 2816
rect 516 2813 525 2816
rect 570 2813 580 2816
rect 618 2813 660 2816
rect 716 2813 733 2816
rect 770 2813 788 2816
rect 844 2813 861 2816
rect 898 2813 925 2816
rect 932 2813 949 2816
rect 186 2805 189 2813
rect 258 2803 268 2806
rect 282 2805 285 2813
rect 330 2803 340 2806
rect 426 2803 436 2806
rect 522 2805 525 2813
rect 556 2803 573 2806
rect 578 2803 588 2806
rect 618 2803 627 2806
rect 686 2803 701 2806
rect 722 2803 732 2806
rect 770 2803 780 2806
rect 838 2803 853 2806
rect 892 2803 901 2806
rect 946 2805 949 2813
rect 994 2813 1012 2816
rect 1076 2813 1101 2816
rect 1132 2813 1149 2816
rect 1226 2813 1243 2816
rect 1260 2814 1277 2817
rect 1626 2816 1629 2836
rect 1698 2816 1701 2826
rect 1794 2816 1797 2846
rect 1282 2813 1300 2816
rect 1330 2813 1340 2816
rect 1402 2813 1420 2816
rect 1458 2814 1468 2816
rect 1458 2813 1469 2814
rect 1498 2813 1516 2816
rect 1554 2813 1581 2816
rect 1586 2813 1596 2816
rect 1626 2813 1652 2816
rect 1698 2813 1724 2816
rect 1738 2813 1748 2816
rect 1794 2813 1805 2816
rect 1842 2813 1851 2816
rect 2026 2813 2060 2816
rect 2074 2813 2108 2816
rect 2122 2813 2156 2816
rect 2220 2813 2229 2816
rect 2282 2813 2316 2816
rect 2388 2813 2405 2816
rect 2476 2813 2493 2816
rect 2580 2813 2605 2816
rect 2668 2813 2685 2816
rect 2756 2813 2765 2816
rect 2868 2813 2893 2816
rect 2924 2813 2949 2816
rect 3092 2813 3117 2816
rect 3148 2813 3173 2816
rect 3226 2813 3252 2816
rect 3282 2813 3292 2816
rect 3386 2813 3396 2816
rect 3476 2813 3485 2816
rect 3532 2813 3541 2816
rect 3580 2813 3589 2816
rect 3764 2813 3773 2816
rect 3836 2813 3845 2816
rect 3850 2813 3860 2816
rect 3994 2813 4020 2816
rect 4060 2813 4077 2816
rect 4124 2813 4133 2816
rect 4138 2813 4148 2816
rect 994 2806 997 2813
rect 980 2803 997 2806
rect 1146 2806 1149 2813
rect 1466 2806 1469 2813
rect 1554 2806 1557 2813
rect 1698 2806 1701 2813
rect 1146 2803 1154 2806
rect 1324 2803 1341 2806
rect 1370 2803 1380 2806
rect 1444 2803 1469 2806
rect 1490 2803 1524 2806
rect 1540 2803 1557 2806
rect 1578 2803 1588 2806
rect 1634 2803 1642 2806
rect 1684 2803 1701 2806
rect 1730 2803 1739 2806
rect 1802 2805 1805 2813
rect 1858 2803 1876 2806
rect 1908 2803 1925 2806
rect 2042 2803 2052 2806
rect 2332 2803 2341 2806
rect 2482 2803 2492 2806
rect 2674 2803 2684 2806
rect 2954 2803 2964 2806
rect 2986 2803 3012 2806
rect 3170 2805 3173 2813
rect 3220 2803 3237 2806
rect 3298 2803 3324 2806
rect 3354 2803 3372 2806
rect 3538 2803 3556 2806
rect 3578 2803 3604 2806
rect 3778 2803 3796 2806
rect 3818 2803 3828 2806
rect 3994 2803 4012 2806
rect 4058 2803 4076 2806
rect 690 2793 699 2796
rect 818 2793 828 2796
rect 850 2793 853 2803
rect 898 2793 901 2803
rect 2980 2793 2997 2796
rect 3538 2793 3541 2803
rect 38 2767 4410 2773
rect 666 2743 675 2746
rect 170 2733 180 2736
rect 402 2726 405 2735
rect 562 2733 572 2736
rect 738 2733 754 2736
rect 778 2733 794 2736
rect 812 2733 821 2736
rect 826 2733 844 2736
rect 860 2733 869 2736
rect 1170 2726 1173 2735
rect 108 2723 125 2726
rect 164 2723 181 2726
rect 250 2723 268 2726
rect 332 2723 357 2726
rect 388 2723 405 2726
rect 412 2723 421 2726
rect 500 2723 525 2726
rect 556 2723 573 2726
rect 610 2723 636 2726
rect 698 2723 707 2726
rect 868 2723 877 2726
rect 954 2723 964 2726
rect 1110 2723 1133 2726
rect 1164 2723 1173 2726
rect 1202 2723 1205 2734
rect 1252 2733 1261 2736
rect 1322 2733 1331 2736
rect 1466 2733 1474 2736
rect 1354 2726 1357 2733
rect 1498 2731 1501 2733
rect 1506 2726 1509 2756
rect 2186 2743 2196 2746
rect 2420 2743 2429 2746
rect 3802 2743 3821 2746
rect 3802 2736 3805 2743
rect 4034 2736 4037 2746
rect 1666 2733 1674 2736
rect 1962 2733 1972 2736
rect 2186 2733 2203 2736
rect 2236 2733 2253 2736
rect 2290 2733 2308 2736
rect 2314 2733 2332 2736
rect 2610 2733 2620 2736
rect 1642 2726 1645 2733
rect 1212 2723 1221 2726
rect 1306 2723 1315 2726
rect 1316 2723 1325 2726
rect 1330 2723 1338 2726
rect 1354 2723 1365 2726
rect 1460 2723 1469 2726
rect 1498 2723 1509 2726
rect 1610 2723 1628 2726
rect 1642 2723 1653 2726
rect 1662 2723 1669 2726
rect 1362 2703 1365 2723
rect 1498 2717 1501 2723
rect 1610 2713 1613 2723
rect 1698 2721 1701 2724
rect 1804 2723 1813 2726
rect 2020 2723 2029 2726
rect 2220 2723 2229 2726
rect 1810 2703 1813 2723
rect 2250 2706 2253 2733
rect 2314 2725 2317 2733
rect 2770 2726 2773 2735
rect 2842 2733 2860 2736
rect 3004 2733 3028 2736
rect 3058 2733 3076 2736
rect 3090 2733 3116 2736
rect 3250 2733 3261 2736
rect 3418 2733 3436 2736
rect 3468 2733 3477 2736
rect 3258 2726 3261 2733
rect 3474 2726 3477 2733
rect 3506 2733 3524 2736
rect 3546 2733 3581 2736
rect 3604 2733 3613 2736
rect 3626 2733 3636 2736
rect 3650 2733 3668 2736
rect 3788 2733 3805 2736
rect 3810 2733 3828 2736
rect 3842 2733 3860 2736
rect 3898 2733 3940 2736
rect 4034 2733 4052 2736
rect 4082 2733 4092 2736
rect 4154 2733 4164 2736
rect 3506 2726 3509 2733
rect 3578 2726 3581 2733
rect 2322 2723 2338 2726
rect 2386 2723 2396 2726
rect 2548 2723 2573 2726
rect 2610 2723 2628 2726
rect 2708 2723 2733 2726
rect 2764 2723 2773 2726
rect 2780 2723 2789 2726
rect 2826 2723 2836 2726
rect 2922 2723 2941 2726
rect 3010 2723 3020 2726
rect 3044 2723 3053 2726
rect 3092 2723 3101 2726
rect 3132 2723 3149 2726
rect 3188 2723 3213 2726
rect 3244 2723 3253 2726
rect 3258 2723 3276 2726
rect 3426 2723 3444 2726
rect 3474 2723 3509 2726
rect 3618 2723 3644 2726
rect 3650 2723 3676 2726
rect 3706 2723 3748 2726
rect 3754 2723 3764 2726
rect 3802 2723 3836 2726
rect 3842 2723 3868 2726
rect 3964 2723 3981 2726
rect 2262 2713 2269 2716
rect 3348 2713 3365 2716
rect 3994 2706 3997 2725
rect 4146 2723 4172 2726
rect 4324 2723 4341 2726
rect 2250 2703 2276 2706
rect 3970 2703 3997 2706
rect 14 2667 4434 2673
rect 570 2623 573 2646
rect 116 2613 125 2616
rect 236 2613 261 2616
rect 292 2613 317 2616
rect 324 2613 333 2616
rect 428 2613 453 2616
rect 490 2613 516 2616
rect 546 2613 555 2616
rect 674 2613 685 2616
rect 314 2605 317 2613
rect 490 2593 493 2613
rect 674 2606 677 2613
rect 762 2606 765 2656
rect 810 2613 852 2616
rect 914 2613 924 2616
rect 1036 2613 1061 2616
rect 1132 2613 1141 2616
rect 1146 2607 1149 2616
rect 562 2603 588 2606
rect 661 2603 677 2606
rect 682 2603 692 2606
rect 706 2603 715 2606
rect 748 2603 757 2606
rect 762 2603 772 2606
rect 826 2603 844 2606
rect 882 2603 900 2606
rect 930 2603 948 2606
rect 980 2603 989 2606
rect 1186 2603 1189 2626
rect 1236 2613 1245 2616
rect 1338 2607 1341 2616
rect 1325 2603 1333 2606
rect 1378 2603 1381 2626
rect 1690 2616 1693 2636
rect 1386 2613 1404 2616
rect 1466 2613 1474 2616
rect 666 2593 683 2596
rect 1106 2593 1116 2596
rect 1306 2593 1315 2596
rect 1330 2593 1333 2603
rect 1386 2583 1389 2613
rect 1434 2596 1437 2613
rect 1442 2603 1466 2606
rect 1514 2603 1522 2606
rect 1594 2596 1597 2616
rect 1612 2613 1621 2616
rect 1626 2607 1629 2616
rect 1666 2606 1669 2616
rect 1685 2613 1693 2616
rect 1797 2613 1813 2616
rect 1818 2607 1821 2616
rect 1858 2613 1876 2616
rect 1890 2613 1900 2616
rect 1858 2606 1861 2613
rect 1930 2606 1933 2626
rect 2194 2616 2197 2623
rect 2234 2616 2237 2636
rect 2298 2633 2317 2636
rect 2266 2616 2269 2623
rect 1980 2613 1997 2616
rect 2036 2613 2053 2616
rect 2162 2613 2186 2616
rect 2194 2613 2210 2616
rect 2226 2613 2237 2616
rect 2242 2613 2252 2616
rect 2266 2613 2277 2616
rect 2294 2613 2301 2616
rect 2162 2607 2165 2613
rect 2226 2607 2229 2613
rect 1604 2603 1621 2606
rect 1666 2603 1674 2606
rect 1810 2603 1820 2606
rect 1852 2603 1861 2606
rect 1882 2603 1892 2606
rect 1930 2603 1956 2606
rect 1972 2603 1989 2606
rect 2098 2603 2115 2606
rect 2194 2603 2203 2606
rect 2234 2603 2243 2606
rect 1410 2593 1418 2596
rect 1434 2593 1445 2596
rect 1810 2593 1813 2603
rect 2274 2596 2277 2613
rect 2306 2606 2309 2626
rect 2314 2616 2317 2633
rect 2314 2613 2322 2616
rect 2326 2613 2340 2616
rect 2420 2613 2437 2616
rect 2362 2606 2365 2613
rect 2458 2606 2461 2625
rect 2922 2623 2925 2646
rect 3514 2633 3533 2636
rect 3130 2623 3140 2626
rect 3410 2616 3413 2626
rect 3452 2623 3469 2626
rect 2492 2613 2516 2616
rect 2594 2613 2612 2616
rect 2764 2613 2781 2616
rect 2826 2613 2844 2616
rect 2906 2613 2940 2616
rect 2978 2613 2996 2616
rect 3060 2613 3077 2616
rect 3196 2613 3205 2616
rect 3034 2606 3037 2613
rect 3202 2606 3205 2613
rect 3314 2613 3332 2616
rect 3410 2613 3436 2616
rect 3466 2613 3476 2616
rect 3500 2613 3517 2616
rect 3530 2615 3533 2633
rect 3778 2633 3797 2636
rect 4018 2633 4045 2636
rect 3660 2613 3685 2616
rect 3314 2606 3317 2613
rect 2290 2603 2314 2606
rect 2330 2603 2346 2606
rect 2362 2603 2388 2606
rect 2412 2603 2437 2606
rect 2458 2603 2468 2606
rect 2708 2603 2725 2606
rect 2850 2603 2868 2606
rect 2922 2603 2931 2606
rect 2964 2603 2997 2606
rect 3018 2603 3037 2606
rect 3170 2603 3188 2606
rect 3202 2603 3220 2606
rect 3236 2603 3261 2606
rect 3300 2603 3317 2606
rect 3322 2603 3340 2606
rect 3354 2603 3387 2606
rect 3410 2603 3428 2606
rect 3554 2603 3580 2606
rect 3596 2603 3613 2606
rect 3722 2603 3748 2606
rect 3322 2596 3325 2603
rect 3020 2593 3029 2596
rect 3060 2593 3085 2596
rect 3306 2593 3325 2596
rect 3356 2593 3373 2596
rect 3500 2593 3517 2596
rect 3778 2593 3781 2633
rect 3818 2613 3828 2616
rect 4042 2615 4045 2633
rect 4106 2613 4116 2616
rect 4154 2613 4180 2616
rect 4332 2613 4341 2616
rect 4106 2606 4109 2613
rect 4098 2603 4109 2606
rect 4114 2603 4124 2606
rect 4140 2603 4165 2606
rect 4100 2593 4109 2596
rect 38 2567 4410 2573
rect 178 2527 181 2535
rect 194 2533 204 2536
rect 346 2527 349 2535
rect 562 2533 572 2536
rect 116 2523 141 2526
rect 172 2524 181 2527
rect 188 2523 205 2526
rect 284 2523 309 2526
rect 340 2524 349 2527
rect 356 2523 365 2526
rect 514 2523 524 2526
rect 556 2523 573 2526
rect 596 2523 605 2526
rect 602 2522 605 2523
rect 610 2493 613 2556
rect 2234 2553 2245 2556
rect 1486 2543 1509 2546
rect 1818 2543 1829 2546
rect 1826 2536 1829 2543
rect 1906 2536 1909 2545
rect 2178 2543 2186 2546
rect 2234 2536 2237 2553
rect 2250 2546 2253 2556
rect 2242 2543 2253 2546
rect 2410 2545 2420 2546
rect 2410 2543 2421 2545
rect 2434 2543 2460 2546
rect 2658 2543 2676 2546
rect 2690 2543 2708 2546
rect 658 2533 675 2536
rect 708 2533 715 2536
rect 740 2533 757 2536
rect 938 2533 948 2536
rect 1138 2533 1155 2536
rect 1226 2533 1235 2536
rect 1290 2533 1315 2536
rect 1350 2533 1373 2536
rect 1404 2533 1428 2536
rect 1458 2533 1466 2536
rect 1506 2533 1516 2536
rect 1548 2533 1565 2536
rect 1690 2533 1708 2536
rect 1740 2533 1765 2536
rect 1804 2533 1821 2536
rect 1826 2533 1836 2536
rect 1884 2533 1909 2536
rect 1980 2533 1997 2536
rect 2018 2533 2027 2536
rect 2052 2533 2069 2536
rect 2074 2533 2092 2536
rect 2106 2533 2115 2536
rect 2164 2533 2196 2536
rect 2234 2533 2253 2536
rect 2378 2533 2388 2536
rect 754 2526 757 2533
rect 786 2526 789 2533
rect 1138 2526 1141 2533
rect 658 2523 683 2526
rect 754 2523 765 2526
rect 786 2523 797 2526
rect 898 2523 924 2526
rect 978 2523 1004 2526
rect 1018 2523 1029 2526
rect 1076 2523 1101 2526
rect 1132 2523 1141 2526
rect 1218 2523 1243 2526
rect 1274 2523 1284 2526
rect 1362 2523 1386 2526
rect 1410 2523 1436 2526
rect 1450 2523 1459 2526
rect 972 2513 981 2516
rect 1026 2506 1029 2523
rect 1404 2513 1413 2516
rect 1450 2513 1453 2523
rect 1506 2516 1509 2533
rect 1562 2526 1565 2533
rect 1770 2526 1773 2533
rect 1514 2523 1524 2526
rect 1562 2523 1580 2526
rect 1628 2523 1645 2526
rect 1706 2523 1716 2526
rect 1746 2523 1773 2526
rect 1810 2523 1844 2526
rect 1850 2523 1868 2526
rect 1930 2523 1956 2526
rect 1986 2523 2021 2526
rect 2140 2523 2173 2526
rect 2378 2525 2381 2533
rect 2418 2526 2421 2543
rect 2850 2536 2853 2546
rect 3188 2543 3205 2546
rect 3554 2543 3564 2546
rect 3706 2543 3724 2546
rect 4074 2536 4077 2545
rect 2442 2533 2468 2536
rect 2490 2533 2500 2536
rect 2634 2533 2644 2536
rect 2684 2533 2701 2536
rect 2706 2533 2716 2536
rect 2746 2533 2764 2536
rect 2796 2533 2813 2536
rect 2834 2533 2860 2536
rect 2914 2533 2924 2536
rect 3100 2533 3125 2536
rect 3554 2533 3572 2536
rect 3602 2533 3612 2536
rect 3636 2533 3645 2536
rect 3650 2533 3668 2536
rect 3706 2533 3732 2536
rect 3794 2533 3804 2536
rect 3860 2533 3869 2536
rect 3978 2533 3996 2536
rect 4028 2533 4045 2536
rect 4074 2533 4085 2536
rect 4140 2533 4149 2536
rect 2698 2526 2701 2533
rect 4154 2526 4157 2534
rect 1490 2513 1509 2516
rect 1026 2503 1037 2506
rect 1850 2503 1853 2523
rect 2018 2503 2021 2523
rect 2052 2513 2061 2516
rect 2234 2513 2259 2516
rect 2266 2506 2269 2524
rect 2396 2523 2421 2526
rect 2436 2523 2453 2526
rect 2476 2523 2485 2526
rect 2524 2523 2533 2526
rect 2562 2523 2572 2526
rect 2594 2523 2612 2526
rect 2634 2523 2652 2526
rect 2698 2523 2709 2526
rect 2730 2523 2772 2526
rect 2802 2523 2828 2526
rect 2850 2523 2868 2526
rect 2886 2523 2931 2526
rect 3058 2523 3076 2526
rect 3154 2523 3164 2526
rect 3348 2523 3357 2526
rect 3412 2523 3437 2526
rect 3580 2523 3589 2526
rect 3634 2523 3676 2526
rect 3746 2523 3772 2526
rect 3794 2523 3805 2526
rect 3812 2523 3821 2526
rect 3978 2523 4004 2526
rect 4106 2523 4124 2526
rect 4146 2523 4157 2526
rect 4202 2523 4205 2534
rect 4242 2523 4252 2526
rect 4364 2523 4373 2526
rect 3794 2516 3797 2523
rect 2290 2513 2308 2516
rect 3236 2513 3245 2516
rect 3636 2513 3661 2516
rect 3788 2513 3797 2516
rect 2258 2503 2269 2506
rect 2290 2503 2309 2506
rect 2834 2483 2837 2506
rect 14 2467 4434 2473
rect 1386 2453 1413 2456
rect 1626 2453 1645 2456
rect 842 2426 845 2436
rect 636 2423 645 2426
rect 730 2423 741 2426
rect 818 2423 845 2426
rect 116 2413 141 2416
rect 196 2413 205 2416
rect 178 2403 188 2406
rect 202 2405 205 2413
rect 242 2413 260 2416
rect 370 2413 396 2416
rect 426 2413 444 2416
rect 532 2413 549 2416
rect 588 2413 597 2416
rect 242 2406 245 2413
rect 426 2406 429 2413
rect 236 2403 245 2406
rect 378 2403 388 2406
rect 420 2403 429 2406
rect 594 2393 597 2413
rect 730 2406 733 2423
rect 738 2413 754 2416
rect 812 2413 821 2416
rect 826 2413 852 2416
rect 858 2413 861 2425
rect 866 2416 869 2436
rect 1418 2433 1436 2436
rect 1450 2433 1490 2436
rect 1834 2433 1868 2436
rect 1882 2433 1893 2436
rect 2258 2433 2269 2436
rect 2290 2433 2322 2436
rect 2338 2433 2373 2436
rect 884 2423 893 2426
rect 1325 2423 1333 2426
rect 866 2413 875 2416
rect 924 2413 949 2416
rect 994 2413 1018 2416
rect 1042 2413 1077 2416
rect 1212 2413 1237 2416
rect 1242 2413 1251 2416
rect 636 2403 645 2406
rect 660 2403 669 2406
rect 674 2403 692 2406
rect 724 2403 733 2406
rect 738 2403 747 2406
rect 804 2403 829 2406
rect 858 2403 868 2406
rect 938 2403 956 2406
rect 994 2403 1012 2406
rect 1042 2403 1045 2413
rect 1122 2403 1147 2406
rect 1210 2403 1243 2406
rect 1277 2403 1285 2406
rect 666 2396 669 2403
rect 738 2396 741 2403
rect 666 2393 677 2396
rect 730 2393 741 2396
rect 1330 2396 1333 2423
rect 1338 2416 1341 2426
rect 1386 2423 1418 2426
rect 1446 2423 1453 2426
rect 1466 2423 1476 2426
rect 1506 2423 1525 2426
rect 1878 2423 1885 2426
rect 1338 2413 1347 2416
rect 1382 2413 1397 2416
rect 1402 2406 1405 2416
rect 1338 2403 1354 2406
rect 1386 2403 1405 2406
rect 1330 2393 1341 2396
rect 1386 2393 1389 2403
rect 1450 2393 1453 2423
rect 1506 2396 1509 2423
rect 1685 2413 1693 2416
rect 1749 2413 1773 2416
rect 1804 2413 1821 2416
rect 1514 2403 1540 2406
rect 1556 2403 1573 2406
rect 1626 2403 1659 2406
rect 1676 2403 1685 2406
rect 1818 2405 1821 2413
rect 1890 2406 1893 2433
rect 2250 2423 2259 2426
rect 2266 2417 2269 2433
rect 2298 2423 2317 2426
rect 2346 2423 2364 2426
rect 2370 2417 2373 2433
rect 2530 2423 2541 2426
rect 1996 2413 2029 2416
rect 2100 2413 2125 2416
rect 2156 2413 2165 2416
rect 2204 2413 2213 2416
rect 2434 2413 2444 2416
rect 2466 2413 2475 2416
rect 2498 2413 2507 2416
rect 1930 2406 1933 2413
rect 2530 2406 2533 2423
rect 2930 2416 2933 2426
rect 3852 2423 3877 2426
rect 4108 2423 4133 2426
rect 2538 2413 2556 2416
rect 2562 2413 2572 2416
rect 2644 2413 2653 2416
rect 2708 2413 2749 2416
rect 2802 2413 2821 2416
rect 1890 2403 1901 2406
rect 1930 2403 1965 2406
rect 2010 2403 2027 2406
rect 2082 2403 2092 2406
rect 2098 2403 2124 2406
rect 2138 2403 2148 2406
rect 2170 2403 2196 2406
rect 2524 2403 2533 2406
rect 2538 2403 2548 2406
rect 2626 2403 2636 2406
rect 2674 2403 2684 2406
rect 2738 2403 2748 2406
rect 2780 2403 2813 2406
rect 2818 2405 2821 2413
rect 2874 2413 2885 2416
rect 2890 2413 2900 2416
rect 2924 2413 2933 2416
rect 2938 2413 2972 2416
rect 3002 2413 3036 2416
rect 3084 2413 3093 2416
rect 3180 2413 3204 2416
rect 3348 2413 3379 2416
rect 3410 2413 3443 2416
rect 3444 2413 3453 2416
rect 3570 2413 3604 2416
rect 3610 2413 3620 2416
rect 3634 2413 3660 2416
rect 3946 2413 3956 2416
rect 3970 2413 3996 2416
rect 4114 2413 4148 2416
rect 4178 2413 4213 2416
rect 2874 2406 2877 2413
rect 2852 2403 2877 2406
rect 2882 2403 2892 2406
rect 2916 2403 2925 2406
rect 2930 2403 2964 2406
rect 2996 2403 3013 2406
rect 3186 2403 3196 2406
rect 3314 2403 3340 2406
rect 3354 2403 3372 2406
rect 2170 2396 2173 2403
rect 2538 2396 2541 2403
rect 2922 2396 2925 2403
rect 1506 2393 1525 2396
rect 2074 2393 2084 2396
rect 2154 2393 2173 2396
rect 2530 2393 2541 2396
rect 2650 2393 2676 2396
rect 2922 2393 2949 2396
rect 3410 2393 3429 2396
rect 3410 2383 3429 2386
rect 3490 2383 3493 2406
rect 3570 2403 3596 2406
rect 3626 2403 3652 2406
rect 3802 2403 3828 2406
rect 3852 2403 3861 2406
rect 3866 2403 3884 2406
rect 3930 2403 3948 2406
rect 4020 2403 4053 2406
rect 4060 2403 4069 2406
rect 4074 2403 4084 2406
rect 4202 2403 4212 2406
rect 3562 2383 3589 2386
rect 38 2367 4410 2373
rect 666 2343 684 2346
rect 818 2336 821 2345
rect 1290 2343 1308 2346
rect 1386 2343 1397 2346
rect 242 2333 268 2336
rect 322 2333 348 2336
rect 514 2333 540 2336
rect 564 2333 573 2336
rect 604 2333 621 2336
rect 660 2333 669 2336
rect 692 2333 709 2336
rect 754 2333 780 2336
rect 804 2333 821 2336
rect 876 2333 893 2336
rect 1178 2333 1188 2336
rect 1220 2333 1237 2336
rect 1284 2333 1309 2336
rect 1322 2333 1347 2336
rect 1382 2333 1389 2336
rect 170 2323 188 2326
rect 194 2323 204 2326
rect 258 2323 276 2326
rect 306 2323 316 2326
rect 322 2313 325 2333
rect 706 2326 709 2333
rect 346 2323 356 2326
rect 386 2323 396 2326
rect 562 2323 588 2326
rect 610 2323 636 2326
rect 706 2323 717 2326
rect 932 2323 957 2326
rect 1044 2323 1061 2326
rect 1100 2323 1125 2326
rect 1162 2323 1195 2326
rect 1338 2323 1354 2326
rect 804 2313 813 2316
rect 1338 2283 1341 2323
rect 1394 2306 1397 2343
rect 1402 2336 1405 2356
rect 1532 2343 1541 2346
rect 1594 2343 1605 2346
rect 2874 2343 2884 2346
rect 1602 2336 1605 2343
rect 2898 2336 2901 2346
rect 1402 2333 1418 2336
rect 1482 2333 1516 2336
rect 1538 2333 1555 2336
rect 1588 2333 1597 2336
rect 1602 2333 1620 2336
rect 1685 2333 1693 2336
rect 1740 2333 1749 2336
rect 1804 2333 1813 2336
rect 1842 2333 1858 2336
rect 1892 2333 1925 2336
rect 1978 2333 1996 2336
rect 2386 2333 2396 2336
rect 2426 2333 2436 2336
rect 1442 2323 1450 2326
rect 1394 2303 1405 2306
rect 1498 2303 1501 2333
rect 1532 2323 1549 2326
rect 1690 2303 1693 2333
rect 2602 2326 2605 2336
rect 2642 2326 2645 2335
rect 2893 2333 2901 2336
rect 2906 2333 2924 2336
rect 2954 2333 2972 2336
rect 2996 2333 3013 2336
rect 3018 2333 3028 2336
rect 3052 2333 3069 2336
rect 3100 2333 3117 2336
rect 3282 2333 3300 2336
rect 3332 2333 3349 2336
rect 3354 2333 3364 2336
rect 3538 2333 3547 2336
rect 3580 2333 3589 2336
rect 3602 2333 3612 2336
rect 3836 2333 3845 2336
rect 3882 2326 3885 2335
rect 3890 2333 3908 2336
rect 4074 2333 4084 2336
rect 4132 2333 4149 2336
rect 4170 2326 4173 2335
rect 1746 2323 1779 2326
rect 1978 2323 2004 2326
rect 2100 2323 2109 2326
rect 2122 2323 2140 2326
rect 2202 2323 2220 2326
rect 2226 2323 2253 2326
rect 2404 2323 2413 2326
rect 2444 2323 2468 2326
rect 2514 2323 2524 2326
rect 2570 2323 2596 2326
rect 2602 2323 2645 2326
rect 2652 2323 2669 2326
rect 2708 2323 2733 2326
rect 2812 2323 2829 2326
rect 2868 2323 2885 2326
rect 2946 2323 2980 2326
rect 3050 2323 3084 2326
rect 3098 2323 3117 2326
rect 3156 2323 3181 2326
rect 2250 2313 2259 2316
rect 2266 2306 2269 2323
rect 2338 2313 2356 2316
rect 2362 2306 2365 2323
rect 2412 2313 2437 2316
rect 1946 2303 1964 2306
rect 2242 2303 2269 2306
rect 2354 2303 2365 2306
rect 2458 2293 2461 2323
rect 2948 2313 2957 2316
rect 2954 2303 2957 2313
rect 3226 2303 3229 2326
rect 3234 2323 3244 2326
rect 3298 2323 3308 2326
rect 3524 2323 3533 2326
rect 3586 2323 3620 2326
rect 3692 2323 3701 2326
rect 3842 2323 3868 2326
rect 3882 2323 3893 2326
rect 3898 2323 3916 2326
rect 4098 2323 4108 2326
rect 4138 2323 4173 2326
rect 4210 2323 4228 2326
rect 4258 2323 4268 2326
rect 3530 2303 3533 2323
rect 3890 2303 3893 2323
rect 14 2267 4434 2273
rect 1098 2236 1101 2246
rect 746 2233 765 2236
rect 850 2233 869 2236
rect 116 2213 141 2216
rect 172 2213 181 2216
rect 236 2213 261 2216
rect 292 2213 309 2216
rect 354 2213 372 2216
rect 428 2213 445 2216
rect 484 2213 501 2216
rect 636 2213 653 2216
rect 690 2213 707 2216
rect 762 2215 765 2233
rect 780 2223 797 2226
rect 794 2213 797 2223
rect 866 2216 869 2233
rect 1002 2233 1013 2236
rect 1098 2233 1124 2236
rect 884 2223 901 2226
rect 802 2213 812 2216
rect 354 2206 357 2213
rect 348 2203 357 2206
rect 498 2203 501 2213
rect 546 2203 572 2206
rect 586 2203 611 2206
rect 628 2203 645 2206
rect 690 2203 715 2206
rect 732 2203 741 2206
rect 786 2203 820 2206
rect 842 2203 845 2214
rect 890 2213 915 2216
rect 972 2213 981 2216
rect 586 2183 589 2203
rect 890 2183 893 2213
rect 1002 2206 1005 2233
rect 1132 2223 1157 2226
rect 1418 2216 1421 2236
rect 1818 2226 1821 2236
rect 2138 2233 2172 2236
rect 2282 2226 2285 2236
rect 1780 2223 1789 2226
rect 1804 2223 1829 2226
rect 2156 2223 2165 2226
rect 2277 2223 2285 2226
rect 2364 2223 2389 2226
rect 2404 2223 2413 2226
rect 2893 2223 2917 2226
rect 1010 2213 1028 2216
rect 1098 2213 1116 2216
rect 1196 2213 1221 2216
rect 1330 2213 1348 2216
rect 1418 2213 1445 2216
rect 1098 2206 1101 2213
rect 1330 2206 1333 2213
rect 1442 2207 1445 2213
rect 1466 2213 1485 2216
rect 1524 2213 1541 2216
rect 1634 2213 1645 2216
rect 1730 2213 1741 2216
rect 1466 2207 1469 2213
rect 898 2203 907 2206
rect 954 2197 957 2206
rect 946 2193 955 2196
rect 970 2193 973 2206
rect 978 2197 981 2206
rect 988 2203 1005 2206
rect 1052 2203 1077 2206
rect 1084 2203 1101 2206
rect 1252 2203 1261 2206
rect 1274 2203 1284 2206
rect 1316 2203 1333 2206
rect 1414 2203 1421 2206
rect 1474 2203 1500 2206
rect 1506 2203 1509 2213
rect 946 2183 949 2193
rect 1530 2183 1533 2206
rect 1594 2203 1620 2206
rect 1602 2193 1612 2196
rect 1626 2193 1629 2213
rect 1642 2207 1645 2213
rect 1724 2203 1733 2206
rect 1738 2186 1741 2213
rect 1786 2203 1789 2213
rect 1826 2207 1829 2223
rect 1874 2213 1900 2216
rect 1930 2213 1940 2216
rect 1946 2213 1980 2216
rect 2010 2213 2028 2216
rect 2186 2213 2203 2216
rect 2218 2213 2228 2216
rect 2234 2213 2243 2216
rect 2244 2213 2261 2216
rect 2306 2213 2324 2216
rect 2378 2213 2396 2216
rect 2428 2213 2445 2216
rect 2516 2213 2541 2216
rect 2572 2213 2589 2216
rect 2596 2213 2613 2216
rect 2700 2213 2725 2216
rect 2762 2213 2788 2216
rect 2834 2213 2844 2216
rect 2922 2213 2931 2216
rect 2970 2213 2988 2216
rect 3084 2213 3093 2216
rect 3098 2213 3116 2216
rect 3162 2213 3180 2216
rect 3332 2213 3357 2216
rect 3370 2213 3379 2216
rect 3516 2213 3533 2216
rect 3540 2213 3573 2216
rect 3730 2213 3748 2216
rect 3826 2213 3852 2216
rect 3882 2213 3900 2216
rect 3924 2213 3941 2216
rect 4130 2213 4148 2216
rect 4308 2213 4325 2216
rect 4364 2213 4373 2216
rect 2010 2206 2013 2213
rect 1868 2203 1885 2206
rect 2004 2203 2013 2206
rect 2162 2203 2165 2213
rect 2210 2203 2220 2206
rect 2370 2203 2388 2206
rect 2402 2203 2420 2206
rect 2586 2205 2589 2213
rect 2610 2203 2620 2206
rect 2812 2203 2821 2206
rect 1746 2193 1755 2196
rect 1738 2183 1749 2186
rect 2610 2183 2613 2203
rect 2834 2193 2837 2213
rect 2970 2206 2973 2213
rect 3162 2206 3165 2213
rect 3826 2206 3829 2213
rect 3882 2206 3885 2213
rect 2956 2203 2973 2206
rect 3098 2203 3108 2206
rect 3140 2203 3165 2206
rect 3308 2203 3317 2206
rect 3338 2203 3372 2206
rect 3562 2203 3571 2206
rect 3730 2203 3740 2206
rect 3820 2203 3829 2206
rect 3876 2203 3885 2206
rect 3906 2203 3916 2206
rect 4050 2203 4068 2206
rect 4130 2203 4140 2206
rect 3290 2193 3300 2196
rect 38 2167 4410 2173
rect 514 2153 525 2156
rect 186 2126 189 2135
rect 266 2133 276 2136
rect 442 2133 460 2136
rect 514 2133 517 2153
rect 556 2143 573 2146
rect 522 2133 540 2136
rect 116 2123 141 2126
rect 172 2123 189 2126
rect 202 2123 212 2126
rect 242 2123 260 2126
rect 274 2123 284 2126
rect 314 2123 324 2126
rect 450 2123 468 2126
rect 498 2123 508 2126
rect 570 2103 573 2143
rect 610 2133 629 2136
rect 738 2133 741 2156
rect 1882 2143 1901 2146
rect 2948 2143 2957 2146
rect 3234 2143 3252 2146
rect 3578 2136 3581 2156
rect 770 2133 781 2136
rect 866 2133 883 2136
rect 938 2133 948 2136
rect 610 2125 613 2133
rect 618 2123 636 2126
rect 714 2123 725 2126
rect 778 2125 781 2133
rect 1082 2126 1085 2135
rect 1178 2133 1195 2136
rect 1234 2133 1251 2136
rect 1402 2133 1418 2136
rect 1434 2133 1450 2136
rect 812 2123 829 2126
rect 874 2123 892 2126
rect 1004 2123 1021 2126
rect 1060 2123 1085 2126
rect 1186 2123 1204 2126
rect 1242 2123 1260 2126
rect 1428 2123 1437 2126
rect 714 2116 717 2123
rect 674 2113 684 2116
rect 708 2113 717 2116
rect 722 2113 732 2116
rect 756 2113 773 2116
rect 874 2113 877 2123
rect 1434 2113 1437 2123
rect 1474 2106 1477 2136
rect 1522 2133 1533 2136
rect 1770 2133 1786 2136
rect 1820 2133 1837 2136
rect 1860 2133 1869 2136
rect 2396 2133 2405 2136
rect 2508 2133 2525 2136
rect 2596 2133 2605 2136
rect 2610 2133 2628 2136
rect 2660 2133 2677 2136
rect 2714 2133 2740 2136
rect 1482 2113 1492 2116
rect 1498 2106 1501 2124
rect 1516 2113 1525 2116
rect 1530 2106 1533 2133
rect 2674 2126 2677 2133
rect 2762 2126 2765 2134
rect 2770 2133 2788 2136
rect 2818 2126 2821 2136
rect 2860 2133 2893 2136
rect 2946 2133 2996 2136
rect 3034 2133 3066 2136
rect 3082 2133 3101 2136
rect 3146 2133 3180 2136
rect 3332 2133 3349 2136
rect 3354 2133 3364 2136
rect 3396 2133 3429 2136
rect 3474 2133 3508 2136
rect 3570 2133 3581 2136
rect 3802 2133 3827 2136
rect 3850 2133 3861 2136
rect 2890 2126 2893 2133
rect 1578 2123 1597 2126
rect 1676 2123 1693 2126
rect 1738 2123 1748 2126
rect 1786 2123 1795 2126
rect 2002 2123 2012 2126
rect 2026 2123 2044 2126
rect 2346 2123 2356 2126
rect 2402 2123 2412 2126
rect 2434 2123 2444 2126
rect 2450 2123 2468 2126
rect 2514 2123 2548 2126
rect 2570 2123 2580 2126
rect 2602 2123 2636 2126
rect 2674 2123 2692 2126
rect 2698 2123 2708 2126
rect 2730 2123 2748 2126
rect 2762 2123 2789 2126
rect 2796 2123 2821 2126
rect 2826 2123 2836 2126
rect 2890 2123 2908 2126
rect 2914 2123 2924 2126
rect 2948 2123 2957 2126
rect 2978 2123 2981 2133
rect 3082 2125 3085 2133
rect 3228 2123 3253 2126
rect 3268 2123 3285 2126
rect 3290 2123 3308 2126
rect 3516 2123 3525 2126
rect 3572 2123 3589 2126
rect 3636 2123 3661 2126
rect 3692 2123 3701 2126
rect 3740 2123 3749 2126
rect 3802 2123 3805 2133
rect 3858 2127 3861 2133
rect 3858 2124 3876 2127
rect 3898 2126 3901 2146
rect 3946 2133 3972 2136
rect 3898 2123 3916 2126
rect 4018 2123 4044 2126
rect 4220 2123 4229 2126
rect 1474 2103 1501 2106
rect 1522 2103 1533 2106
rect 1738 2083 1741 2123
rect 2116 2113 2125 2116
rect 2164 2113 2173 2116
rect 2178 2113 2186 2116
rect 2218 2113 2236 2116
rect 2274 2113 2284 2116
rect 2122 2093 2125 2113
rect 2170 2106 2173 2113
rect 2138 2103 2156 2106
rect 2170 2103 2181 2106
rect 2186 2103 2204 2106
rect 2226 2103 2252 2106
rect 2274 2103 2277 2113
rect 2346 2103 2349 2123
rect 2570 2103 2573 2123
rect 3892 2113 3901 2116
rect 4020 2113 4037 2116
rect 14 2067 4434 2073
rect 1026 2043 1037 2046
rect 164 2013 181 2016
rect 188 2013 197 2016
rect 276 2013 301 2016
rect 332 2013 349 2016
rect 386 2013 396 2016
rect 402 2013 420 2016
rect 450 2013 460 2016
rect 618 2013 636 2016
rect 660 2013 669 2016
rect 690 2013 716 2016
rect 748 2013 757 2016
rect 762 2013 780 2016
rect 908 2013 917 2016
rect 978 2013 988 2016
rect 178 2005 181 2013
rect 1026 2006 1029 2043
rect 3170 2036 3173 2046
rect 1132 2013 1157 2016
rect 1188 2013 1197 2016
rect 338 2003 348 2006
rect 402 2003 412 2006
rect 562 2003 580 2006
rect 612 2003 629 2006
rect 682 2003 724 2006
rect 746 2003 788 2006
rect 970 2003 980 2006
rect 1012 2003 1029 2006
rect 1034 2003 1044 2006
rect 402 1983 405 2003
rect 682 1993 685 2003
rect 1194 1986 1197 2013
rect 1202 1996 1205 2026
rect 1458 2023 1477 2026
rect 2298 2016 2301 2036
rect 3170 2033 3189 2036
rect 3506 2033 3517 2036
rect 1266 2013 1292 2016
rect 1332 2013 1341 2016
rect 1394 2013 1427 2016
rect 1458 2013 1500 2016
rect 1562 2013 1588 2016
rect 1618 2013 1650 2016
rect 1756 2013 1765 2016
rect 1794 2013 1802 2016
rect 1804 2013 1829 2016
rect 1266 2006 1269 2013
rect 1626 2006 1629 2013
rect 1210 2003 1220 2006
rect 1252 2003 1269 2006
rect 1274 2003 1284 2006
rect 1458 2003 1492 2006
rect 1554 2003 1580 2006
rect 1612 2003 1629 2006
rect 1634 2003 1642 2006
rect 1826 2005 1829 2013
rect 1866 2013 1892 2016
rect 2004 2013 2013 2016
rect 2164 2013 2173 2016
rect 2298 2013 2308 2016
rect 2386 2013 2396 2016
rect 1866 2006 1869 2013
rect 2442 2006 2445 2026
rect 2978 2023 2989 2026
rect 2978 2016 2981 2023
rect 2450 2013 2460 2016
rect 2532 2013 2549 2016
rect 2644 2013 2653 2016
rect 2700 2013 2717 2016
rect 2906 2013 2931 2016
rect 2964 2013 2981 2016
rect 2986 2013 2996 2016
rect 3042 2013 3066 2016
rect 3090 2013 3093 2026
rect 3164 2013 3181 2016
rect 3186 2006 3189 2033
rect 3290 2023 3300 2026
rect 3468 2023 3501 2026
rect 3250 2013 3268 2016
rect 3354 2013 3364 2016
rect 3396 2013 3405 2016
rect 3418 2013 3452 2016
rect 3514 2015 3517 2033
rect 3604 2013 3613 2016
rect 3618 2013 3652 2016
rect 3666 2013 3684 2016
rect 3738 2013 3746 2016
rect 3818 2013 3851 2016
rect 3890 2013 3917 2016
rect 4124 2013 4133 2016
rect 4204 2013 4213 2016
rect 4250 2013 4292 2016
rect 4322 2013 4332 2016
rect 1861 2003 1869 2006
rect 1898 2003 1916 2006
rect 2284 2003 2293 2006
rect 2380 2003 2389 2006
rect 2442 2003 2453 2006
rect 2500 2003 2509 2006
rect 2524 2003 2533 2006
rect 2597 2003 2605 2006
rect 2748 2003 2781 2006
rect 2788 2003 2797 2006
rect 2914 2003 2940 2006
rect 2978 2003 3004 2006
rect 3034 2003 3060 2006
rect 3084 2003 3117 2006
rect 3124 2003 3133 2006
rect 3156 2003 3165 2006
rect 3186 2003 3202 2006
rect 3236 2003 3245 2006
rect 3284 2003 3293 2006
rect 3338 2003 3372 2006
rect 3388 2003 3413 2006
rect 3474 2003 3501 2006
rect 3538 2003 3579 2006
rect 1202 1993 1213 1996
rect 1194 1983 1205 1986
rect 2602 1983 2605 2003
rect 3090 1993 3116 1996
rect 3610 1993 3613 2013
rect 3890 2006 3893 2013
rect 3634 2003 3644 2006
rect 3730 2003 3740 2006
rect 3876 2003 3893 2006
rect 3914 1983 3917 2013
rect 3922 2003 3940 2006
rect 3972 2003 3997 2006
rect 4098 2003 4116 2006
rect 4178 2003 4196 2006
rect 4274 2003 4284 2006
rect 38 1967 4410 1973
rect 1202 1953 1213 1956
rect 732 1943 749 1946
rect 1018 1943 1036 1946
rect 178 1933 188 1936
rect 434 1933 452 1936
rect 738 1933 780 1936
rect 802 1933 844 1936
rect 906 1933 915 1936
rect 938 1933 980 1936
rect 1004 1933 1037 1936
rect 1044 1933 1085 1936
rect 178 1926 181 1933
rect 434 1926 437 1933
rect 116 1923 141 1926
rect 172 1923 181 1926
rect 196 1923 205 1926
rect 244 1923 269 1926
rect 306 1923 324 1926
rect 372 1923 397 1926
rect 428 1923 437 1926
rect 442 1923 460 1926
rect 500 1923 509 1926
rect 556 1923 581 1926
rect 612 1923 621 1926
rect 626 1923 644 1926
rect 682 1923 707 1926
rect 732 1923 741 1926
rect 804 1923 829 1926
rect 868 1923 901 1926
rect 940 1923 965 1926
rect 1132 1923 1141 1926
rect 1202 1923 1205 1953
rect 1346 1943 1365 1946
rect 1218 1933 1228 1936
rect 1260 1933 1269 1936
rect 1274 1933 1308 1936
rect 1340 1933 1357 1936
rect 1266 1926 1269 1933
rect 1210 1923 1235 1926
rect 1266 1923 1277 1926
rect 1282 1923 1309 1926
rect 1138 1916 1141 1923
rect 1004 1913 1021 1916
rect 1138 1913 1149 1916
rect 1210 1886 1213 1923
rect 1362 1913 1365 1943
rect 1706 1936 1709 1956
rect 3074 1946 3077 1956
rect 1538 1933 1555 1936
rect 1670 1933 1709 1936
rect 1404 1923 1421 1926
rect 1618 1923 1637 1926
rect 1754 1903 1757 1946
rect 2042 1943 2060 1946
rect 1762 1933 1786 1936
rect 1820 1933 1845 1936
rect 2026 1933 2068 1936
rect 2114 1935 2132 1936
rect 2114 1933 2133 1935
rect 1842 1926 1845 1933
rect 1786 1923 1795 1926
rect 1842 1923 1858 1926
rect 1964 1923 1973 1926
rect 2020 1923 2053 1926
rect 2082 1923 2092 1926
rect 2130 1923 2133 1933
rect 2186 1926 2189 1945
rect 2316 1943 2325 1946
rect 2196 1933 2213 1936
rect 2268 1933 2277 1936
rect 2282 1933 2300 1936
rect 2140 1923 2149 1926
rect 2156 1923 2189 1926
rect 2210 1926 2213 1933
rect 2346 1926 2349 1945
rect 2356 1933 2397 1936
rect 2442 1926 2445 1945
rect 3074 1943 3084 1946
rect 2452 1933 2461 1936
rect 2466 1933 2493 1936
rect 2692 1933 2709 1936
rect 2938 1933 2964 1936
rect 3066 1933 3092 1936
rect 3106 1933 3133 1936
rect 3156 1933 3181 1936
rect 2210 1923 2228 1926
rect 2316 1923 2349 1926
rect 2364 1923 2389 1926
rect 2420 1923 2445 1926
rect 2460 1923 2485 1926
rect 2490 1925 2493 1933
rect 2706 1926 2709 1933
rect 3186 1926 3189 1946
rect 3618 1943 3629 1946
rect 3228 1933 3245 1936
rect 3250 1933 3260 1936
rect 3266 1933 3277 1936
rect 3426 1933 3452 1936
rect 3548 1933 3573 1936
rect 3604 1933 3621 1936
rect 3250 1926 3253 1933
rect 2524 1923 2533 1926
rect 2580 1923 2597 1926
rect 2706 1923 2724 1926
rect 2772 1923 2781 1926
rect 3100 1923 3109 1926
rect 3114 1923 3130 1926
rect 3186 1923 3202 1926
rect 3242 1923 3253 1926
rect 3274 1893 3277 1933
rect 3372 1923 3389 1926
rect 3460 1923 3469 1926
rect 3490 1923 3524 1926
rect 3420 1913 3445 1916
rect 1202 1883 1213 1886
rect 3618 1883 3621 1933
rect 3626 1926 3629 1943
rect 3682 1933 3716 1936
rect 3730 1933 3740 1936
rect 3778 1933 3789 1936
rect 3786 1926 3789 1933
rect 3898 1926 3901 1946
rect 3940 1933 3957 1936
rect 3954 1926 3957 1933
rect 3994 1933 4004 1936
rect 4034 1933 4052 1936
rect 4146 1933 4172 1936
rect 4244 1933 4253 1936
rect 3994 1926 3997 1933
rect 4250 1926 4253 1933
rect 3626 1923 3652 1926
rect 3738 1923 3746 1926
rect 3766 1923 3781 1926
rect 3786 1923 3804 1926
rect 3898 1923 3909 1926
rect 3954 1923 3965 1926
rect 3986 1923 3997 1926
rect 4034 1923 4044 1926
rect 4076 1923 4085 1926
rect 4146 1923 4180 1926
rect 4250 1923 4276 1926
rect 4372 1923 4381 1926
rect 3778 1916 3781 1923
rect 3778 1913 3789 1916
rect 3852 1913 3869 1916
rect 3946 1893 3949 1916
rect 4378 1913 4381 1923
rect 14 1867 4434 1873
rect 90 1853 133 1856
rect 1130 1833 1149 1836
rect 1338 1823 1341 1846
rect 1634 1843 1653 1846
rect 3234 1823 3261 1826
rect 3234 1816 3237 1823
rect 170 1813 180 1816
rect 210 1813 236 1816
rect 258 1813 276 1816
rect 330 1813 340 1816
rect 370 1813 388 1816
rect 508 1813 525 1816
rect 564 1813 581 1816
rect 586 1813 612 1816
rect 658 1813 676 1816
rect 682 1813 716 1816
rect 762 1813 780 1816
rect 884 1813 917 1816
rect 1125 1813 1157 1816
rect 1212 1813 1221 1816
rect 1322 1813 1354 1816
rect 1402 1813 1418 1816
rect 1506 1813 1525 1816
rect 1628 1813 1637 1816
rect 1642 1813 1659 1816
rect 1692 1813 1709 1816
rect 1756 1813 1773 1816
rect 1812 1813 1837 1816
rect 1884 1813 1925 1816
rect 1946 1813 1964 1816
rect 2010 1813 2020 1816
rect 2148 1813 2157 1816
rect 2242 1813 2252 1816
rect 2274 1813 2292 1816
rect 2354 1813 2364 1816
rect 2564 1813 2589 1816
rect 2620 1813 2653 1816
rect 2660 1813 2693 1816
rect 2810 1813 2828 1816
rect 2914 1813 2932 1816
rect 3018 1813 3036 1816
rect 3140 1813 3149 1816
rect 3228 1813 3237 1816
rect 3242 1813 3276 1816
rect 3322 1813 3340 1816
rect 3388 1813 3413 1816
rect 3466 1813 3476 1816
rect 3572 1813 3597 1816
rect 3630 1813 3637 1816
rect 3644 1813 3677 1816
rect 3730 1813 3763 1816
rect 3802 1813 3827 1816
rect 3866 1813 3884 1816
rect 3914 1813 3931 1816
rect 370 1806 373 1813
rect 658 1806 661 1813
rect 762 1806 765 1813
rect 210 1803 228 1806
rect 242 1803 268 1806
rect 300 1803 309 1806
rect 314 1803 332 1806
rect 364 1803 373 1806
rect 394 1803 412 1806
rect 594 1803 604 1806
rect 636 1803 661 1806
rect 740 1803 765 1806
rect 898 1803 916 1806
rect 940 1803 965 1806
rect 972 1803 981 1806
rect 986 1803 1020 1806
rect 1044 1803 1061 1806
rect 1118 1803 1133 1806
rect 1146 1803 1154 1806
rect 1180 1803 1189 1806
rect 1194 1803 1204 1806
rect 210 1783 213 1803
rect 978 1796 981 1803
rect 1130 1796 1133 1803
rect 954 1793 964 1796
rect 978 1793 1013 1796
rect 1050 1793 1068 1796
rect 1130 1793 1149 1796
rect 1194 1783 1197 1803
rect 1322 1783 1325 1813
rect 1402 1806 1405 1813
rect 1506 1806 1509 1813
rect 1834 1806 1837 1813
rect 2650 1806 2653 1813
rect 2810 1806 2813 1813
rect 2914 1806 2917 1813
rect 3018 1806 3021 1813
rect 3322 1806 3325 1813
rect 1338 1803 1347 1806
rect 1380 1803 1405 1806
rect 1484 1803 1509 1806
rect 1514 1803 1524 1806
rect 1650 1803 1668 1806
rect 1685 1803 1693 1806
rect 1834 1803 1844 1806
rect 1876 1803 1893 1806
rect 1906 1803 1924 1806
rect 1948 1803 1957 1806
rect 1980 1803 1989 1806
rect 2002 1803 2012 1806
rect 2036 1803 2061 1806
rect 2114 1803 2140 1806
rect 2162 1803 2172 1806
rect 2268 1803 2277 1806
rect 2330 1803 2372 1806
rect 2442 1803 2476 1806
rect 2634 1805 2653 1806
rect 2634 1803 2652 1805
rect 2666 1803 2692 1806
rect 2730 1803 2764 1806
rect 2796 1803 2813 1806
rect 2834 1803 2860 1806
rect 2892 1803 2917 1806
rect 2954 1803 2964 1806
rect 2996 1803 3021 1806
rect 3154 1803 3173 1806
rect 3202 1803 3219 1806
rect 3220 1803 3261 1806
rect 3300 1803 3325 1806
rect 3634 1805 3637 1813
rect 3730 1806 3733 1813
rect 3866 1806 3869 1813
rect 3658 1803 3676 1806
rect 3708 1803 3733 1806
rect 3746 1803 3754 1806
rect 3802 1803 3820 1806
rect 3852 1803 3869 1806
rect 1514 1793 1517 1803
rect 2146 1793 2164 1796
rect 2492 1793 2509 1796
rect 3170 1795 3173 1803
rect 3186 1793 3210 1796
rect 3234 1793 3253 1796
rect 3250 1783 3253 1793
rect 3306 1783 3325 1786
rect 3914 1783 3917 1813
rect 3938 1793 3941 1816
rect 4044 1813 4053 1816
rect 4100 1813 4125 1816
rect 4186 1813 4196 1816
rect 4202 1813 4220 1816
rect 4250 1813 4268 1816
rect 4250 1806 4253 1813
rect 4162 1803 4172 1806
rect 4202 1803 4212 1806
rect 4244 1803 4253 1806
rect 4162 1793 4165 1803
rect 38 1767 4410 1773
rect 1034 1743 1044 1746
rect 2186 1743 2196 1746
rect 2316 1743 2325 1746
rect 2452 1743 2477 1746
rect 2474 1736 2477 1743
rect 2554 1736 2557 1746
rect 178 1733 204 1736
rect 236 1733 261 1736
rect 394 1733 420 1736
rect 498 1733 508 1736
rect 540 1733 565 1736
rect 618 1733 652 1736
rect 684 1733 709 1736
rect 850 1733 876 1736
rect 900 1733 917 1736
rect 948 1733 973 1736
rect 978 1733 988 1736
rect 1012 1733 1045 1736
rect 1052 1733 1093 1736
rect 1116 1733 1157 1736
rect 1202 1733 1244 1736
rect 1268 1733 1277 1736
rect 1468 1733 1509 1736
rect 1540 1733 1573 1736
rect 1578 1733 1588 1736
rect 1668 1733 1677 1736
rect 1738 1733 1755 1736
rect 2076 1733 2085 1736
rect 2180 1733 2189 1736
rect 2204 1733 2213 1736
rect 2236 1733 2245 1736
rect 2268 1733 2285 1736
rect 2322 1733 2356 1736
rect 2404 1733 2413 1736
rect 2418 1733 2436 1736
rect 2474 1733 2485 1736
rect 2540 1733 2557 1736
rect 2572 1733 2597 1736
rect 2634 1733 2660 1736
rect 2684 1733 2693 1736
rect 2796 1733 2813 1736
rect 2882 1733 2924 1736
rect 2954 1733 2988 1736
rect 3018 1733 3052 1736
rect 3082 1733 3085 1756
rect 3106 1736 3109 1746
rect 3106 1733 3140 1736
rect 3220 1733 3245 1736
rect 258 1726 261 1733
rect 562 1726 565 1733
rect 706 1726 709 1733
rect 116 1723 141 1726
rect 172 1723 205 1726
rect 258 1723 276 1726
rect 332 1723 349 1726
rect 418 1723 428 1726
rect 458 1723 468 1726
rect 482 1723 516 1726
rect 562 1723 588 1726
rect 604 1723 629 1726
rect 706 1723 732 1726
rect 874 1723 883 1726
rect 1090 1725 1093 1733
rect 1578 1726 1581 1733
rect 1674 1726 1677 1733
rect 2810 1726 2813 1733
rect 3250 1726 3253 1734
rect 3266 1726 3269 1756
rect 3442 1743 3452 1746
rect 3314 1733 3348 1736
rect 3364 1733 3389 1736
rect 1124 1723 1141 1726
rect 1146 1723 1171 1726
rect 1204 1723 1229 1726
rect 1290 1723 1300 1726
rect 1364 1723 1373 1726
rect 1434 1723 1443 1726
rect 1490 1723 1524 1726
rect 1554 1723 1581 1726
rect 1596 1723 1605 1726
rect 1610 1723 1620 1726
rect 1642 1723 1652 1726
rect 1674 1723 1684 1726
rect 1766 1723 1773 1726
rect 1946 1723 1956 1726
rect 2034 1723 2052 1726
rect 2084 1723 2093 1726
rect 2276 1723 2285 1726
rect 2372 1723 2389 1726
rect 2452 1723 2469 1726
rect 2508 1723 2533 1726
rect 2580 1723 2589 1726
rect 2634 1723 2668 1726
rect 2810 1723 2828 1726
rect 2906 1723 2916 1726
rect 3060 1723 3069 1726
rect 3114 1723 3130 1726
rect 3165 1723 3173 1726
rect 3186 1723 3195 1726
rect 3229 1723 3253 1726
rect 3260 1723 3269 1726
rect 3274 1723 3283 1726
rect 3314 1723 3340 1726
rect 3372 1723 3389 1726
rect 900 1713 933 1716
rect 1268 1713 1285 1716
rect 1882 1713 1900 1716
rect 2628 1713 2653 1716
rect 2906 1713 2909 1723
rect 3066 1713 3076 1716
rect 3100 1713 3109 1716
rect 3114 1713 3117 1723
rect 3442 1716 3445 1743
rect 3450 1733 3460 1736
rect 3490 1733 3508 1736
rect 3690 1733 3716 1736
rect 3746 1733 3779 1736
rect 3834 1733 3844 1736
rect 3858 1733 3868 1736
rect 3900 1733 3909 1736
rect 4076 1733 4093 1736
rect 3906 1726 3909 1733
rect 4098 1726 4101 1734
rect 4250 1727 4253 1734
rect 3474 1723 3500 1726
rect 3532 1723 3541 1726
rect 3580 1723 3589 1726
rect 3630 1723 3637 1726
rect 3698 1723 3708 1726
rect 3740 1723 3765 1726
rect 3842 1723 3851 1726
rect 3906 1723 3924 1726
rect 4028 1723 4045 1726
rect 4090 1723 4101 1726
rect 4138 1723 4148 1726
rect 4244 1724 4253 1727
rect 3378 1713 3412 1716
rect 3436 1713 3445 1716
rect 1882 1703 1916 1706
rect 14 1667 4434 1673
rect 1482 1633 1508 1636
rect 1682 1633 1725 1636
rect 3746 1633 3765 1636
rect 1364 1623 1381 1626
rect 228 1613 253 1616
rect 284 1613 309 1616
rect 330 1613 348 1616
rect 378 1613 404 1616
rect 516 1613 525 1616
rect 530 1613 572 1616
rect 618 1613 644 1616
rect 658 1613 684 1616
rect 730 1613 756 1616
rect 996 1613 1021 1616
rect 306 1605 309 1613
rect 618 1606 621 1613
rect 730 1606 733 1613
rect 1042 1606 1045 1614
rect 1076 1613 1101 1616
rect 1180 1613 1189 1616
rect 1282 1613 1292 1616
rect 1322 1613 1347 1616
rect 1434 1613 1444 1616
rect 322 1603 340 1606
rect 386 1603 396 1606
rect 596 1603 621 1606
rect 626 1603 636 1606
rect 650 1603 676 1606
rect 708 1603 733 1606
rect 898 1603 916 1606
rect 994 1603 1045 1606
rect 1242 1603 1268 1606
rect 1308 1603 1317 1606
rect 1322 1596 1325 1613
rect 1364 1603 1405 1606
rect 954 1593 980 1596
rect 1314 1593 1325 1596
rect 1386 1593 1404 1596
rect 1482 1583 1485 1633
rect 1516 1623 1549 1626
rect 1682 1623 1716 1626
rect 1618 1613 1628 1616
rect 1650 1613 1668 1616
rect 1674 1613 1709 1616
rect 1722 1615 1725 1633
rect 1754 1613 1788 1616
rect 1820 1613 1837 1616
rect 1954 1613 1964 1616
rect 2010 1613 2036 1616
rect 2170 1613 2180 1616
rect 2290 1613 2316 1616
rect 2388 1613 2397 1616
rect 2452 1613 2493 1616
rect 2170 1606 2173 1613
rect 2498 1606 2501 1614
rect 2524 1613 2557 1616
rect 2562 1613 2572 1616
rect 2668 1613 2685 1616
rect 2690 1613 2708 1616
rect 2812 1613 2829 1616
rect 2874 1613 2908 1616
rect 3028 1613 3045 1616
rect 3154 1613 3202 1616
rect 3284 1613 3293 1616
rect 3346 1613 3373 1616
rect 1530 1603 1564 1606
rect 1754 1603 1781 1606
rect 2004 1603 2013 1606
rect 2076 1603 2101 1606
rect 2148 1603 2173 1606
rect 2220 1603 2229 1606
rect 2332 1603 2349 1606
rect 2354 1603 2372 1606
rect 2402 1603 2436 1606
rect 2490 1603 2501 1606
rect 2626 1603 2660 1606
rect 2748 1603 2765 1606
rect 2924 1603 2965 1606
rect 3148 1603 3157 1606
rect 3229 1603 3245 1606
rect 2284 1593 2309 1596
rect 2452 1593 2461 1596
rect 2524 1593 2533 1596
rect 2618 1593 2652 1596
rect 2954 1593 2964 1596
rect 3346 1583 3349 1613
rect 3354 1603 3379 1606
rect 3386 1593 3389 1615
rect 3420 1613 3429 1616
rect 3476 1613 3501 1616
rect 3532 1613 3541 1616
rect 3546 1613 3571 1616
rect 3602 1606 3605 1626
rect 3634 1616 3637 1626
rect 3746 1623 3754 1626
rect 3618 1613 3626 1616
rect 3634 1613 3652 1616
rect 3682 1613 3716 1616
rect 3762 1615 3765 1633
rect 3786 1613 3812 1616
rect 4074 1613 4092 1616
rect 4140 1613 4157 1616
rect 4236 1613 4253 1616
rect 4306 1613 4316 1616
rect 4346 1613 4364 1616
rect 3602 1603 3619 1606
rect 3634 1603 3644 1606
rect 3676 1603 3685 1606
rect 3690 1593 3693 1613
rect 4346 1606 4349 1613
rect 3740 1603 3749 1606
rect 3794 1603 3804 1606
rect 4298 1603 4308 1606
rect 4340 1603 4349 1606
rect 4298 1583 4301 1603
rect 38 1567 4410 1573
rect 1130 1553 1149 1556
rect 3058 1553 3077 1556
rect 3506 1553 3533 1556
rect 3578 1553 3613 1556
rect 978 1543 1004 1546
rect 1130 1536 1133 1553
rect 1146 1543 1156 1546
rect 1818 1543 1844 1546
rect 2482 1543 2516 1546
rect 186 1526 189 1535
rect 244 1533 253 1536
rect 322 1533 348 1536
rect 386 1533 412 1536
rect 450 1533 476 1536
rect 508 1533 533 1536
rect 762 1526 765 1535
rect 930 1533 948 1536
rect 972 1533 997 1536
rect 1018 1533 1052 1536
rect 1076 1533 1101 1536
rect 1116 1533 1133 1536
rect 1138 1533 1164 1536
rect 1460 1533 1477 1536
rect 1732 1533 1749 1536
rect 1812 1533 1829 1536
rect 1834 1533 1852 1536
rect 1882 1533 1892 1536
rect 2164 1533 2173 1536
rect 2170 1526 2173 1533
rect 2442 1533 2451 1536
rect 2442 1526 2445 1533
rect 116 1523 133 1526
rect 172 1523 189 1526
rect 196 1523 205 1526
rect 274 1523 292 1526
rect 338 1523 356 1526
rect 474 1523 484 1526
rect 572 1523 581 1526
rect 692 1523 709 1526
rect 748 1523 765 1526
rect 772 1523 781 1526
rect 828 1523 853 1526
rect 884 1523 901 1526
rect 1026 1523 1060 1526
rect 1172 1523 1213 1526
rect 1218 1523 1228 1526
rect 1298 1523 1308 1526
rect 1412 1523 1421 1526
rect 1468 1523 1493 1526
rect 1740 1523 1749 1526
rect 1860 1523 1893 1526
rect 1914 1523 1941 1526
rect 2170 1523 2188 1526
rect 2364 1523 2389 1526
rect 2420 1523 2445 1526
rect 2474 1526 2477 1534
rect 2506 1533 2524 1536
rect 2636 1533 2653 1536
rect 2914 1533 2956 1536
rect 2962 1533 2997 1536
rect 2474 1523 2485 1526
rect 2490 1523 2509 1526
rect 2578 1523 2588 1526
rect 2610 1523 2620 1526
rect 2770 1523 2796 1526
rect 2842 1523 2868 1526
rect 2962 1525 2965 1533
rect 3002 1526 3005 1534
rect 3037 1533 3053 1536
rect 2986 1523 3005 1526
rect 2482 1516 2485 1523
rect 2482 1513 2493 1516
rect 3058 1506 3061 1553
rect 3116 1533 3149 1536
rect 3154 1533 3164 1536
rect 3218 1533 3236 1536
rect 3260 1533 3269 1536
rect 3332 1533 3357 1536
rect 3362 1533 3396 1536
rect 3418 1533 3453 1536
rect 3458 1533 3468 1536
rect 3514 1533 3556 1536
rect 3586 1533 3619 1536
rect 3652 1533 3669 1536
rect 3732 1533 3741 1536
rect 3762 1533 3771 1536
rect 3796 1533 3805 1536
rect 3810 1533 3827 1536
rect 3842 1533 3868 1536
rect 3914 1533 3924 1536
rect 4026 1533 4036 1536
rect 4050 1533 4059 1536
rect 4202 1533 4212 1536
rect 4244 1533 4253 1536
rect 3362 1526 3365 1533
rect 3802 1526 3805 1533
rect 3042 1503 3061 1506
rect 3074 1523 3092 1526
rect 3122 1523 3172 1526
rect 3218 1523 3244 1526
rect 3298 1523 3306 1526
rect 3340 1523 3349 1526
rect 3354 1523 3365 1526
rect 3378 1523 3387 1526
rect 3420 1523 3445 1526
rect 3466 1523 3476 1526
rect 3564 1523 3613 1526
rect 3618 1523 3626 1526
rect 3658 1523 3700 1526
rect 3770 1523 3779 1526
rect 3802 1523 3813 1526
rect 3836 1523 3869 1526
rect 3932 1523 3941 1526
rect 3978 1523 3988 1526
rect 3074 1496 3077 1523
rect 3058 1493 3077 1496
rect 3122 1493 3125 1523
rect 3346 1516 3349 1523
rect 3188 1513 3213 1516
rect 3260 1513 3301 1516
rect 3346 1513 3365 1516
rect 3442 1513 3445 1523
rect 3732 1513 3749 1516
rect 4050 1513 4053 1533
rect 4250 1526 4253 1533
rect 4250 1523 4276 1526
rect 3738 1503 3757 1506
rect 14 1467 4434 1473
rect 3330 1433 3349 1436
rect 3442 1433 3461 1436
rect 738 1416 741 1426
rect 948 1423 965 1426
rect 3346 1423 3349 1433
rect 3458 1423 3461 1433
rect 4066 1416 4069 1426
rect 116 1413 133 1416
rect 172 1413 181 1416
rect 188 1413 197 1416
rect 236 1413 261 1416
rect 292 1413 301 1416
rect 308 1413 317 1416
rect 356 1413 381 1416
rect 412 1413 421 1416
rect 468 1413 485 1416
rect 524 1413 533 1416
rect 596 1413 621 1416
rect 652 1413 661 1416
rect 668 1413 693 1416
rect 738 1413 764 1416
rect 890 1413 908 1416
rect 994 1413 1028 1416
rect 1082 1413 1109 1416
rect 1212 1413 1253 1416
rect 1404 1413 1429 1416
rect 1460 1413 1477 1416
rect 1484 1413 1509 1416
rect 1514 1413 1524 1416
rect 1570 1413 1580 1416
rect 1634 1413 1659 1416
rect 1690 1413 1724 1416
rect 1762 1413 1779 1416
rect 1810 1413 1821 1416
rect 1900 1413 1917 1416
rect 1922 1413 1932 1416
rect 1996 1413 2013 1416
rect 2130 1413 2140 1416
rect 2162 1413 2180 1416
rect 2284 1413 2309 1416
rect 2354 1413 2396 1416
rect 2442 1413 2460 1416
rect 2524 1413 2549 1416
rect 2682 1413 2700 1416
rect 2714 1413 2740 1416
rect 2818 1413 2844 1416
rect 2882 1413 2900 1416
rect 3026 1413 3036 1416
rect 3124 1413 3133 1416
rect 3156 1413 3173 1416
rect 3317 1413 3341 1416
rect 3356 1413 3405 1416
rect 3442 1413 3476 1416
rect 3482 1413 3508 1416
rect 3570 1413 3579 1416
rect 3666 1413 3676 1416
rect 3778 1413 3804 1416
rect 3834 1413 3884 1416
rect 4034 1413 4059 1416
rect 4066 1413 4084 1416
rect 4130 1413 4148 1416
rect 4178 1413 4212 1416
rect 4242 1413 4260 1416
rect 178 1405 181 1413
rect 298 1405 301 1413
rect 418 1405 421 1413
rect 530 1405 533 1413
rect 658 1405 661 1413
rect 890 1406 893 1413
rect 674 1403 692 1406
rect 738 1403 756 1406
rect 818 1403 836 1406
rect 868 1403 893 1406
rect 948 1403 965 1406
rect 980 1403 989 1406
rect 994 1403 1020 1406
rect 1044 1403 1053 1406
rect 1068 1403 1101 1406
rect 1106 1405 1109 1413
rect 1132 1403 1157 1406
rect 1164 1403 1189 1406
rect 1194 1403 1204 1406
rect 1276 1403 1285 1406
rect 1348 1403 1357 1406
rect 1474 1405 1477 1413
rect 1506 1403 1516 1406
rect 1618 1403 1652 1406
rect 1684 1403 1693 1406
rect 1698 1403 1716 1406
rect 1740 1403 1749 1406
rect 1754 1403 1772 1406
rect 1805 1403 1813 1406
rect 986 1396 989 1403
rect 1818 1396 1821 1413
rect 2442 1406 2445 1413
rect 2682 1406 2685 1413
rect 2882 1406 2885 1413
rect 3834 1406 3837 1413
rect 4242 1406 4245 1413
rect 1882 1403 1892 1406
rect 1906 1403 1924 1406
rect 1970 1403 1988 1406
rect 2090 1403 2108 1406
rect 2156 1403 2165 1406
rect 2236 1403 2245 1406
rect 2266 1403 2276 1406
rect 2370 1403 2388 1406
rect 2420 1403 2445 1406
rect 2466 1403 2500 1406
rect 2516 1403 2541 1406
rect 2602 1403 2628 1406
rect 2660 1403 2685 1406
rect 2706 1403 2732 1406
rect 2756 1403 2781 1406
rect 2794 1403 2836 1406
rect 2868 1403 2885 1406
rect 3010 1403 3044 1406
rect 3060 1403 3116 1406
rect 3170 1403 3195 1406
rect 3229 1403 3237 1406
rect 3242 1403 3260 1406
rect 3274 1403 3306 1406
rect 3322 1403 3348 1406
rect 3362 1403 3404 1406
rect 3436 1403 3453 1406
rect 3458 1403 3468 1406
rect 3532 1403 3541 1406
rect 3546 1403 3572 1406
rect 3618 1403 3636 1406
rect 3658 1403 3668 1406
rect 3700 1403 3717 1406
rect 3764 1403 3789 1406
rect 3828 1403 3837 1406
rect 3858 1403 3876 1406
rect 3908 1403 3933 1406
rect 4042 1403 4052 1406
rect 4114 1403 4140 1406
rect 4172 1403 4181 1406
rect 4236 1403 4245 1406
rect 986 1393 1013 1396
rect 1810 1393 1821 1396
rect 2258 1393 2268 1396
rect 2762 1393 2780 1396
rect 3130 1393 3140 1396
rect 3450 1393 3453 1403
rect 38 1367 4410 1373
rect 1194 1343 1204 1346
rect 1556 1343 1565 1346
rect 2402 1343 2428 1346
rect 2442 1343 2468 1346
rect 178 1333 188 1336
rect 458 1333 476 1336
rect 834 1333 852 1336
rect 884 1333 893 1336
rect 972 1333 981 1336
rect 1146 1333 1156 1336
rect 1180 1333 1189 1336
rect 178 1326 181 1333
rect 890 1326 893 1333
rect 978 1326 981 1333
rect 1194 1326 1197 1343
rect 2490 1336 2493 1356
rect 3378 1346 3381 1356
rect 2756 1343 2781 1346
rect 3130 1343 3155 1346
rect 3378 1343 3387 1346
rect 4010 1343 4020 1346
rect 1212 1333 1237 1336
rect 1276 1333 1301 1336
rect 116 1323 125 1326
rect 172 1323 181 1326
rect 196 1323 205 1326
rect 292 1323 301 1326
rect 396 1323 421 1326
rect 452 1323 461 1326
rect 514 1323 524 1326
rect 572 1323 581 1326
rect 652 1323 677 1326
rect 772 1323 789 1326
rect 828 1323 837 1326
rect 842 1323 860 1326
rect 890 1323 908 1326
rect 930 1323 948 1326
rect 978 1323 996 1326
rect 1186 1323 1197 1326
rect 1242 1323 1252 1326
rect 1298 1293 1301 1333
rect 1410 1326 1413 1335
rect 1426 1333 1460 1336
rect 1498 1333 1540 1336
rect 1618 1333 1628 1336
rect 1642 1333 1668 1336
rect 1836 1333 1853 1336
rect 1954 1333 1988 1336
rect 2020 1333 2045 1336
rect 2066 1333 2084 1336
rect 2108 1333 2117 1336
rect 1340 1323 1349 1326
rect 1396 1323 1413 1326
rect 1450 1323 1468 1326
rect 1498 1313 1501 1333
rect 2042 1326 2045 1333
rect 2322 1326 2325 1335
rect 2476 1333 2493 1336
rect 2546 1333 2564 1336
rect 2578 1333 2596 1336
rect 2650 1333 2676 1336
rect 2682 1333 2692 1336
rect 2714 1333 2740 1336
rect 2754 1333 2796 1336
rect 2828 1333 2853 1336
rect 3028 1333 3045 1336
rect 3050 1333 3060 1336
rect 3082 1333 3100 1336
rect 3124 1333 3157 1336
rect 3165 1333 3181 1336
rect 3210 1333 3220 1336
rect 1506 1323 1532 1326
rect 1578 1323 1596 1326
rect 1676 1323 1693 1326
rect 1740 1323 1765 1326
rect 1802 1323 1820 1326
rect 1892 1323 1917 1326
rect 2042 1323 2060 1326
rect 2122 1323 2140 1326
rect 2252 1323 2269 1326
rect 2308 1323 2325 1326
rect 2332 1323 2357 1326
rect 2362 1323 2372 1326
rect 2484 1323 2509 1326
rect 2514 1323 2524 1326
rect 2572 1323 2589 1326
rect 2690 1323 2700 1326
rect 2722 1323 2732 1326
rect 2754 1325 2757 1333
rect 2850 1326 2853 1333
rect 3050 1326 3053 1333
rect 2794 1323 2803 1326
rect 2850 1323 2868 1326
rect 2978 1323 3012 1326
rect 3026 1323 3053 1326
rect 3242 1326 3245 1336
rect 3274 1333 3284 1336
rect 3306 1333 3333 1336
rect 3364 1333 3381 1336
rect 3396 1333 3445 1336
rect 3842 1333 3868 1336
rect 3892 1333 3917 1336
rect 3948 1333 3973 1336
rect 3988 1333 3997 1336
rect 4028 1333 4053 1336
rect 4236 1333 4245 1336
rect 3274 1326 3277 1333
rect 3242 1323 3260 1326
rect 3261 1323 3277 1326
rect 3330 1326 3333 1333
rect 4242 1326 4245 1333
rect 3330 1323 3348 1326
rect 3410 1323 3443 1326
rect 3468 1323 3493 1326
rect 3532 1323 3541 1326
rect 3652 1323 3677 1326
rect 3708 1323 3717 1326
rect 3780 1323 3805 1326
rect 3858 1323 3876 1326
rect 3890 1323 3932 1326
rect 4180 1323 4197 1326
rect 4242 1323 4269 1326
rect 1506 1313 1509 1323
rect 2108 1313 2133 1316
rect 2540 1313 2557 1316
rect 3124 1313 3141 1316
rect 3300 1313 3325 1316
rect 3892 1313 3901 1316
rect 14 1267 4434 1273
rect 210 1253 237 1256
rect 2418 1253 2429 1256
rect 140 1213 165 1216
rect 210 1213 260 1216
rect 282 1213 316 1216
rect 354 1213 372 1216
rect 450 1213 468 1216
rect 474 1213 516 1216
rect 652 1213 669 1216
rect 716 1213 725 1216
rect 778 1213 804 1216
rect 948 1213 957 1216
rect 962 1213 979 1216
rect 354 1206 357 1213
rect 450 1206 453 1213
rect 202 1203 252 1206
rect 266 1203 308 1206
rect 340 1203 357 1206
rect 378 1203 404 1206
rect 436 1203 453 1206
rect 498 1203 508 1206
rect 580 1203 597 1206
rect 644 1203 669 1206
rect 802 1203 812 1206
rect 828 1203 837 1206
rect 842 1203 876 1206
rect 930 1203 940 1206
rect 962 1196 965 1213
rect 1004 1203 1029 1206
rect 1034 1196 1037 1226
rect 1618 1223 1637 1226
rect 1042 1213 1052 1216
rect 1090 1213 1117 1216
rect 1132 1213 1149 1216
rect 1180 1213 1221 1216
rect 1250 1213 1284 1216
rect 1316 1213 1341 1216
rect 1356 1213 1397 1216
rect 1516 1213 1541 1216
rect 1618 1213 1621 1223
rect 1634 1213 1644 1216
rect 1676 1213 1693 1216
rect 1732 1213 1757 1216
rect 1788 1213 1797 1216
rect 1804 1213 1821 1216
rect 1882 1213 1892 1216
rect 1924 1213 1949 1216
rect 1956 1213 1981 1216
rect 2100 1213 2117 1216
rect 2156 1213 2165 1216
rect 2212 1213 2237 1216
rect 2356 1213 2373 1216
rect 1042 1203 1060 1206
rect 1114 1196 1117 1213
rect 1162 1203 1172 1206
rect 1228 1203 1292 1206
rect 1322 1203 1348 1206
rect 1450 1203 1492 1206
rect 1530 1203 1540 1206
rect 1554 1203 1580 1206
rect 1642 1203 1652 1206
rect 1794 1205 1797 1213
rect 2418 1206 2421 1253
rect 3124 1223 3141 1226
rect 3170 1216 3173 1246
rect 3354 1233 3357 1256
rect 2426 1213 2436 1216
rect 2482 1213 2500 1216
rect 2588 1213 2613 1216
rect 2644 1213 2653 1216
rect 2748 1213 2780 1216
rect 2834 1213 2852 1216
rect 2882 1213 2900 1216
rect 2906 1213 2924 1216
rect 2956 1213 2973 1216
rect 3020 1213 3029 1216
rect 3076 1213 3085 1216
rect 3090 1213 3108 1216
rect 3165 1213 3173 1216
rect 3260 1213 3277 1216
rect 3316 1213 3333 1216
rect 3470 1214 3477 1217
rect 3658 1213 3676 1216
rect 3732 1213 3741 1216
rect 3748 1213 3765 1216
rect 3810 1213 3827 1216
rect 3852 1213 3869 1216
rect 3914 1213 3924 1216
rect 3954 1213 3972 1216
rect 4020 1213 4029 1216
rect 4212 1213 4221 1216
rect 2882 1206 2885 1213
rect 1818 1203 1827 1206
rect 1874 1203 1900 1206
rect 1922 1203 1948 1206
rect 1970 1203 1988 1206
rect 2034 1203 2044 1206
rect 2292 1203 2301 1206
rect 2418 1203 2429 1206
rect 2434 1203 2443 1206
rect 2460 1203 2493 1206
rect 2754 1203 2787 1206
rect 2805 1203 2821 1206
rect 2834 1203 2844 1206
rect 2876 1203 2885 1206
rect 2914 1203 2932 1206
rect 2954 1203 2973 1206
rect 3124 1203 3149 1206
rect 3156 1203 3181 1206
rect 3330 1205 3333 1213
rect 3954 1206 3957 1213
rect 3410 1203 3420 1206
rect 3482 1203 3516 1206
rect 3570 1203 3588 1206
rect 3692 1203 3717 1206
rect 3810 1203 3820 1206
rect 3858 1203 3868 1206
rect 3948 1203 3957 1206
rect 554 1193 572 1196
rect 922 1193 932 1196
rect 954 1193 965 1196
rect 1026 1193 1037 1196
rect 1818 1183 1821 1203
rect 3410 1183 3413 1203
rect 38 1167 4410 1173
rect 914 1153 933 1156
rect 602 1143 628 1146
rect 666 1136 669 1146
rect 914 1143 940 1146
rect 1004 1143 1021 1146
rect 1122 1143 1147 1146
rect 1170 1143 1180 1146
rect 1378 1143 1396 1146
rect 1476 1143 1493 1146
rect 1642 1143 1660 1146
rect 1770 1143 1780 1146
rect 1810 1136 1813 1156
rect 2106 1136 2109 1156
rect 2778 1143 2787 1146
rect 2818 1136 2821 1146
rect 3058 1136 3061 1146
rect 3186 1143 3210 1146
rect 3234 1143 3244 1146
rect 170 1133 188 1136
rect 636 1133 669 1136
rect 674 1133 684 1136
rect 706 1133 741 1136
rect 802 1133 820 1136
rect 842 1133 876 1136
rect 938 1133 948 1136
rect 1018 1133 1036 1136
rect 1042 1133 1053 1136
rect 1074 1133 1084 1136
rect 1117 1133 1149 1136
rect 1156 1133 1181 1136
rect 1188 1133 1221 1136
rect 1378 1133 1453 1136
rect 1516 1133 1525 1136
rect 1668 1133 1677 1136
rect 1690 1133 1716 1136
rect 1788 1133 1813 1136
rect 1852 1133 1877 1136
rect 1978 1133 1996 1136
rect 2028 1133 2053 1136
rect 2090 1133 2109 1136
rect 2114 1133 2124 1136
rect 2242 1133 2252 1136
rect 2346 1133 2356 1136
rect 2388 1133 2405 1136
rect 2458 1133 2492 1136
rect 2506 1133 2532 1136
rect 2634 1133 2643 1136
rect 2700 1133 2709 1136
rect 2772 1133 2789 1136
rect 2798 1133 2821 1136
rect 2978 1133 2996 1136
rect 3052 1133 3061 1136
rect 156 1123 181 1126
rect 284 1123 309 1126
rect 340 1123 365 1126
rect 410 1123 420 1126
rect 532 1123 541 1126
rect 666 1123 676 1126
rect 708 1123 725 1126
rect 738 1125 741 1133
rect 772 1123 781 1126
rect 786 1123 812 1126
rect 844 1123 853 1126
rect 914 1123 933 1126
rect 962 1123 979 1126
rect 962 1113 965 1123
rect 1018 1083 1021 1133
rect 1042 1125 1045 1133
rect 1050 1123 1092 1126
rect 1196 1123 1221 1126
rect 1316 1123 1341 1126
rect 1450 1125 1453 1133
rect 1476 1123 1501 1126
rect 1524 1123 1541 1126
rect 1580 1123 1597 1126
rect 1676 1123 1709 1126
rect 1796 1123 1813 1126
rect 1916 1123 1941 1126
rect 1986 1123 2003 1126
rect 2034 1123 2060 1126
rect 2090 1125 2093 1133
rect 2402 1126 2405 1133
rect 2706 1126 2709 1133
rect 2826 1126 2829 1133
rect 2106 1123 2132 1126
rect 2260 1123 2285 1126
rect 2290 1123 2300 1126
rect 2354 1123 2364 1126
rect 2402 1123 2420 1126
rect 2460 1123 2485 1126
rect 2500 1123 2517 1126
rect 2572 1123 2581 1126
rect 2586 1123 2603 1126
rect 2634 1123 2652 1126
rect 2706 1123 2724 1126
rect 2818 1123 2829 1126
rect 2866 1123 2876 1126
rect 2972 1123 2988 1126
rect 3020 1123 3029 1126
rect 3066 1123 3069 1135
rect 3106 1133 3130 1136
rect 3220 1133 3237 1136
rect 3242 1133 3252 1136
rect 3274 1133 3283 1136
rect 3317 1133 3341 1136
rect 3402 1133 3405 1143
rect 3410 1136 3413 1156
rect 3461 1143 3469 1146
rect 4026 1143 4044 1146
rect 3410 1133 3443 1136
rect 3836 1133 3853 1136
rect 3970 1133 3980 1136
rect 4042 1133 4052 1136
rect 4058 1133 4075 1136
rect 4090 1133 4108 1136
rect 1218 1106 1221 1123
rect 1218 1103 1237 1106
rect 2514 1103 2517 1123
rect 2578 1116 2581 1123
rect 2578 1113 2589 1116
rect 2634 1113 2637 1123
rect 3234 1113 3237 1133
rect 3274 1103 3277 1133
rect 3338 1113 3341 1133
rect 3426 1123 3436 1126
rect 3508 1123 3517 1126
rect 3732 1123 3749 1126
rect 3900 1123 3925 1126
rect 3970 1093 3973 1133
rect 3978 1123 3988 1126
rect 4116 1123 4125 1126
rect 4212 1123 4221 1126
rect 4308 1123 4317 1126
rect 14 1067 4434 1073
rect 810 1033 827 1036
rect 1650 1033 1668 1036
rect 658 1023 668 1026
rect 692 1023 709 1026
rect 812 1023 821 1026
rect 836 1023 853 1026
rect 172 1013 181 1016
rect 194 1013 204 1016
rect 234 1013 284 1016
rect 402 1013 420 1016
rect 426 1013 436 1016
rect 492 1013 501 1016
rect 548 1013 573 1016
rect 914 1013 924 1016
rect 402 1006 405 1013
rect 178 1003 196 1006
rect 308 1003 325 1006
rect 332 1003 349 1006
rect 396 1003 405 1006
rect 570 1005 573 1013
rect 604 1003 613 1006
rect 626 1003 644 1006
rect 706 1003 716 1006
rect 842 1003 868 1006
rect 954 996 957 1026
rect 1652 1023 1661 1026
rect 1010 1013 1019 1016
rect 1090 1013 1099 1016
rect 1124 1013 1149 1016
rect 1194 1013 1220 1016
rect 1308 1013 1333 1016
rect 1364 1013 1373 1016
rect 1380 1013 1405 1016
rect 1458 1013 1468 1016
rect 1492 1013 1501 1016
rect 1522 1013 1532 1016
rect 1682 1013 1708 1016
rect 1762 1013 1772 1016
rect 1826 1013 1852 1016
rect 1924 1013 1949 1016
rect 1980 1013 1997 1016
rect 2004 1013 2013 1016
rect 2018 1013 2028 1016
rect 994 1003 1011 1006
rect 1044 1003 1053 1006
rect 1066 1003 1076 1006
rect 1090 1003 1106 1006
rect 1122 1003 1156 1006
rect 1188 1003 1221 1006
rect 1370 1005 1373 1013
rect 1394 1003 1412 1006
rect 1556 1003 1581 1006
rect 1596 1003 1613 1006
rect 1834 1003 1844 1006
rect 1876 1003 1885 1006
rect 1994 1005 1997 1013
rect 2058 1006 2061 1036
rect 2706 1033 2725 1036
rect 2970 1023 2980 1026
rect 2100 1013 2125 1016
rect 2596 1013 2613 1016
rect 2652 1013 2677 1016
rect 2706 1013 2717 1016
rect 2754 1013 2772 1016
rect 2786 1013 2796 1016
rect 2058 1003 2092 1006
rect 2156 1003 2189 1006
rect 2228 1003 2245 1006
rect 2354 1003 2364 1006
rect 2396 1003 2413 1006
rect 2490 1003 2500 1006
rect 2674 1003 2692 1006
rect 314 993 324 996
rect 618 993 636 996
rect 778 993 788 996
rect 948 993 957 996
rect 1570 993 1588 996
rect 2242 993 2260 996
rect 2324 993 2341 996
rect 2354 983 2357 1003
rect 2666 993 2684 996
rect 2706 993 2709 1013
rect 2754 1006 2757 1013
rect 2866 1006 2869 1014
rect 2946 1013 2964 1016
rect 3034 1013 3044 1016
rect 3082 1013 3108 1016
rect 3138 1013 3155 1016
rect 3220 1013 3229 1016
rect 3268 1013 3293 1016
rect 2946 1006 2949 1013
rect 3306 1006 3309 1036
rect 3354 1006 3357 1036
rect 3362 1016 3365 1036
rect 3850 1033 3876 1036
rect 3834 1023 3860 1026
rect 3884 1023 3893 1026
rect 3362 1013 3387 1016
rect 3490 1013 3508 1016
rect 3514 1013 3532 1016
rect 3636 1013 3661 1016
rect 3764 1013 3789 1016
rect 3490 1006 3493 1013
rect 3946 1006 3949 1014
rect 4026 1013 4052 1016
rect 4082 1013 4116 1016
rect 4132 1013 4141 1016
rect 4146 1013 4156 1016
rect 4250 1013 4268 1016
rect 4354 1013 4372 1016
rect 4250 1006 4253 1013
rect 4354 1006 4357 1013
rect 2714 1003 2740 1006
rect 2746 1003 2757 1006
rect 2794 1003 2803 1006
rect 2834 1003 2852 1006
rect 2866 1003 2900 1006
rect 2932 1003 2949 1006
rect 3010 1003 3036 1006
rect 3082 1003 3099 1006
rect 3133 1003 3141 1006
rect 3146 1003 3157 1006
rect 3202 1003 3210 1006
rect 3274 1003 3292 1006
rect 3306 1003 3324 1006
rect 3340 1003 3357 1006
rect 3412 1003 3421 1006
rect 3426 1003 3444 1006
rect 3476 1003 3493 1006
rect 3556 1003 3573 1006
rect 3634 1003 3676 1006
rect 3746 1003 3756 1006
rect 3778 1003 3796 1006
rect 3906 1003 3924 1006
rect 3946 1003 3980 1006
rect 4012 1003 4029 1006
rect 4034 1003 4044 1006
rect 4082 1003 4108 1006
rect 4186 1003 4212 1006
rect 4244 1003 4253 1006
rect 4274 1003 4300 1006
rect 4332 1003 4357 1006
rect 2722 993 2732 996
rect 2402 983 2421 986
rect 2874 983 2877 1003
rect 3146 983 3149 1003
rect 3181 993 3197 996
rect 3268 993 3277 996
rect 3714 993 3732 996
rect 3746 993 3749 1003
rect 3194 983 3197 993
rect 38 967 4410 973
rect 586 953 605 956
rect 410 943 420 946
rect 498 943 516 946
rect 602 936 605 953
rect 1114 943 1124 946
rect 1986 936 1989 956
rect 3146 946 3149 956
rect 3146 943 3172 946
rect 3194 943 3204 946
rect 3698 943 3708 946
rect 194 933 205 936
rect 124 923 149 926
rect 194 906 197 933
rect 234 926 237 935
rect 268 933 285 936
rect 306 933 316 936
rect 362 933 372 936
rect 404 933 413 936
rect 202 923 237 926
rect 282 926 285 933
rect 282 923 324 926
rect 410 923 413 933
rect 434 933 453 936
rect 492 933 517 936
rect 524 933 541 936
rect 572 933 597 936
rect 602 933 620 936
rect 636 933 661 936
rect 700 933 717 936
rect 914 933 948 936
rect 1002 933 1011 936
rect 434 925 437 933
rect 442 923 468 926
rect 532 923 541 926
rect 650 923 676 926
rect 708 923 725 926
rect 866 923 884 926
rect 914 925 917 933
rect 922 923 956 926
rect 194 903 205 906
rect 538 893 541 923
rect 764 913 773 916
rect 714 903 756 906
rect 922 903 925 923
rect 1002 903 1005 933
rect 1370 926 1373 935
rect 1394 933 1412 936
rect 1514 933 1532 936
rect 1634 933 1660 936
rect 1682 933 1716 936
rect 1890 933 1900 936
rect 1922 926 1925 936
rect 1938 933 1948 936
rect 1986 933 1996 936
rect 2314 933 2340 936
rect 2372 933 2397 936
rect 2394 926 2397 933
rect 2450 933 2469 936
rect 2492 933 2509 936
rect 2514 933 2524 936
rect 1140 923 1157 926
rect 1194 923 1220 926
rect 1308 923 1333 926
rect 1364 923 1373 926
rect 1380 923 1405 926
rect 1410 923 1420 926
rect 1514 923 1525 926
rect 1564 923 1573 926
rect 1626 923 1652 926
rect 1684 923 1701 926
rect 1724 923 1733 926
rect 1772 923 1797 926
rect 1882 923 1892 926
rect 1956 923 1965 926
rect 1978 923 2003 926
rect 2196 923 2221 926
rect 2252 923 2277 926
rect 2394 923 2412 926
rect 1154 906 1157 923
rect 1514 916 1517 923
rect 1500 913 1517 916
rect 1834 913 1844 916
rect 1868 913 1877 916
rect 1882 913 1885 923
rect 2450 913 2453 933
rect 2506 926 2509 933
rect 2506 923 2525 926
rect 2532 923 2549 926
rect 1154 903 1173 906
rect 1458 903 1492 906
rect 1834 903 1837 913
rect 2586 896 2589 936
rect 2770 933 2787 936
rect 2820 933 2837 936
rect 2874 933 2892 936
rect 3050 933 3068 936
rect 3084 933 3109 936
rect 3140 933 3173 936
rect 3181 933 3189 936
rect 3530 933 3548 936
rect 3562 933 3580 936
rect 3716 933 3733 936
rect 3906 933 3924 936
rect 3946 933 3980 936
rect 4004 933 4021 936
rect 4210 933 4236 936
rect 2754 923 2763 926
rect 2786 923 2796 926
rect 2826 913 2844 916
rect 2850 906 2853 924
rect 2882 923 2900 926
rect 2980 923 2989 926
rect 3050 916 3053 933
rect 3092 923 3101 926
rect 3106 916 3109 933
rect 3138 923 3173 926
rect 3220 923 3245 926
rect 3284 923 3309 926
rect 3354 923 3371 926
rect 3556 923 3573 926
rect 3780 923 3805 926
rect 3948 923 3981 926
rect 4002 923 4044 926
rect 4116 923 4141 926
rect 4172 923 4181 926
rect 4188 923 4197 926
rect 4218 923 4244 926
rect 2868 913 2885 916
rect 3042 913 3053 916
rect 3098 913 3109 916
rect 2842 903 2853 906
rect 2586 893 2597 896
rect 3242 893 3245 923
rect 14 867 4434 873
rect 116 813 141 816
rect 172 813 189 816
rect 244 813 253 816
rect 292 813 317 816
rect 348 813 357 816
rect 410 813 428 816
rect 410 806 413 813
rect 178 803 196 806
rect 396 803 413 806
rect 466 806 469 846
rect 666 833 700 836
rect 714 833 748 836
rect 834 833 868 836
rect 554 823 565 826
rect 652 823 661 826
rect 674 823 684 826
rect 756 823 773 826
rect 826 823 852 826
rect 876 823 909 826
rect 1084 823 1101 826
rect 482 813 492 816
rect 562 806 565 823
rect 948 813 957 816
rect 972 813 1005 816
rect 1212 813 1221 816
rect 1316 813 1333 816
rect 1372 813 1405 816
rect 1548 813 1573 816
rect 1610 813 1636 816
rect 1658 806 1661 856
rect 1986 833 2005 836
rect 1796 823 1805 826
rect 1700 813 1717 816
rect 1844 813 1853 816
rect 1924 813 1941 816
rect 2002 815 2005 833
rect 2026 826 2029 846
rect 2482 833 2493 836
rect 2538 833 2565 836
rect 2586 833 2597 836
rect 2810 833 2821 836
rect 2020 823 2029 826
rect 2276 823 2285 826
rect 2476 823 2485 826
rect 2034 813 2052 816
rect 2090 813 2100 816
rect 2180 813 2205 816
rect 2236 813 2245 816
rect 2250 813 2260 816
rect 2362 813 2396 816
rect 2450 813 2460 816
rect 2490 806 2493 833
rect 2546 823 2556 826
rect 2562 815 2565 833
rect 2594 815 2597 833
rect 2612 823 2621 826
rect 2804 823 2813 826
rect 2660 813 2669 816
rect 2708 813 2733 816
rect 2818 806 2821 833
rect 2994 833 3020 836
rect 3274 833 3285 836
rect 3738 833 3757 836
rect 2860 813 2869 816
rect 2932 813 2941 816
rect 466 803 484 806
rect 532 803 557 806
rect 562 803 580 806
rect 652 803 677 806
rect 762 803 796 806
rect 890 803 924 806
rect 978 803 1004 806
rect 1042 803 1060 806
rect 1148 803 1173 806
rect 1394 803 1404 806
rect 1652 803 1661 806
rect 1906 803 1916 806
rect 2026 803 2044 806
rect 2068 803 2085 806
rect 2242 803 2252 806
rect 2314 803 2324 806
rect 2356 803 2381 806
rect 2490 803 2508 806
rect 2805 803 2821 806
rect 2826 803 2836 806
rect 466 783 469 803
rect 2242 793 2245 803
rect 2994 783 2997 833
rect 3004 823 3013 826
rect 3266 823 3276 826
rect 3074 806 3077 814
rect 3170 813 3196 816
rect 3226 813 3237 816
rect 3260 813 3269 816
rect 3282 815 3285 833
rect 3300 823 3309 826
rect 3404 823 3413 826
rect 3418 823 3436 826
rect 3466 823 3477 826
rect 3580 823 3589 826
rect 3410 816 3413 823
rect 3378 813 3387 816
rect 3410 813 3429 816
rect 3234 806 3237 813
rect 3034 803 3052 806
rect 3074 803 3100 806
rect 3132 803 3149 806
rect 3220 803 3229 806
rect 3234 803 3252 806
rect 3348 803 3365 806
rect 3138 793 3148 796
rect 3466 783 3469 823
rect 3474 813 3484 816
rect 3564 813 3573 816
rect 3610 813 3628 816
rect 3754 815 3757 833
rect 3658 806 3661 814
rect 3794 813 3812 816
rect 3842 813 3860 816
rect 3892 813 3901 816
rect 3924 813 3941 816
rect 4020 813 4037 816
rect 4116 813 4133 816
rect 4204 813 4213 816
rect 4364 813 4373 816
rect 3482 803 3492 806
rect 3618 803 3636 806
rect 3658 803 3692 806
rect 3858 803 3868 806
rect 3930 803 3948 806
rect 3986 803 4012 806
rect 4042 803 4052 806
rect 4090 803 4108 806
rect 4122 803 4140 806
rect 4172 803 4181 806
rect 4186 803 4196 806
rect 38 767 4410 773
rect 338 743 356 746
rect 442 743 460 746
rect 474 743 501 746
rect 1642 743 1652 746
rect 2554 743 2572 746
rect 2962 743 2980 746
rect 258 726 261 735
rect 332 733 357 736
rect 364 733 397 736
rect 172 723 189 726
rect 228 723 261 726
rect 268 723 277 726
rect 282 723 308 726
rect 442 713 445 743
rect 498 736 501 743
rect 450 713 453 736
rect 468 733 493 736
rect 498 733 516 736
rect 532 733 557 736
rect 596 733 613 736
rect 706 733 748 736
rect 764 733 797 736
rect 866 733 892 736
rect 906 733 932 736
rect 962 733 980 736
rect 1018 733 1044 736
rect 1202 733 1212 736
rect 1242 733 1252 736
rect 1290 733 1308 736
rect 1322 733 1340 736
rect 1378 733 1412 736
rect 1444 733 1461 736
rect 1482 733 1500 736
rect 1570 733 1580 736
rect 1594 733 1620 736
rect 1674 733 1692 736
rect 1706 733 1724 736
rect 1810 733 1820 736
rect 1866 733 1884 736
rect 1916 733 1933 736
rect 2220 733 2237 736
rect 2266 733 2276 736
rect 2308 733 2317 736
rect 2426 733 2436 736
rect 2506 733 2524 736
rect 2570 733 2580 736
rect 2650 733 2660 736
rect 2674 733 2684 736
rect 2698 733 2708 736
rect 1202 726 1205 733
rect 1458 726 1461 733
rect 1570 726 1573 733
rect 1930 726 1933 733
rect 2234 726 2237 733
rect 2426 726 2429 733
rect 2738 726 2741 735
rect 2772 733 2781 736
rect 2914 733 2924 736
rect 2956 733 2965 736
rect 2988 733 2997 736
rect 3100 733 3109 736
rect 3274 733 3284 736
rect 3308 733 3317 736
rect 3562 733 3572 736
rect 3700 733 3733 736
rect 3772 733 3781 736
rect 4074 733 4100 736
rect 4226 733 4244 736
rect 602 723 628 726
rect 642 723 676 726
rect 708 723 717 726
rect 722 723 740 726
rect 772 723 805 726
rect 834 723 860 726
rect 914 723 940 726
rect 1018 723 1052 726
rect 1082 723 1101 726
rect 1140 723 1157 726
rect 1196 723 1205 726
rect 1220 723 1253 726
rect 1386 723 1420 726
rect 1458 723 1476 726
rect 1538 723 1573 726
rect 1602 723 1628 726
rect 1668 723 1693 726
rect 1882 723 1892 726
rect 1930 723 1948 726
rect 1996 723 2021 726
rect 2052 723 2061 726
rect 2108 723 2125 726
rect 2164 723 2181 726
rect 2234 723 2277 726
rect 2420 723 2429 726
rect 2444 723 2468 726
rect 2498 723 2532 726
rect 2594 723 2612 726
rect 2634 723 2668 726
rect 2674 723 2692 726
rect 2716 723 2741 726
rect 2778 726 2781 733
rect 3106 726 3109 733
rect 3562 726 3565 733
rect 2778 723 2796 726
rect 2844 723 2853 726
rect 2922 723 2932 726
rect 3106 723 3124 726
rect 3172 723 3189 726
rect 3266 723 3292 726
rect 3372 723 3381 726
rect 3492 723 3517 726
rect 3548 723 3565 726
rect 3570 723 3580 726
rect 3730 723 3733 733
rect 3738 723 3756 726
rect 3802 723 3812 726
rect 3884 723 3909 726
rect 4012 723 4037 726
rect 4108 723 4117 726
rect 4252 723 4269 726
rect 4308 723 4333 726
rect 4364 723 4373 726
rect 722 716 725 723
rect 714 713 725 716
rect 908 713 933 716
rect 1524 713 1533 716
rect 2628 713 2661 716
rect 3042 713 3061 716
rect 1378 683 1405 686
rect 14 667 4434 673
rect 444 623 461 626
rect 116 613 141 616
rect 172 613 181 616
rect 194 613 204 616
rect 242 613 252 616
rect 308 613 324 616
rect 604 613 613 616
rect 676 613 693 616
rect 732 613 741 616
rect 186 603 196 606
rect 228 603 237 606
rect 276 603 285 606
rect 354 603 372 606
rect 404 603 413 606
rect 450 603 468 606
rect 546 603 580 606
rect 738 605 741 613
rect 754 606 757 626
rect 1916 623 1933 626
rect 2642 616 2645 626
rect 3220 623 3237 626
rect 3458 616 3461 636
rect 828 613 837 616
rect 884 613 909 616
rect 940 613 949 616
rect 988 613 1005 616
rect 1148 613 1173 616
rect 1188 613 1197 616
rect 1220 613 1245 616
rect 1498 613 1524 616
rect 1556 613 1565 616
rect 1578 613 1588 616
rect 1594 613 1620 616
rect 1682 613 1692 616
rect 1794 613 1804 616
rect 1882 613 1900 616
rect 1986 613 2004 616
rect 2092 613 2117 616
rect 2148 613 2165 616
rect 2172 613 2181 616
rect 2234 613 2260 616
rect 2290 613 2324 616
rect 2354 613 2372 616
rect 2404 613 2437 616
rect 2548 613 2557 616
rect 2570 613 2588 616
rect 2602 613 2628 616
rect 2642 613 2668 616
rect 2738 613 2757 616
rect 2842 613 2869 616
rect 754 603 780 606
rect 796 603 805 606
rect 810 603 820 606
rect 1098 603 1124 606
rect 1162 603 1180 606
rect 1276 603 1301 606
rect 1340 603 1349 606
rect 1388 603 1413 606
rect 1458 603 1484 606
rect 1530 603 1548 606
rect 1570 603 1580 606
rect 1644 603 1661 606
rect 1666 603 1684 606
rect 1764 603 1781 606
rect 1786 603 1796 606
rect 1858 603 1868 606
rect 1882 603 1892 606
rect 1922 603 1940 606
rect 1986 603 2012 606
rect 2028 603 2037 606
rect 2162 605 2165 613
rect 2234 606 2237 613
rect 2220 603 2237 606
rect 2284 603 2309 606
rect 2354 603 2380 606
rect 2426 603 2444 606
rect 2476 603 2501 606
rect 2506 603 2524 606
rect 2540 603 2549 606
rect 2594 603 2620 606
rect 2634 603 2660 606
rect 2724 603 2741 606
rect 1778 596 1781 603
rect 2506 596 2509 603
rect 1154 593 1172 596
rect 1186 593 1204 596
rect 1458 593 1476 596
rect 1778 593 1789 596
rect 1850 593 1860 596
rect 2418 593 2436 596
rect 2450 593 2468 596
rect 2498 593 2509 596
rect 2754 583 2757 613
rect 2828 603 2861 606
rect 2866 605 2869 613
rect 3058 613 3076 616
rect 3180 613 3197 616
rect 3212 613 3229 616
rect 3244 613 3269 616
rect 3284 613 3301 616
rect 3316 613 3341 616
rect 3354 613 3371 616
rect 3452 613 3461 616
rect 3484 613 3501 616
rect 3554 613 3572 616
rect 3658 613 3677 616
rect 3698 613 3716 616
rect 3754 613 3780 616
rect 3980 613 4005 616
rect 4036 613 4061 616
rect 4068 613 4085 616
rect 4122 613 4148 616
rect 4306 613 4324 616
rect 3058 606 3061 613
rect 3554 606 3557 613
rect 3658 606 3661 613
rect 2932 603 2957 606
rect 2980 603 2989 606
rect 3052 603 3061 606
rect 3194 603 3204 606
rect 3218 603 3236 606
rect 3250 603 3276 606
rect 3290 603 3308 606
rect 3322 603 3340 606
rect 3458 603 3476 606
rect 3482 603 3508 606
rect 3540 603 3557 606
rect 3610 603 3628 606
rect 3644 603 3661 606
rect 3666 603 3684 606
rect 3690 603 3708 606
rect 3746 603 3772 606
rect 4058 605 4061 613
rect 4122 603 4140 606
rect 4306 603 4316 606
rect 2802 593 2820 596
rect 2906 593 2924 596
rect 3458 593 3468 596
rect 3658 593 3676 596
rect 38 567 4410 573
rect 1266 553 1285 556
rect 2018 543 2036 546
rect 3306 543 3316 546
rect 202 526 205 535
rect 218 533 228 536
rect 332 533 349 536
rect 388 533 412 536
rect 436 533 445 536
rect 498 533 516 536
rect 540 533 557 536
rect 658 533 676 536
rect 940 533 957 536
rect 1052 533 1061 536
rect 1124 533 1133 536
rect 1196 533 1236 536
rect 1266 533 1292 536
rect 1316 533 1325 536
rect 1386 533 1420 536
rect 1452 533 1461 536
rect 1586 533 1604 536
rect 1700 533 1717 536
rect 1834 533 1852 536
rect 1884 533 1901 536
rect 1906 533 1924 536
rect 2004 533 2037 536
rect 2050 533 2068 536
rect 2202 533 2228 536
rect 2244 533 2277 536
rect 954 526 957 533
rect 1058 526 1061 533
rect 1458 526 1461 533
rect 1714 526 1717 533
rect 2282 526 2285 535
rect 2316 533 2333 536
rect 2370 533 2388 536
rect 124 523 149 526
rect 180 523 205 526
rect 212 523 221 526
rect 282 523 308 526
rect 434 523 468 526
rect 498 523 524 526
rect 666 523 684 526
rect 756 523 781 526
rect 812 523 829 526
rect 874 523 884 526
rect 954 523 972 526
rect 988 523 1005 526
rect 1058 523 1100 526
rect 1138 523 1172 526
rect 1210 523 1244 526
rect 1282 523 1300 526
rect 1394 523 1428 526
rect 1458 523 1476 526
rect 1524 523 1533 526
rect 1658 523 1676 526
rect 1714 523 1732 526
rect 1970 523 1988 526
rect 2052 523 2061 526
rect 2132 523 2157 526
rect 2188 523 2213 526
rect 2266 523 2285 526
rect 2330 526 2333 533
rect 2594 526 2597 535
rect 2602 533 2612 536
rect 2634 526 2637 535
rect 2642 533 2652 536
rect 2682 533 2692 536
rect 2802 533 2828 536
rect 2906 533 2932 536
rect 2970 533 2996 536
rect 3028 533 3037 536
rect 3234 533 3268 536
rect 3324 533 3333 536
rect 3338 533 3364 536
rect 3410 533 3420 536
rect 3434 533 3444 536
rect 3476 533 3508 536
rect 3532 533 3541 536
rect 3578 533 3604 536
rect 3650 533 3660 536
rect 3778 533 3796 536
rect 3826 533 3852 536
rect 3868 533 3909 536
rect 4202 533 4212 536
rect 4244 533 4253 536
rect 3034 526 3037 533
rect 4250 526 4253 533
rect 2330 523 2348 526
rect 2354 523 2364 526
rect 2386 523 2396 526
rect 2426 523 2460 526
rect 2490 523 2516 526
rect 2562 523 2580 526
rect 2594 523 2605 526
rect 2634 523 2645 526
rect 2730 523 2756 526
rect 2908 523 2925 526
rect 2978 523 3004 526
rect 3034 523 3052 526
rect 3100 523 3109 526
rect 3188 523 3197 526
rect 3242 523 3276 526
rect 3332 523 3357 526
rect 3362 523 3371 526
rect 3428 523 3452 526
rect 3546 523 3556 526
rect 3642 523 3668 526
rect 3716 523 3741 526
rect 3972 523 3981 526
rect 4076 523 4085 526
rect 4202 523 4220 526
rect 4250 523 4268 526
rect 282 513 285 523
rect 1210 483 1213 523
rect 1658 513 1661 523
rect 2602 513 2605 523
rect 3354 513 3357 523
rect 14 467 4434 473
rect 290 416 293 436
rect 124 413 149 416
rect 202 413 212 416
rect 242 413 268 416
rect 290 413 324 416
rect 354 413 372 416
rect 434 413 452 416
rect 474 413 484 416
rect 514 413 540 416
rect 596 413 621 416
rect 652 413 685 416
rect 692 413 701 416
rect 796 413 813 416
rect 852 413 877 416
rect 1036 413 1061 416
rect 1092 413 1109 416
rect 1116 413 1141 416
rect 1202 413 1220 416
rect 1268 413 1293 416
rect 1324 413 1341 416
rect 1380 413 1405 416
rect 1436 413 1461 416
rect 1484 413 1509 416
rect 1548 413 1573 416
rect 1604 413 1613 416
rect 1620 413 1653 416
rect 1818 413 1836 416
rect 1866 413 1884 416
rect 1914 413 1924 416
rect 2012 413 2021 416
rect 2124 413 2149 416
rect 2180 413 2197 416
rect 2204 413 2221 416
rect 2282 413 2300 416
rect 2546 413 2564 416
rect 2748 413 2773 416
rect 2834 413 2844 416
rect 2874 413 2892 416
rect 2906 413 2932 416
rect 2962 413 2980 416
rect 3140 413 3165 416
rect 3252 413 3277 416
rect 3308 413 3317 416
rect 3324 413 3341 416
rect 3436 413 3461 416
rect 3506 413 3524 416
rect 3554 413 3588 416
rect 3602 413 3621 416
rect 3636 413 3669 416
rect 3876 413 3909 416
rect 3946 413 3997 416
rect 4002 413 4012 416
rect 4058 413 4076 416
rect 4132 413 4149 416
rect 4186 413 4220 416
rect 4250 413 4268 416
rect 4364 413 4373 416
rect 354 406 357 413
rect 434 406 437 413
rect 514 406 517 413
rect 186 403 204 406
rect 236 403 253 406
rect 290 403 316 406
rect 348 403 357 406
rect 378 403 396 406
rect 428 403 437 406
rect 458 403 476 406
rect 508 403 517 406
rect 682 405 685 413
rect 1106 405 1109 413
rect 1122 403 1148 406
rect 1450 403 1460 406
rect 1610 405 1613 413
rect 1866 406 1869 413
rect 1684 403 1701 406
rect 1802 403 1828 406
rect 1860 403 1869 406
rect 1890 403 1916 406
rect 2194 405 2197 413
rect 2874 406 2877 413
rect 2962 406 2965 413
rect 2266 403 2292 406
rect 2324 403 2341 406
rect 2810 403 2836 406
rect 2868 403 2877 406
rect 2898 403 2924 406
rect 2956 403 2965 406
rect 3314 405 3317 413
rect 3380 403 3397 406
rect 3498 403 3516 406
rect 3554 403 3580 406
rect 3602 405 3605 413
rect 4250 406 4253 413
rect 3610 403 3628 406
rect 3634 403 3668 406
rect 3706 403 3732 406
rect 3770 403 3804 406
rect 3836 403 3853 406
rect 3868 403 3893 406
rect 3898 403 3908 406
rect 3940 403 3965 406
rect 3986 403 4004 406
rect 4042 403 4068 406
rect 4114 403 4124 406
rect 4138 403 4148 406
rect 4244 403 4253 406
rect 3898 396 3901 403
rect 3610 393 3620 396
rect 3842 393 3860 396
rect 3890 393 3901 396
rect 3946 383 3949 403
rect 38 367 4410 373
rect 2434 336 2437 346
rect 3674 336 3677 346
rect 3850 343 3860 346
rect 652 333 661 336
rect 682 333 700 336
rect 732 333 749 336
rect 874 333 892 336
rect 924 333 933 336
rect 658 326 661 333
rect 746 326 749 333
rect 930 326 933 333
rect 1082 326 1085 335
rect 1106 333 1116 336
rect 1148 333 1157 336
rect 1354 333 1372 336
rect 1402 333 1412 336
rect 1444 333 1453 336
rect 1458 333 1484 336
rect 1522 333 1556 336
rect 1586 333 1620 336
rect 1698 333 1716 336
rect 1874 333 1892 336
rect 1924 333 1941 336
rect 1938 326 1941 333
rect 2194 326 2197 335
rect 2266 333 2292 336
rect 2338 333 2356 336
rect 2388 333 2405 336
rect 2434 333 2444 336
rect 2476 333 2501 336
rect 2540 333 2557 336
rect 2692 333 2701 336
rect 2402 326 2405 333
rect 2810 327 2813 335
rect 2938 333 2956 336
rect 3226 327 3229 335
rect 3242 333 3260 336
rect 3298 333 3316 336
rect 3354 333 3371 336
rect 3404 333 3421 336
rect 3522 327 3525 335
rect 3554 333 3564 336
rect 3668 333 3677 336
rect 3682 333 3692 336
rect 3722 333 3756 336
rect 3802 333 3812 336
rect 3868 333 3885 336
rect 3890 333 3908 336
rect 3946 333 3980 336
rect 164 323 189 326
rect 292 323 317 326
rect 348 323 357 326
rect 532 323 541 326
rect 610 323 628 326
rect 658 323 676 326
rect 690 323 708 326
rect 746 323 764 326
rect 780 323 805 326
rect 850 323 893 326
rect 930 323 948 326
rect 1004 323 1029 326
rect 1060 323 1085 326
rect 1092 323 1101 326
rect 1220 323 1245 326
rect 1290 323 1324 326
rect 1380 323 1413 326
rect 1530 323 1564 326
rect 1580 323 1613 326
rect 1618 323 1628 326
rect 1692 323 1717 326
rect 1812 323 1829 326
rect 1882 323 1900 326
rect 1938 323 1956 326
rect 2124 323 2149 326
rect 2180 323 2197 326
rect 2204 323 2229 326
rect 2290 323 2300 326
rect 2346 323 2364 326
rect 2402 323 2420 326
rect 2482 323 2516 326
rect 2546 323 2572 326
rect 2588 323 2597 326
rect 2634 323 2668 326
rect 2804 324 2813 327
rect 2820 323 2829 326
rect 2994 323 3004 326
rect 3164 323 3189 326
rect 3220 324 3229 327
rect 3250 323 3268 326
rect 3306 323 3324 326
rect 3362 323 3380 326
rect 3516 324 3525 327
rect 3674 326 3677 333
rect 4298 326 4301 335
rect 4332 333 4357 336
rect 3562 323 3572 326
rect 3626 323 3644 326
rect 3674 323 3700 326
rect 3794 323 3820 326
rect 3876 323 3909 326
rect 3962 323 3988 326
rect 4250 323 4301 326
rect 4354 326 4357 333
rect 4354 323 4372 326
rect 14 267 4434 273
rect 124 213 149 216
rect 194 213 245 216
rect 540 213 557 216
rect 620 213 645 216
rect 682 213 700 216
rect 748 213 765 216
rect 810 213 836 216
rect 866 213 876 216
rect 930 213 940 216
rect 1004 213 1029 216
rect 1060 213 1069 216
rect 1082 213 1108 216
rect 1138 213 1164 216
rect 1218 213 1228 216
rect 1276 213 1301 216
rect 1346 213 1364 216
rect 1420 213 1445 216
rect 1482 213 1524 216
rect 1596 213 1621 216
rect 1682 213 1692 216
rect 1738 213 1773 216
rect 1778 213 1796 216
rect 1826 213 1852 216
rect 1938 213 1965 216
rect 2116 213 2141 216
rect 2172 213 2197 216
rect 2290 213 2300 216
rect 2492 213 2517 216
rect 2548 213 2565 216
rect 2642 213 2668 216
rect 2674 213 2684 216
rect 2700 213 2733 216
rect 2850 213 2893 216
rect 2938 213 2972 216
rect 2988 213 3029 216
rect 3074 213 3108 216
rect 3146 213 3164 216
rect 3170 213 3212 216
rect 3258 213 3293 216
rect 3338 213 3372 216
rect 3378 213 3388 216
rect 3402 213 3436 216
rect 3482 213 3517 216
rect 3628 213 3653 216
rect 3690 213 3716 216
rect 3722 213 3748 216
rect 3922 213 3948 216
rect 3954 213 3988 216
rect 4018 213 4060 216
rect 4066 213 4092 216
rect 4098 213 4116 216
rect 4122 213 4148 216
rect 4178 213 4220 216
rect 4308 213 4317 216
rect 242 205 245 213
rect 282 203 316 206
rect 370 203 388 206
rect 420 203 445 206
rect 554 205 557 213
rect 818 203 828 206
rect 1066 205 1069 213
rect 1738 206 1741 213
rect 1826 206 1829 213
rect 1938 206 1941 213
rect 1138 203 1156 206
rect 1338 203 1356 206
rect 1434 203 1444 206
rect 1490 203 1516 206
rect 1666 203 1684 206
rect 1716 203 1741 206
rect 1762 203 1788 206
rect 1820 203 1829 206
rect 1874 203 1884 206
rect 1916 203 1941 206
rect 2194 205 2197 213
rect 2252 203 2277 206
rect 2282 203 2292 206
rect 2562 205 2565 213
rect 2850 206 2853 213
rect 2938 206 2941 213
rect 3146 206 3149 213
rect 3258 206 3261 213
rect 3482 206 3485 213
rect 3922 206 3925 213
rect 4018 206 4021 213
rect 2578 203 2604 206
rect 2636 203 2653 206
rect 2706 203 2732 206
rect 2770 203 2804 206
rect 2836 203 2853 206
rect 2882 203 2892 206
rect 2924 203 2941 206
rect 2994 203 3028 206
rect 3066 203 3100 206
rect 3132 203 3149 206
rect 3178 203 3204 206
rect 3236 203 3261 206
rect 3332 203 3357 206
rect 3394 203 3428 206
rect 3460 203 3485 206
rect 3506 203 3532 206
rect 3794 203 3804 206
rect 3842 203 3876 206
rect 3908 203 3925 206
rect 3954 203 3980 206
rect 4012 203 4021 206
rect 4034 203 4052 206
rect 4074 203 4084 206
rect 4122 203 4140 206
rect 38 167 4410 173
rect 266 126 269 135
rect 1138 126 1141 135
rect 1274 126 1277 135
rect 1298 133 1308 136
rect 1466 133 1484 136
rect 1516 133 1533 136
rect 1882 133 1892 136
rect 1924 133 1941 136
rect 1530 126 1533 133
rect 1938 126 1941 133
rect 2194 126 2197 135
rect 2322 126 2325 135
rect 2458 126 2461 135
rect 2650 126 2653 135
rect 196 123 221 126
rect 252 123 269 126
rect 452 123 477 126
rect 508 123 533 126
rect 570 123 580 126
rect 620 123 629 126
rect 836 123 845 126
rect 1060 123 1085 126
rect 1116 123 1141 126
rect 1148 123 1165 126
rect 1204 123 1221 126
rect 1260 123 1277 126
rect 1284 123 1309 126
rect 1404 123 1421 126
rect 1474 123 1492 126
rect 1530 123 1548 126
rect 1874 123 1900 126
rect 1938 123 1956 126
rect 2116 123 2133 126
rect 2172 123 2197 126
rect 2204 123 2213 126
rect 2308 123 2325 126
rect 2380 123 2405 126
rect 2436 123 2461 126
rect 2468 123 2493 126
rect 2580 123 2605 126
rect 2636 123 2653 126
rect 2716 123 2741 126
rect 3036 123 3045 126
rect 3708 123 3733 126
rect 14 67 4434 73
rect 38 37 4410 57
rect 14 13 4434 33
<< metal2 >>
rect 338 4337 381 4340
rect 14 13 34 4327
rect 38 37 58 4303
rect 82 4263 117 4266
rect 66 4116 69 4216
rect 82 4203 85 4263
rect 106 4206 109 4246
rect 114 4213 117 4263
rect 170 4233 197 4236
rect 98 4203 109 4206
rect 74 4126 77 4196
rect 98 4156 101 4203
rect 98 4153 109 4156
rect 82 4133 93 4136
rect 74 4123 85 4126
rect 98 4116 101 4126
rect 66 4113 101 4116
rect 106 4106 109 4153
rect 114 4136 117 4206
rect 122 4203 125 4226
rect 170 4213 173 4233
rect 178 4213 181 4226
rect 138 4193 141 4206
rect 170 4146 173 4206
rect 154 4143 165 4146
rect 170 4143 181 4146
rect 162 4136 165 4143
rect 114 4133 141 4136
rect 66 4033 69 4106
rect 74 4103 109 4106
rect 114 4123 133 4126
rect 74 4026 77 4103
rect 66 4023 77 4026
rect 82 4023 85 4096
rect 114 4036 117 4123
rect 122 4113 133 4116
rect 122 4083 125 4106
rect 98 4033 117 4036
rect 66 3916 69 4023
rect 98 4016 101 4033
rect 106 4023 125 4026
rect 90 4013 117 4016
rect 82 3933 85 3946
rect 90 3923 93 4013
rect 106 4003 117 4006
rect 122 3956 125 4023
rect 130 3993 133 4113
rect 138 4066 141 4133
rect 146 4113 149 4126
rect 154 4106 157 4136
rect 162 4133 173 4136
rect 178 4126 181 4143
rect 186 4136 189 4226
rect 194 4213 197 4233
rect 202 4223 205 4236
rect 226 4166 229 4226
rect 242 4193 245 4206
rect 290 4176 293 4216
rect 290 4173 317 4176
rect 226 4163 269 4166
rect 194 4143 197 4156
rect 186 4133 197 4136
rect 146 4103 157 4106
rect 162 4123 181 4126
rect 194 4126 197 4133
rect 194 4123 213 4126
rect 146 4083 149 4103
rect 162 4096 165 4123
rect 218 4116 221 4136
rect 154 4093 165 4096
rect 178 4113 221 4116
rect 138 4063 145 4066
rect 142 3986 145 4063
rect 154 4013 157 4093
rect 178 4056 181 4113
rect 170 4053 181 4056
rect 170 4013 173 4053
rect 186 4033 213 4036
rect 186 4013 189 4033
rect 178 4003 197 4006
rect 178 3986 181 4003
rect 218 3996 221 4106
rect 106 3953 125 3956
rect 138 3983 145 3986
rect 170 3983 181 3986
rect 186 3993 221 3996
rect 66 3913 77 3916
rect 74 3866 77 3913
rect 66 3863 77 3866
rect 66 3843 69 3863
rect 106 3856 109 3953
rect 138 3933 141 3983
rect 90 3853 109 3856
rect 90 3806 93 3853
rect 82 3803 93 3806
rect 98 3803 101 3816
rect 106 3813 109 3846
rect 114 3803 117 3876
rect 130 3873 133 3926
rect 146 3886 149 3926
rect 170 3906 173 3983
rect 186 3913 189 3993
rect 210 3973 213 3986
rect 226 3963 229 4016
rect 170 3903 181 3906
rect 138 3883 149 3886
rect 130 3793 133 3806
rect 138 3803 141 3883
rect 178 3873 181 3903
rect 202 3873 205 3936
rect 234 3873 237 4146
rect 258 4096 261 4156
rect 266 4146 269 4163
rect 266 4143 273 4146
rect 250 4093 261 4096
rect 242 3923 245 4026
rect 250 3993 253 4093
rect 270 4086 273 4143
rect 266 4083 273 4086
rect 282 4086 285 4126
rect 314 4123 317 4173
rect 322 4133 333 4136
rect 338 4133 341 4337
rect 394 4216 397 4236
rect 386 4213 397 4216
rect 354 4156 357 4206
rect 346 4153 357 4156
rect 386 4156 389 4213
rect 402 4166 405 4216
rect 402 4163 445 4166
rect 386 4153 397 4156
rect 322 4086 325 4126
rect 282 4083 325 4086
rect 266 3943 269 4083
rect 298 4023 309 4026
rect 314 4023 317 4036
rect 322 4033 325 4046
rect 330 4023 333 4133
rect 306 4016 309 4023
rect 338 4016 341 4126
rect 346 4096 349 4153
rect 362 4133 365 4146
rect 346 4093 353 4096
rect 298 4003 301 4016
rect 306 4013 341 4016
rect 314 3966 317 4006
rect 338 3983 341 4006
rect 350 3976 353 4093
rect 394 4086 397 4153
rect 394 4083 405 4086
rect 362 4003 365 4046
rect 370 4013 373 4026
rect 386 3993 389 4006
rect 306 3963 317 3966
rect 346 3973 353 3976
rect 146 3863 181 3866
rect 146 3813 149 3863
rect 162 3786 165 3806
rect 178 3803 181 3863
rect 186 3793 189 3826
rect 194 3823 221 3826
rect 194 3813 197 3823
rect 202 3786 205 3816
rect 162 3783 205 3786
rect 242 3776 245 3806
rect 258 3803 261 3876
rect 290 3823 293 3936
rect 298 3923 301 3936
rect 306 3923 309 3963
rect 346 3896 349 3973
rect 394 3963 397 4016
rect 402 3973 405 4083
rect 410 4013 413 4126
rect 442 4123 445 4163
rect 450 4146 453 4340
rect 586 4326 589 4340
rect 578 4323 589 4326
rect 466 4203 469 4226
rect 514 4203 517 4216
rect 530 4166 533 4286
rect 526 4163 533 4166
rect 450 4143 469 4146
rect 450 4133 453 4143
rect 450 4026 453 4126
rect 474 4026 477 4136
rect 482 4123 485 4156
rect 498 4133 501 4146
rect 526 4096 529 4163
rect 514 4093 529 4096
rect 418 4013 421 4026
rect 450 4023 469 4026
rect 474 4023 509 4026
rect 466 4016 469 4023
rect 442 4013 453 4016
rect 466 4013 477 4016
rect 442 4006 445 4013
rect 426 4003 445 4006
rect 450 3993 453 4006
rect 458 3983 461 4006
rect 474 3993 477 4013
rect 370 3923 373 3936
rect 426 3923 429 3976
rect 466 3933 469 3946
rect 466 3923 477 3926
rect 338 3893 349 3896
rect 282 3776 285 3816
rect 338 3786 341 3893
rect 362 3853 405 3856
rect 362 3813 365 3853
rect 402 3813 405 3853
rect 378 3786 381 3806
rect 338 3783 381 3786
rect 242 3773 285 3776
rect 378 3753 381 3783
rect 90 3546 93 3746
rect 154 3733 157 3746
rect 290 3733 293 3746
rect 90 3543 101 3546
rect 82 3503 85 3536
rect 98 3496 101 3543
rect 114 3536 117 3616
rect 170 3546 173 3616
rect 178 3596 181 3726
rect 210 3623 213 3646
rect 234 3626 237 3726
rect 314 3636 317 3726
rect 218 3623 237 3626
rect 194 3613 213 3616
rect 186 3603 197 3606
rect 210 3596 213 3606
rect 178 3593 213 3596
rect 218 3593 221 3623
rect 242 3613 245 3626
rect 274 3613 277 3636
rect 306 3633 317 3636
rect 290 3613 293 3626
rect 154 3543 173 3546
rect 114 3533 125 3536
rect 90 3493 101 3496
rect 90 3176 93 3493
rect 114 3423 117 3526
rect 130 3463 133 3526
rect 154 3503 157 3543
rect 162 3523 165 3536
rect 178 3533 181 3586
rect 218 3543 221 3556
rect 234 3546 237 3606
rect 266 3603 277 3606
rect 306 3603 309 3633
rect 314 3623 349 3626
rect 266 3586 269 3603
rect 274 3593 285 3596
rect 266 3583 277 3586
rect 226 3543 237 3546
rect 250 3543 253 3556
rect 186 3533 205 3536
rect 226 3533 229 3543
rect 186 3526 189 3533
rect 170 3523 189 3526
rect 138 3403 141 3416
rect 162 3413 173 3416
rect 178 3403 181 3426
rect 186 3416 189 3466
rect 210 3423 213 3526
rect 234 3503 237 3536
rect 266 3533 269 3546
rect 266 3496 269 3516
rect 258 3493 269 3496
rect 258 3446 261 3493
rect 258 3443 269 3446
rect 186 3413 213 3416
rect 202 3403 213 3406
rect 218 3403 221 3416
rect 234 3413 237 3426
rect 266 3423 269 3443
rect 274 3433 277 3583
rect 282 3533 285 3593
rect 314 3583 317 3616
rect 338 3606 341 3616
rect 346 3613 349 3623
rect 354 3613 357 3626
rect 370 3613 373 3726
rect 322 3563 325 3606
rect 338 3603 349 3606
rect 402 3603 405 3746
rect 426 3686 429 3736
rect 450 3703 453 3826
rect 458 3783 461 3846
rect 466 3793 469 3836
rect 474 3803 477 3923
rect 482 3913 485 4016
rect 490 3993 493 4006
rect 498 3933 501 4016
rect 506 4003 509 4023
rect 514 4013 517 4093
rect 538 4016 541 4226
rect 554 4206 557 4256
rect 578 4246 581 4323
rect 602 4253 605 4340
rect 634 4283 637 4340
rect 706 4326 709 4340
rect 698 4323 709 4326
rect 698 4266 701 4323
rect 698 4263 709 4266
rect 578 4243 589 4246
rect 706 4243 709 4263
rect 586 4223 589 4243
rect 722 4233 725 4340
rect 746 4243 749 4340
rect 794 4326 797 4340
rect 786 4323 797 4326
rect 786 4266 789 4323
rect 786 4263 797 4266
rect 562 4213 573 4216
rect 554 4203 565 4206
rect 562 4166 565 4203
rect 578 4193 581 4216
rect 586 4196 589 4216
rect 610 4213 613 4226
rect 626 4213 645 4216
rect 594 4203 605 4206
rect 610 4196 613 4206
rect 586 4193 613 4196
rect 562 4163 573 4166
rect 546 4103 549 4126
rect 570 4086 573 4163
rect 610 4136 613 4193
rect 618 4143 621 4196
rect 626 4193 629 4206
rect 634 4136 637 4166
rect 642 4146 645 4213
rect 658 4146 661 4216
rect 682 4213 685 4226
rect 674 4203 685 4206
rect 674 4186 677 4203
rect 698 4196 701 4216
rect 682 4193 701 4196
rect 714 4186 717 4206
rect 730 4193 733 4206
rect 674 4183 701 4186
rect 714 4183 733 4186
rect 642 4143 653 4146
rect 658 4143 685 4146
rect 610 4133 645 4136
rect 650 4133 653 4143
rect 610 4123 645 4126
rect 610 4113 613 4123
rect 626 4093 629 4106
rect 554 4083 573 4086
rect 538 4013 549 4016
rect 514 4003 533 4006
rect 506 3923 509 3956
rect 514 3933 517 4003
rect 530 3856 533 3946
rect 538 3933 541 4006
rect 546 3936 549 4013
rect 554 3996 557 4083
rect 570 4013 573 4046
rect 586 4023 589 4036
rect 578 4013 589 4016
rect 578 4006 581 4013
rect 562 4003 581 4006
rect 554 3993 565 3996
rect 546 3933 557 3936
rect 522 3853 533 3856
rect 522 3823 525 3853
rect 522 3803 525 3816
rect 546 3813 549 3926
rect 554 3843 557 3933
rect 562 3906 565 3993
rect 570 3923 573 4003
rect 586 3953 589 4006
rect 594 4003 597 4026
rect 610 4003 613 4046
rect 634 4043 637 4116
rect 642 4113 645 4123
rect 658 4103 661 4136
rect 666 4133 677 4136
rect 682 4133 685 4143
rect 666 4123 677 4126
rect 690 4106 693 4146
rect 698 4123 701 4183
rect 706 4123 725 4126
rect 706 4113 709 4123
rect 690 4103 717 4106
rect 722 4103 725 4116
rect 730 4103 733 4183
rect 738 4113 741 4126
rect 714 4096 717 4103
rect 746 4096 749 4136
rect 714 4093 749 4096
rect 658 4013 669 4016
rect 578 3916 581 3936
rect 586 3933 597 3936
rect 626 3933 629 3956
rect 642 3933 645 3986
rect 674 3936 677 4006
rect 682 3953 685 4026
rect 690 4023 693 4036
rect 698 4026 701 4036
rect 698 4023 709 4026
rect 698 3963 701 4016
rect 674 3933 685 3936
rect 578 3913 613 3916
rect 562 3903 569 3906
rect 566 3826 569 3903
rect 666 3856 669 3926
rect 562 3823 569 3826
rect 634 3853 669 3856
rect 562 3803 565 3823
rect 634 3813 637 3853
rect 554 3733 557 3756
rect 426 3683 453 3686
rect 450 3656 453 3683
rect 442 3653 453 3656
rect 338 3593 349 3596
rect 338 3553 341 3593
rect 282 3516 285 3526
rect 298 3523 301 3546
rect 306 3516 309 3526
rect 282 3513 309 3516
rect 322 3446 325 3536
rect 346 3533 349 3586
rect 426 3583 429 3616
rect 442 3606 445 3653
rect 506 3636 509 3726
rect 602 3723 605 3796
rect 634 3723 637 3806
rect 650 3733 653 3846
rect 682 3836 685 3933
rect 706 3926 709 4023
rect 714 4013 717 4093
rect 754 4086 757 4196
rect 762 4123 765 4156
rect 770 4126 773 4216
rect 778 4133 781 4166
rect 770 4123 781 4126
rect 746 4083 757 4086
rect 746 3983 749 4083
rect 770 3993 773 4016
rect 778 3963 781 4116
rect 786 3956 789 4136
rect 794 3966 797 4263
rect 802 4126 805 4246
rect 810 4213 813 4340
rect 826 4326 829 4340
rect 826 4323 837 4326
rect 834 4256 837 4323
rect 882 4256 885 4340
rect 1018 4256 1021 4340
rect 834 4253 853 4256
rect 882 4253 897 4256
rect 1018 4253 1053 4256
rect 810 4133 813 4156
rect 826 4143 829 4216
rect 850 4196 853 4253
rect 842 4193 853 4196
rect 802 4123 813 4126
rect 802 4093 805 4116
rect 810 4056 813 4123
rect 826 4106 829 4126
rect 818 4103 829 4106
rect 810 4053 817 4056
rect 814 4006 817 4053
rect 810 4003 817 4006
rect 810 3973 813 4003
rect 826 3993 829 4016
rect 834 4013 837 4136
rect 842 4126 845 4193
rect 874 4183 877 4216
rect 894 4186 897 4253
rect 906 4193 909 4216
rect 922 4203 925 4216
rect 894 4183 901 4186
rect 850 4133 869 4136
rect 842 4123 849 4126
rect 794 3963 801 3966
rect 778 3953 789 3956
rect 730 3933 733 3946
rect 746 3943 765 3946
rect 762 3936 765 3943
rect 762 3933 773 3936
rect 778 3933 781 3953
rect 706 3923 725 3926
rect 762 3903 765 3926
rect 770 3886 773 3933
rect 786 3923 789 3946
rect 674 3833 685 3836
rect 762 3883 773 3886
rect 762 3836 765 3883
rect 762 3833 773 3836
rect 674 3813 677 3833
rect 698 3776 701 3816
rect 730 3793 733 3816
rect 770 3813 773 3833
rect 778 3803 781 3906
rect 798 3896 801 3963
rect 818 3933 821 3986
rect 834 3963 837 4006
rect 846 3966 849 4123
rect 858 4076 861 4126
rect 866 4093 869 4133
rect 858 4073 869 4076
rect 846 3963 853 3966
rect 842 3923 845 3946
rect 850 3933 853 3963
rect 858 3926 861 4066
rect 866 4013 869 4073
rect 874 4023 877 4116
rect 882 4003 885 4156
rect 890 4123 893 4146
rect 898 4036 901 4183
rect 922 4133 925 4186
rect 954 4126 957 4216
rect 970 4146 973 4216
rect 962 4133 965 4146
rect 970 4143 997 4146
rect 1002 4143 1005 4216
rect 1018 4203 1021 4216
rect 1050 4196 1053 4253
rect 1066 4203 1069 4216
rect 1098 4213 1101 4340
rect 1186 4326 1189 4340
rect 1178 4323 1189 4326
rect 1178 4266 1181 4323
rect 1202 4276 1205 4340
rect 1282 4326 1285 4340
rect 1194 4273 1205 4276
rect 1274 4323 1285 4326
rect 1178 4263 1185 4266
rect 1114 4203 1117 4216
rect 994 4133 997 4143
rect 906 4123 941 4126
rect 954 4123 965 4126
rect 922 4086 925 4116
rect 930 4103 933 4116
rect 938 4113 957 4116
rect 938 4086 941 4113
rect 962 4106 965 4123
rect 922 4083 941 4086
rect 946 4036 949 4106
rect 890 4033 901 4036
rect 938 4033 949 4036
rect 954 4103 965 4106
rect 890 3996 893 4033
rect 898 4013 909 4016
rect 898 4003 909 4006
rect 938 4003 941 4033
rect 954 4003 957 4103
rect 978 4023 981 4126
rect 1002 4103 1005 4136
rect 1018 4133 1021 4196
rect 1042 4193 1053 4196
rect 1010 4123 1021 4126
rect 1026 4113 1029 4126
rect 1042 4086 1045 4193
rect 1058 4113 1061 4136
rect 1022 4083 1045 4086
rect 1066 4106 1069 4146
rect 1082 4123 1085 4156
rect 1114 4146 1117 4196
rect 1090 4143 1117 4146
rect 1090 4116 1093 4143
rect 1082 4113 1093 4116
rect 1066 4103 1077 4106
rect 978 4003 981 4016
rect 890 3993 901 3996
rect 850 3923 861 3926
rect 798 3893 805 3896
rect 786 3793 789 3816
rect 802 3786 805 3893
rect 850 3813 853 3923
rect 786 3783 805 3786
rect 698 3773 709 3776
rect 682 3733 701 3736
rect 698 3706 701 3726
rect 706 3723 709 3773
rect 738 3706 741 3736
rect 786 3723 789 3783
rect 866 3753 869 3806
rect 498 3633 509 3636
rect 442 3603 453 3606
rect 450 3576 453 3603
rect 450 3573 461 3576
rect 354 3533 437 3536
rect 458 3533 461 3573
rect 330 3523 349 3526
rect 322 3443 333 3446
rect 258 3413 269 3416
rect 258 3406 261 3413
rect 242 3403 261 3406
rect 146 3303 149 3346
rect 194 3323 197 3346
rect 226 3323 229 3356
rect 266 3343 269 3406
rect 274 3363 277 3406
rect 290 3346 293 3436
rect 330 3413 333 3443
rect 338 3413 341 3506
rect 354 3503 357 3516
rect 370 3513 373 3526
rect 386 3523 397 3526
rect 402 3523 421 3526
rect 402 3516 405 3523
rect 394 3513 405 3516
rect 402 3493 405 3506
rect 410 3503 413 3516
rect 434 3506 437 3533
rect 434 3503 461 3506
rect 378 3393 381 3406
rect 402 3396 405 3416
rect 458 3413 461 3503
rect 482 3493 485 3616
rect 498 3553 501 3633
rect 538 3613 541 3706
rect 698 3703 741 3706
rect 698 3656 701 3703
rect 698 3653 705 3656
rect 514 3566 517 3606
rect 506 3563 517 3566
rect 506 3476 509 3563
rect 578 3533 581 3586
rect 530 3523 541 3526
rect 602 3523 605 3596
rect 498 3473 509 3476
rect 402 3393 413 3396
rect 354 3353 381 3356
rect 290 3343 297 3346
rect 266 3303 269 3336
rect 294 3296 297 3343
rect 290 3293 297 3296
rect 90 3173 101 3176
rect 98 3133 101 3173
rect 130 3166 133 3246
rect 138 3213 141 3226
rect 126 3163 133 3166
rect 126 3046 129 3163
rect 126 3043 133 3046
rect 82 3003 85 3016
rect 114 2846 117 2866
rect 114 2843 121 2846
rect 90 2766 93 2806
rect 118 2796 121 2843
rect 82 2763 93 2766
rect 114 2793 121 2796
rect 66 1896 69 2686
rect 82 2636 85 2763
rect 114 2756 117 2793
rect 110 2753 117 2756
rect 110 2656 113 2753
rect 122 2723 125 2746
rect 110 2653 117 2656
rect 74 2633 85 2636
rect 74 2436 77 2633
rect 90 2553 93 2606
rect 90 2533 93 2546
rect 74 2433 85 2436
rect 90 2413 93 2526
rect 90 2393 93 2406
rect 74 2346 77 2366
rect 74 2343 81 2346
rect 78 2266 81 2343
rect 74 2263 81 2266
rect 74 2123 77 2263
rect 90 2053 93 2386
rect 106 2306 109 2376
rect 114 2363 117 2653
rect 122 2613 125 2716
rect 130 2676 133 3043
rect 138 3013 141 3156
rect 170 3136 173 3216
rect 186 3213 189 3226
rect 210 3223 253 3226
rect 210 3203 213 3223
rect 226 3153 229 3216
rect 162 3133 173 3136
rect 146 3113 149 3126
rect 162 3086 165 3133
rect 146 3083 165 3086
rect 146 2993 149 3083
rect 178 3036 181 3126
rect 186 3113 189 3126
rect 154 3033 181 3036
rect 154 3003 157 3033
rect 162 3013 165 3026
rect 186 3013 189 3026
rect 210 2946 213 3136
rect 218 3113 221 3136
rect 242 3133 245 3216
rect 250 3213 253 3223
rect 258 3133 261 3206
rect 266 3203 269 3216
rect 290 3206 293 3293
rect 306 3213 309 3326
rect 354 3303 357 3353
rect 378 3333 381 3353
rect 410 3346 413 3393
rect 402 3343 413 3346
rect 362 3306 365 3326
rect 402 3323 405 3343
rect 498 3333 501 3473
rect 618 3446 621 3616
rect 658 3613 661 3626
rect 702 3606 705 3653
rect 834 3623 837 3726
rect 850 3723 853 3736
rect 898 3723 901 3993
rect 938 3933 941 3986
rect 1022 3976 1025 4083
rect 1066 4046 1069 4103
rect 1058 4043 1077 4046
rect 1034 4013 1037 4036
rect 1042 4013 1045 4026
rect 1058 4003 1061 4043
rect 1074 4033 1077 4043
rect 1082 4023 1085 4113
rect 1090 4016 1093 4036
rect 1082 4013 1093 4016
rect 1098 3986 1101 4116
rect 1106 4033 1109 4136
rect 1114 4056 1117 4143
rect 1122 4103 1125 4136
rect 1130 4123 1133 4146
rect 1138 4123 1141 4206
rect 1146 4106 1149 4136
rect 1162 4123 1165 4216
rect 1182 4206 1185 4263
rect 1194 4213 1197 4273
rect 1274 4266 1277 4323
rect 1274 4263 1285 4266
rect 1282 4216 1285 4263
rect 1298 4256 1301 4340
rect 1338 4266 1341 4340
rect 1338 4263 1345 4266
rect 1298 4253 1333 4256
rect 1182 4203 1189 4206
rect 1210 4203 1213 4216
rect 1154 4113 1165 4116
rect 1170 4106 1173 4136
rect 1186 4126 1189 4203
rect 1234 4146 1237 4216
rect 1218 4143 1237 4146
rect 1186 4123 1197 4126
rect 1146 4103 1173 4106
rect 1186 4103 1189 4116
rect 1114 4053 1149 4056
rect 1106 3993 1109 4026
rect 1138 4003 1141 4016
rect 1146 4013 1149 4053
rect 1018 3973 1025 3976
rect 1066 3983 1101 3986
rect 914 3753 917 3816
rect 962 3786 965 3936
rect 986 3886 989 3926
rect 1018 3923 1021 3973
rect 1026 3933 1029 3956
rect 1066 3933 1069 3983
rect 1026 3886 1029 3926
rect 986 3883 1029 3886
rect 954 3783 965 3786
rect 954 3733 957 3783
rect 994 3763 997 3876
rect 1042 3793 1045 3816
rect 1074 3813 1077 3976
rect 1106 3933 1109 3986
rect 1154 3923 1157 4016
rect 1162 4003 1165 4103
rect 1178 4013 1181 4026
rect 1178 3953 1181 4006
rect 1194 3923 1197 4123
rect 1202 4106 1205 4136
rect 1218 4123 1221 4143
rect 1210 4113 1221 4116
rect 1226 4106 1229 4136
rect 1258 4133 1261 4216
rect 1282 4213 1293 4216
rect 1306 4203 1309 4216
rect 1330 4186 1333 4253
rect 1326 4183 1333 4186
rect 1202 4103 1229 4106
rect 1226 4036 1229 4103
rect 1234 4086 1237 4126
rect 1242 4103 1245 4116
rect 1282 4086 1285 4126
rect 1326 4086 1329 4183
rect 1342 4176 1345 4263
rect 1338 4173 1345 4176
rect 1338 4123 1341 4173
rect 1346 4106 1349 4156
rect 1354 4146 1357 4216
rect 1386 4213 1389 4340
rect 1450 4326 1453 4340
rect 1442 4323 1453 4326
rect 1442 4246 1445 4323
rect 1466 4256 1469 4340
rect 1482 4326 1485 4340
rect 1482 4323 1493 4326
rect 1466 4253 1473 4256
rect 1442 4243 1453 4246
rect 1402 4203 1405 4216
rect 1442 4213 1445 4226
rect 1450 4176 1453 4243
rect 1354 4143 1397 4146
rect 1234 4083 1285 4086
rect 1314 4083 1329 4086
rect 1342 4103 1349 4106
rect 1210 4013 1213 4036
rect 1226 4033 1277 4036
rect 1226 4013 1229 4026
rect 1218 3933 1221 3986
rect 1234 3953 1237 4006
rect 1242 3993 1245 4033
rect 1258 4013 1261 4026
rect 1274 4013 1277 4033
rect 1282 4006 1285 4016
rect 1266 4003 1285 4006
rect 1298 4006 1301 4036
rect 1306 4013 1309 4026
rect 1298 4003 1309 4006
rect 1266 3923 1269 4003
rect 1274 3993 1285 3996
rect 1314 3923 1317 4083
rect 1342 4036 1345 4103
rect 1354 4083 1357 4126
rect 1370 4123 1373 4136
rect 1342 4033 1349 4036
rect 1322 4013 1325 4026
rect 1346 4003 1349 4033
rect 1354 3936 1357 4036
rect 1362 4003 1365 4016
rect 1370 4013 1373 4116
rect 1378 4113 1381 4136
rect 1394 4133 1397 4143
rect 1402 4133 1405 4146
rect 1386 4023 1389 4126
rect 1410 4116 1413 4176
rect 1450 4173 1461 4176
rect 1402 4113 1413 4116
rect 1402 4036 1405 4113
rect 1418 4046 1421 4146
rect 1458 4136 1461 4173
rect 1470 4166 1473 4253
rect 1490 4246 1493 4323
rect 1482 4243 1493 4246
rect 1482 4213 1485 4243
rect 1514 4226 1517 4340
rect 1570 4326 1573 4340
rect 1562 4323 1573 4326
rect 1490 4203 1493 4226
rect 1498 4223 1517 4226
rect 1530 4226 1533 4276
rect 1562 4266 1565 4323
rect 1562 4263 1573 4266
rect 1570 4243 1573 4263
rect 1586 4226 1589 4340
rect 1530 4223 1541 4226
rect 1578 4223 1589 4226
rect 1466 4163 1473 4166
rect 1482 4193 1493 4196
rect 1482 4163 1485 4193
rect 1498 4186 1501 4223
rect 1490 4183 1501 4186
rect 1466 4143 1469 4163
rect 1442 4133 1461 4136
rect 1474 4133 1485 4136
rect 1426 4113 1429 4126
rect 1434 4073 1437 4126
rect 1442 4056 1445 4133
rect 1450 4063 1453 4116
rect 1458 4113 1461 4126
rect 1466 4123 1477 4126
rect 1466 4093 1469 4123
rect 1482 4093 1485 4116
rect 1482 4066 1485 4086
rect 1478 4063 1485 4066
rect 1442 4053 1461 4056
rect 1418 4043 1425 4046
rect 1402 4033 1413 4036
rect 1410 4013 1413 4033
rect 1338 3933 1357 3936
rect 1362 3933 1365 3986
rect 1386 3933 1389 3946
rect 1322 3923 1349 3926
rect 1354 3873 1357 3933
rect 1422 3916 1425 4043
rect 1458 3976 1461 4053
rect 1478 3986 1481 4063
rect 1490 4053 1493 4183
rect 1506 4176 1509 4216
rect 1522 4213 1533 4216
rect 1514 4203 1525 4206
rect 1506 4173 1517 4176
rect 1498 4143 1509 4146
rect 1498 4073 1501 4143
rect 1514 4133 1517 4173
rect 1514 4063 1517 4126
rect 1522 4113 1525 4136
rect 1530 4133 1533 4213
rect 1538 4163 1541 4206
rect 1554 4193 1557 4206
rect 1578 4176 1581 4223
rect 1562 4173 1581 4176
rect 1538 4103 1541 4126
rect 1546 4106 1549 4136
rect 1554 4123 1557 4146
rect 1562 4106 1565 4173
rect 1578 4143 1581 4156
rect 1578 4126 1581 4136
rect 1586 4133 1589 4216
rect 1594 4136 1597 4246
rect 1634 4213 1637 4340
rect 1706 4326 1709 4334
rect 1682 4323 1709 4326
rect 1594 4133 1605 4136
rect 1570 4113 1573 4126
rect 1578 4123 1597 4126
rect 1546 4103 1581 4106
rect 1538 4036 1541 4056
rect 1534 4033 1541 4036
rect 1478 3983 1485 3986
rect 1458 3973 1469 3976
rect 1434 3923 1437 3936
rect 1466 3923 1469 3973
rect 1422 3913 1429 3916
rect 634 3583 637 3606
rect 698 3603 705 3606
rect 698 3583 701 3603
rect 674 3513 677 3526
rect 690 3486 693 3556
rect 714 3543 717 3616
rect 762 3553 765 3606
rect 810 3603 813 3616
rect 866 3576 869 3616
rect 858 3573 869 3576
rect 842 3546 845 3556
rect 810 3543 845 3546
rect 738 3523 741 3536
rect 810 3533 813 3543
rect 826 3533 837 3536
rect 842 3526 845 3543
rect 690 3483 717 3486
rect 818 3483 821 3526
rect 834 3523 845 3526
rect 858 3523 861 3573
rect 874 3533 877 3606
rect 898 3563 901 3716
rect 938 3593 941 3726
rect 970 3646 973 3736
rect 994 3733 997 3756
rect 970 3643 977 3646
rect 946 3603 949 3616
rect 922 3553 957 3556
rect 922 3543 925 3553
rect 898 3533 925 3536
rect 618 3443 645 3446
rect 522 3413 525 3426
rect 586 3403 589 3416
rect 602 3393 605 3406
rect 362 3303 381 3306
rect 290 3203 297 3206
rect 282 3133 285 3196
rect 294 3146 297 3203
rect 306 3196 309 3206
rect 354 3203 357 3216
rect 362 3196 365 3216
rect 306 3193 365 3196
rect 290 3143 297 3146
rect 234 3023 237 3126
rect 250 3113 253 3126
rect 266 3103 269 3126
rect 290 3013 293 3143
rect 298 3083 301 3126
rect 338 3116 341 3186
rect 370 3183 373 3206
rect 226 2993 229 3006
rect 306 2996 309 3106
rect 314 3096 317 3116
rect 338 3113 357 3116
rect 314 3093 325 3096
rect 322 3046 325 3093
rect 378 3076 381 3303
rect 410 3213 413 3326
rect 394 3133 397 3206
rect 410 3196 413 3206
rect 450 3203 453 3216
rect 458 3196 461 3216
rect 410 3193 461 3196
rect 402 3103 405 3126
rect 434 3116 437 3186
rect 466 3183 469 3226
rect 474 3203 477 3326
rect 522 3323 525 3366
rect 594 3323 597 3386
rect 642 3336 645 3443
rect 650 3413 653 3446
rect 610 3256 613 3336
rect 642 3333 653 3336
rect 698 3333 701 3416
rect 714 3376 717 3483
rect 762 3393 765 3416
rect 714 3373 733 3376
rect 602 3253 613 3256
rect 514 3203 517 3216
rect 538 3213 541 3246
rect 482 3133 485 3156
rect 490 3123 493 3166
rect 418 3083 421 3116
rect 434 3113 461 3116
rect 506 3103 509 3116
rect 378 3073 421 3076
rect 314 3043 325 3046
rect 314 3023 317 3043
rect 314 3013 341 3016
rect 410 3013 413 3036
rect 314 3003 317 3013
rect 322 3003 349 3006
rect 306 2993 317 2996
rect 410 2993 413 3006
rect 418 2983 421 3073
rect 426 2996 429 3006
rect 442 3003 445 3016
rect 450 2996 453 3006
rect 426 2993 453 2996
rect 514 2983 517 3006
rect 522 2993 525 3206
rect 546 3113 549 3216
rect 562 3196 565 3216
rect 570 3203 573 3226
rect 578 3196 581 3206
rect 562 3193 581 3196
rect 586 3156 589 3216
rect 602 3196 605 3253
rect 634 3246 637 3326
rect 650 3266 653 3333
rect 618 3243 637 3246
rect 642 3263 653 3266
rect 618 3213 621 3243
rect 626 3213 629 3236
rect 642 3233 645 3263
rect 690 3236 693 3326
rect 730 3313 733 3373
rect 834 3363 837 3523
rect 842 3503 845 3516
rect 874 3513 877 3526
rect 914 3516 917 3526
rect 882 3513 917 3516
rect 922 3496 925 3533
rect 914 3493 925 3496
rect 842 3413 845 3426
rect 874 3423 909 3426
rect 882 3406 885 3416
rect 906 3413 909 3423
rect 914 3406 917 3493
rect 930 3473 933 3546
rect 858 3393 861 3406
rect 866 3346 869 3406
rect 882 3403 917 3406
rect 882 3366 885 3386
rect 906 3373 909 3396
rect 882 3363 889 3366
rect 866 3343 877 3346
rect 682 3233 693 3236
rect 642 3223 677 3226
rect 642 3206 645 3223
rect 666 3213 669 3223
rect 674 3206 677 3216
rect 618 3203 645 3206
rect 650 3203 677 3206
rect 602 3193 613 3196
rect 610 3176 613 3193
rect 610 3173 621 3176
rect 682 3156 685 3233
rect 690 3223 725 3226
rect 690 3203 693 3223
rect 698 3203 701 3216
rect 706 3213 725 3216
rect 562 3153 589 3156
rect 658 3153 685 3156
rect 562 3143 565 3153
rect 602 3136 605 3146
rect 578 3133 605 3136
rect 658 3133 661 3153
rect 690 3133 693 3176
rect 562 3123 597 3126
rect 530 2983 533 3006
rect 538 2986 541 3006
rect 554 2993 557 3016
rect 562 2986 565 3123
rect 674 3026 677 3126
rect 722 3123 725 3206
rect 730 3163 733 3206
rect 770 3203 773 3326
rect 778 3286 781 3326
rect 802 3323 813 3326
rect 778 3283 837 3286
rect 794 3203 797 3226
rect 802 3223 829 3226
rect 802 3213 805 3223
rect 810 3203 813 3216
rect 818 3213 829 3216
rect 770 3123 773 3166
rect 818 3136 821 3213
rect 834 3203 837 3283
rect 850 3193 853 3336
rect 874 3233 877 3343
rect 886 3226 889 3363
rect 914 3343 917 3403
rect 898 3286 901 3326
rect 922 3293 925 3416
rect 938 3396 941 3553
rect 954 3543 957 3553
rect 946 3533 957 3536
rect 962 3523 965 3636
rect 974 3566 977 3643
rect 994 3636 997 3716
rect 1034 3713 1037 3736
rect 1082 3646 1085 3726
rect 1082 3643 1109 3646
rect 986 3633 997 3636
rect 986 3613 989 3633
rect 994 3623 1013 3626
rect 1018 3623 1021 3636
rect 1042 3633 1101 3636
rect 994 3613 997 3623
rect 1010 3616 1013 3623
rect 970 3563 977 3566
rect 946 3413 949 3506
rect 938 3393 949 3396
rect 954 3393 957 3446
rect 962 3403 965 3416
rect 946 3373 949 3393
rect 970 3353 973 3563
rect 986 3553 989 3606
rect 1002 3596 1005 3616
rect 1010 3613 1021 3616
rect 1026 3613 1037 3616
rect 1010 3603 1021 3606
rect 1026 3596 1029 3613
rect 1002 3593 1029 3596
rect 1026 3533 1029 3576
rect 1042 3523 1045 3633
rect 1058 3526 1061 3616
rect 1074 3586 1077 3626
rect 1098 3613 1101 3633
rect 1106 3613 1109 3643
rect 1114 3636 1117 3726
rect 1122 3723 1125 3826
rect 1130 3823 1157 3826
rect 1130 3813 1133 3823
rect 1138 3763 1141 3816
rect 1154 3793 1157 3806
rect 1162 3783 1165 3806
rect 1194 3793 1197 3866
rect 1226 3823 1229 3836
rect 1274 3833 1317 3836
rect 1130 3696 1133 3736
rect 1162 3733 1165 3746
rect 1194 3726 1197 3746
rect 1130 3693 1141 3696
rect 1138 3646 1141 3693
rect 1162 3686 1165 3726
rect 1190 3723 1197 3726
rect 1162 3683 1173 3686
rect 1138 3643 1149 3646
rect 1114 3633 1141 3636
rect 1122 3603 1125 3626
rect 1074 3583 1085 3586
rect 1066 3533 1069 3556
rect 1082 3543 1085 3583
rect 1058 3523 1069 3526
rect 1042 3503 1045 3516
rect 1050 3513 1061 3516
rect 978 3383 981 3416
rect 986 3403 989 3486
rect 1002 3386 1005 3456
rect 1050 3443 1053 3513
rect 1066 3453 1069 3523
rect 1090 3483 1093 3586
rect 1130 3576 1133 3606
rect 1114 3573 1133 3576
rect 1098 3513 1101 3546
rect 1074 3433 1077 3446
rect 1050 3423 1061 3426
rect 1050 3413 1053 3423
rect 1066 3406 1069 3416
rect 1082 3413 1085 3426
rect 1050 3403 1061 3406
rect 1066 3403 1093 3406
rect 1098 3403 1101 3426
rect 1002 3383 1029 3386
rect 930 3343 1005 3346
rect 930 3323 933 3343
rect 938 3286 941 3326
rect 954 3316 957 3336
rect 970 3333 973 3343
rect 986 3333 997 3336
rect 1002 3333 1005 3343
rect 970 3323 981 3326
rect 986 3316 989 3326
rect 954 3313 989 3316
rect 898 3283 941 3286
rect 994 3273 997 3333
rect 1010 3323 1013 3346
rect 1018 3236 1021 3356
rect 1026 3323 1029 3383
rect 986 3233 1021 3236
rect 858 3186 861 3206
rect 866 3196 869 3226
rect 882 3223 889 3226
rect 962 3223 1005 3226
rect 874 3203 877 3216
rect 866 3193 877 3196
rect 882 3186 885 3223
rect 890 3186 893 3206
rect 858 3183 893 3186
rect 794 3133 821 3136
rect 826 3123 829 3146
rect 874 3133 877 3156
rect 618 3003 621 3026
rect 634 3013 637 3026
rect 674 3023 701 3026
rect 538 2983 565 2986
rect 186 2933 189 2946
rect 210 2943 221 2946
rect 218 2896 221 2943
rect 234 2903 237 2926
rect 210 2893 221 2896
rect 186 2856 189 2886
rect 210 2863 213 2893
rect 178 2853 189 2856
rect 138 2813 141 2826
rect 178 2796 181 2853
rect 202 2803 205 2846
rect 178 2793 189 2796
rect 130 2673 137 2676
rect 134 2606 137 2673
rect 162 2646 165 2666
rect 130 2603 137 2606
rect 158 2643 165 2646
rect 106 2303 117 2306
rect 82 1956 85 2006
rect 106 2003 109 2016
rect 114 1976 117 2303
rect 122 2226 125 2506
rect 130 2243 133 2603
rect 158 2586 161 2643
rect 170 2613 173 2736
rect 178 2716 181 2726
rect 186 2723 189 2793
rect 194 2716 197 2736
rect 178 2713 197 2716
rect 202 2703 205 2726
rect 186 2636 189 2656
rect 210 2636 213 2806
rect 218 2753 221 2816
rect 226 2803 229 2826
rect 234 2823 261 2826
rect 234 2813 237 2823
rect 234 2803 245 2806
rect 250 2793 253 2816
rect 258 2776 261 2823
rect 234 2773 261 2776
rect 218 2663 221 2726
rect 226 2713 229 2736
rect 182 2633 189 2636
rect 194 2633 213 2636
rect 158 2583 165 2586
rect 162 2566 165 2583
rect 162 2563 173 2566
rect 138 2523 141 2546
rect 154 2536 157 2556
rect 154 2533 161 2536
rect 158 2486 161 2533
rect 154 2483 161 2486
rect 138 2413 141 2426
rect 138 2336 141 2356
rect 138 2333 145 2336
rect 142 2266 145 2333
rect 154 2293 157 2483
rect 170 2456 173 2563
rect 182 2526 185 2633
rect 194 2533 197 2633
rect 210 2603 213 2626
rect 234 2596 237 2773
rect 242 2733 245 2766
rect 250 2626 253 2756
rect 258 2733 261 2766
rect 266 2656 269 2946
rect 330 2933 333 2946
rect 298 2886 301 2906
rect 290 2883 301 2886
rect 306 2886 309 2926
rect 306 2883 317 2886
rect 290 2836 293 2883
rect 290 2833 301 2836
rect 290 2803 293 2816
rect 298 2803 301 2833
rect 306 2813 309 2826
rect 314 2803 317 2883
rect 274 2733 277 2746
rect 282 2723 285 2776
rect 322 2763 325 2816
rect 330 2773 333 2806
rect 290 2703 293 2736
rect 282 2666 285 2696
rect 282 2663 293 2666
rect 266 2653 277 2656
rect 274 2636 277 2653
rect 274 2633 281 2636
rect 226 2593 237 2596
rect 246 2623 253 2626
rect 218 2533 221 2546
rect 182 2523 189 2526
rect 162 2453 173 2456
rect 138 2263 145 2266
rect 122 2223 129 2226
rect 126 2076 129 2223
rect 138 2213 141 2263
rect 138 2113 141 2126
rect 154 2076 157 2286
rect 90 1973 117 1976
rect 90 1956 93 1973
rect 82 1953 93 1956
rect 90 1933 93 1953
rect 66 1893 77 1896
rect 74 1766 77 1893
rect 66 1763 77 1766
rect 66 1296 69 1763
rect 90 1696 93 1856
rect 82 1693 93 1696
rect 82 1596 85 1693
rect 114 1686 117 1973
rect 122 2073 129 2076
rect 150 2073 157 2076
rect 162 2106 165 2453
rect 170 2403 173 2416
rect 178 2403 181 2436
rect 170 2323 173 2336
rect 178 2213 181 2336
rect 186 2286 189 2523
rect 202 2513 205 2526
rect 210 2493 213 2526
rect 226 2523 229 2593
rect 246 2556 249 2623
rect 258 2593 261 2616
rect 278 2566 281 2633
rect 274 2563 281 2566
rect 242 2553 249 2556
rect 234 2513 237 2536
rect 242 2446 245 2553
rect 258 2533 261 2556
rect 274 2543 277 2563
rect 290 2496 293 2663
rect 306 2623 309 2736
rect 346 2636 349 2896
rect 378 2886 381 2926
rect 378 2883 397 2886
rect 362 2803 365 2856
rect 370 2793 373 2816
rect 354 2723 357 2746
rect 314 2633 349 2636
rect 314 2596 317 2633
rect 330 2623 365 2626
rect 330 2613 333 2623
rect 322 2603 333 2606
rect 314 2593 325 2596
rect 306 2523 309 2536
rect 210 2443 245 2446
rect 194 2333 197 2416
rect 210 2363 213 2443
rect 218 2403 221 2426
rect 202 2336 205 2356
rect 226 2346 229 2436
rect 242 2403 253 2406
rect 226 2343 237 2346
rect 202 2333 213 2336
rect 218 2333 229 2336
rect 234 2326 237 2343
rect 242 2333 245 2346
rect 194 2303 197 2326
rect 218 2323 237 2326
rect 234 2303 237 2323
rect 186 2283 193 2286
rect 190 2206 193 2283
rect 186 2203 193 2206
rect 170 2123 173 2136
rect 162 2103 173 2106
rect 122 1836 125 2073
rect 130 1853 133 2056
rect 150 1976 153 2073
rect 150 1973 157 1976
rect 122 1833 129 1836
rect 74 1593 85 1596
rect 98 1683 117 1686
rect 74 1386 77 1593
rect 98 1576 101 1683
rect 126 1676 129 1833
rect 138 1803 141 1926
rect 146 1773 149 1836
rect 138 1723 141 1746
rect 90 1573 101 1576
rect 122 1673 129 1676
rect 90 1413 93 1573
rect 122 1503 125 1673
rect 154 1606 157 1973
rect 162 1733 165 2103
rect 170 1916 173 2036
rect 178 2013 181 2046
rect 178 1933 181 1956
rect 170 1913 177 1916
rect 174 1846 177 1913
rect 170 1843 177 1846
rect 170 1813 173 1843
rect 186 1833 189 2203
rect 194 2123 197 2146
rect 202 2133 205 2176
rect 210 2163 213 2296
rect 250 2226 253 2366
rect 258 2316 261 2496
rect 282 2493 293 2496
rect 282 2436 285 2493
rect 322 2476 325 2593
rect 266 2433 285 2436
rect 318 2473 325 2476
rect 266 2376 269 2433
rect 282 2393 285 2406
rect 306 2376 309 2416
rect 266 2373 273 2376
rect 270 2326 273 2373
rect 290 2373 309 2376
rect 290 2336 293 2373
rect 282 2333 293 2336
rect 298 2326 301 2336
rect 306 2333 309 2356
rect 318 2346 321 2473
rect 330 2356 333 2586
rect 338 2546 341 2616
rect 346 2613 357 2616
rect 346 2593 349 2606
rect 338 2543 345 2546
rect 342 2456 345 2543
rect 342 2453 349 2456
rect 330 2353 341 2356
rect 318 2343 325 2346
rect 322 2326 325 2343
rect 330 2333 333 2346
rect 270 2323 285 2326
rect 258 2313 269 2316
rect 266 2266 269 2313
rect 282 2286 285 2323
rect 290 2303 293 2326
rect 298 2323 309 2326
rect 322 2323 333 2326
rect 322 2306 325 2316
rect 306 2303 325 2306
rect 282 2283 293 2286
rect 266 2263 277 2266
rect 242 2223 253 2226
rect 242 2176 245 2223
rect 258 2183 261 2216
rect 242 2173 253 2176
rect 250 2156 253 2173
rect 210 2153 253 2156
rect 202 2103 205 2126
rect 210 2096 213 2153
rect 218 2113 221 2136
rect 234 2133 237 2146
rect 266 2136 269 2176
rect 250 2133 269 2136
rect 226 2123 245 2126
rect 226 2106 229 2123
rect 242 2113 245 2123
rect 202 2093 213 2096
rect 218 2103 229 2106
rect 194 2013 197 2026
rect 202 2013 205 2093
rect 218 2013 221 2103
rect 250 2086 253 2133
rect 234 2083 253 2086
rect 194 1973 197 2006
rect 202 2003 213 2006
rect 226 2003 229 2026
rect 234 1973 237 2083
rect 250 1976 253 2036
rect 274 1976 277 2263
rect 290 2206 293 2283
rect 306 2236 309 2303
rect 306 2233 317 2236
rect 246 1973 253 1976
rect 258 1973 277 1976
rect 282 2203 293 2206
rect 170 1736 173 1806
rect 178 1803 188 1806
rect 194 1796 197 1816
rect 202 1803 205 1926
rect 210 1796 213 1816
rect 218 1803 221 1936
rect 246 1856 249 1973
rect 246 1853 253 1856
rect 242 1806 245 1836
rect 226 1803 245 1806
rect 194 1793 229 1796
rect 170 1733 181 1736
rect 186 1716 189 1776
rect 178 1713 189 1716
rect 178 1626 181 1713
rect 194 1646 197 1786
rect 202 1783 213 1786
rect 202 1733 205 1783
rect 202 1713 205 1726
rect 210 1656 213 1736
rect 218 1733 221 1746
rect 226 1723 229 1793
rect 250 1763 253 1853
rect 258 1803 261 1973
rect 266 1866 269 1926
rect 282 1873 285 2203
rect 306 2196 309 2216
rect 314 2203 317 2233
rect 306 2193 317 2196
rect 290 2133 293 2186
rect 306 2126 309 2136
rect 314 2133 317 2193
rect 322 2166 325 2296
rect 330 2223 333 2323
rect 338 2313 341 2353
rect 338 2213 341 2306
rect 346 2233 349 2453
rect 354 2346 357 2606
rect 362 2573 365 2623
rect 370 2603 373 2706
rect 378 2566 381 2806
rect 386 2703 389 2816
rect 394 2803 397 2883
rect 402 2636 405 2946
rect 410 2853 413 2926
rect 418 2896 421 2936
rect 442 2933 445 2966
rect 530 2936 533 2976
rect 650 2963 653 3006
rect 530 2933 541 2936
rect 418 2893 429 2896
rect 426 2826 429 2893
rect 418 2823 429 2826
rect 410 2793 413 2806
rect 418 2733 421 2823
rect 426 2783 429 2806
rect 442 2786 445 2916
rect 466 2886 469 2926
rect 522 2886 525 2926
rect 450 2883 469 2886
rect 474 2883 525 2886
rect 450 2803 453 2883
rect 458 2813 461 2826
rect 442 2783 461 2786
rect 466 2783 469 2806
rect 474 2803 477 2883
rect 538 2876 541 2933
rect 562 2903 565 2956
rect 490 2826 493 2876
rect 530 2873 541 2876
rect 486 2823 493 2826
rect 434 2733 437 2746
rect 418 2713 421 2726
rect 362 2563 381 2566
rect 386 2633 405 2636
rect 362 2533 365 2563
rect 370 2533 381 2536
rect 362 2486 365 2526
rect 370 2493 373 2526
rect 386 2523 389 2633
rect 394 2486 397 2556
rect 362 2483 397 2486
rect 402 2476 405 2626
rect 426 2563 429 2726
rect 442 2723 445 2776
rect 450 2643 453 2736
rect 458 2706 461 2783
rect 486 2776 489 2823
rect 498 2783 501 2816
rect 506 2803 509 2866
rect 486 2773 493 2776
rect 490 2746 493 2773
rect 474 2733 477 2746
rect 490 2743 501 2746
rect 458 2703 469 2706
rect 434 2583 437 2626
rect 442 2593 445 2616
rect 450 2613 453 2636
rect 362 2353 365 2416
rect 370 2346 373 2416
rect 354 2343 373 2346
rect 378 2343 381 2406
rect 386 2366 389 2476
rect 394 2473 405 2476
rect 394 2396 397 2473
rect 418 2446 421 2546
rect 418 2443 425 2446
rect 410 2413 413 2436
rect 402 2403 413 2406
rect 394 2393 405 2396
rect 386 2363 397 2366
rect 354 2316 357 2343
rect 362 2333 373 2336
rect 378 2326 381 2336
rect 386 2333 389 2356
rect 354 2313 361 2316
rect 358 2226 361 2313
rect 370 2303 373 2326
rect 378 2323 389 2326
rect 394 2293 397 2363
rect 346 2206 349 2226
rect 330 2173 333 2206
rect 338 2203 349 2206
rect 354 2223 361 2226
rect 322 2163 333 2166
rect 290 1906 293 2126
rect 298 2113 301 2126
rect 306 2123 317 2126
rect 298 2013 301 2026
rect 314 1936 317 2096
rect 298 1933 317 1936
rect 298 1923 301 1933
rect 290 1903 297 1906
rect 266 1863 285 1866
rect 266 1713 269 1776
rect 274 1656 277 1826
rect 282 1803 285 1863
rect 294 1826 297 1903
rect 294 1823 301 1826
rect 290 1793 293 1816
rect 298 1786 301 1823
rect 306 1803 309 1926
rect 322 1923 325 2156
rect 330 2026 333 2163
rect 338 2073 341 2203
rect 354 2153 357 2223
rect 362 2193 365 2206
rect 402 2203 405 2393
rect 422 2386 425 2443
rect 434 2403 437 2486
rect 442 2403 445 2526
rect 450 2466 453 2586
rect 466 2576 469 2703
rect 474 2663 477 2716
rect 482 2626 485 2676
rect 458 2573 469 2576
rect 474 2623 485 2626
rect 458 2473 461 2573
rect 474 2566 477 2623
rect 482 2613 493 2616
rect 498 2606 501 2743
rect 514 2736 517 2816
rect 530 2803 533 2873
rect 570 2843 573 2856
rect 586 2836 589 2926
rect 642 2906 645 2926
rect 634 2903 645 2906
rect 538 2833 589 2836
rect 594 2843 621 2846
rect 538 2803 541 2833
rect 594 2826 597 2843
rect 546 2796 549 2826
rect 546 2793 553 2796
rect 466 2563 477 2566
rect 482 2603 501 2606
rect 506 2733 517 2736
rect 466 2533 469 2563
rect 466 2486 469 2506
rect 466 2483 477 2486
rect 450 2463 469 2466
rect 450 2403 453 2436
rect 458 2393 461 2456
rect 418 2383 425 2386
rect 418 2366 421 2383
rect 466 2376 469 2463
rect 474 2423 477 2483
rect 410 2363 421 2366
rect 462 2373 469 2376
rect 410 2306 413 2363
rect 426 2333 429 2346
rect 450 2323 453 2336
rect 462 2306 465 2373
rect 410 2303 429 2306
rect 462 2303 469 2306
rect 474 2303 477 2406
rect 482 2403 485 2603
rect 490 2563 493 2596
rect 506 2563 509 2733
rect 522 2723 525 2746
rect 514 2673 517 2706
rect 538 2703 541 2776
rect 550 2726 553 2793
rect 546 2723 553 2726
rect 546 2706 549 2723
rect 546 2703 557 2706
rect 546 2686 549 2703
rect 530 2683 549 2686
rect 490 2366 493 2536
rect 514 2533 517 2666
rect 522 2603 525 2636
rect 530 2586 533 2683
rect 562 2673 565 2826
rect 570 2823 597 2826
rect 570 2803 573 2823
rect 578 2793 581 2806
rect 570 2763 589 2766
rect 594 2763 597 2816
rect 602 2803 605 2836
rect 610 2803 613 2816
rect 618 2813 621 2843
rect 634 2826 637 2903
rect 634 2823 645 2826
rect 650 2823 653 2936
rect 690 2933 693 3016
rect 698 2956 701 3023
rect 786 3016 789 3036
rect 858 3033 861 3126
rect 890 3123 893 3136
rect 898 3113 901 3216
rect 922 3196 925 3216
rect 938 3203 941 3216
rect 946 3196 949 3206
rect 922 3193 949 3196
rect 986 3183 989 3206
rect 994 3203 997 3216
rect 1002 3206 1005 3223
rect 1002 3203 1009 3206
rect 1018 3203 1021 3233
rect 906 3126 909 3136
rect 962 3133 965 3176
rect 906 3123 917 3126
rect 946 3123 973 3126
rect 970 3103 973 3123
rect 994 3116 997 3196
rect 1006 3136 1009 3203
rect 1026 3156 1029 3316
rect 1058 3216 1061 3326
rect 1034 3213 1053 3216
rect 1058 3213 1077 3216
rect 1058 3166 1061 3206
rect 1066 3173 1069 3206
rect 1058 3163 1069 3166
rect 1026 3153 1045 3156
rect 1006 3133 1021 3136
rect 1026 3133 1029 3153
rect 990 3113 997 3116
rect 990 3056 993 3113
rect 1002 3103 1005 3126
rect 978 3053 993 3056
rect 722 3013 733 3016
rect 698 2953 709 2956
rect 722 2936 725 3013
rect 754 2963 757 3006
rect 778 2976 781 3016
rect 786 3013 797 3016
rect 762 2973 781 2976
rect 706 2926 709 2936
rect 714 2933 725 2936
rect 746 2933 757 2936
rect 762 2933 765 2973
rect 794 2966 797 3013
rect 786 2963 797 2966
rect 658 2913 661 2926
rect 698 2863 701 2926
rect 706 2923 717 2926
rect 722 2873 725 2933
rect 746 2916 749 2926
rect 754 2923 765 2926
rect 770 2923 773 2946
rect 746 2913 773 2916
rect 658 2823 685 2826
rect 642 2806 645 2823
rect 618 2803 645 2806
rect 562 2636 565 2646
rect 570 2643 573 2763
rect 586 2756 589 2763
rect 578 2723 581 2756
rect 586 2753 613 2756
rect 586 2733 589 2746
rect 602 2726 605 2736
rect 610 2733 613 2753
rect 594 2703 597 2726
rect 602 2723 613 2726
rect 578 2693 605 2696
rect 578 2683 581 2693
rect 594 2636 597 2686
rect 546 2616 549 2636
rect 562 2633 597 2636
rect 538 2613 549 2616
rect 538 2603 541 2613
rect 554 2606 557 2616
rect 546 2603 557 2606
rect 562 2603 565 2633
rect 526 2583 533 2586
rect 498 2483 501 2526
rect 506 2443 509 2496
rect 514 2453 517 2526
rect 526 2506 529 2583
rect 538 2533 541 2596
rect 522 2503 529 2506
rect 538 2503 541 2516
rect 522 2473 525 2503
rect 546 2496 549 2536
rect 534 2493 549 2496
rect 534 2436 537 2493
rect 530 2433 537 2436
rect 506 2403 509 2416
rect 490 2363 497 2366
rect 426 2196 429 2303
rect 466 2283 469 2303
rect 494 2286 497 2363
rect 506 2323 509 2386
rect 530 2376 533 2433
rect 514 2333 517 2376
rect 522 2373 533 2376
rect 522 2316 525 2373
rect 538 2353 541 2416
rect 546 2413 549 2486
rect 554 2343 557 2603
rect 562 2533 565 2566
rect 570 2533 573 2626
rect 578 2613 589 2616
rect 586 2563 589 2613
rect 570 2503 573 2526
rect 578 2413 581 2526
rect 586 2483 589 2536
rect 490 2283 497 2286
rect 514 2313 525 2316
rect 422 2193 429 2196
rect 354 2033 357 2136
rect 378 2123 381 2166
rect 402 2136 405 2156
rect 394 2133 405 2136
rect 378 2036 381 2116
rect 370 2033 381 2036
rect 394 2036 397 2133
rect 422 2106 425 2193
rect 434 2123 437 2266
rect 442 2253 477 2256
rect 442 2213 445 2253
rect 418 2103 425 2106
rect 418 2086 421 2103
rect 410 2083 421 2086
rect 394 2033 405 2036
rect 330 2023 357 2026
rect 314 1803 317 1836
rect 330 1816 333 2023
rect 338 1973 341 2006
rect 346 1996 349 2016
rect 354 2013 357 2023
rect 362 2003 365 2026
rect 370 2013 373 2033
rect 378 2013 389 2016
rect 378 2003 381 2013
rect 386 1996 389 2006
rect 346 1993 389 1996
rect 386 1983 389 1993
rect 346 1933 349 1946
rect 394 1936 397 2016
rect 402 2013 405 2033
rect 402 1973 405 1986
rect 410 1943 413 2083
rect 418 1986 421 2016
rect 434 2013 437 2116
rect 442 2103 445 2186
rect 450 2063 453 2236
rect 474 2176 477 2253
rect 466 2173 477 2176
rect 490 2173 493 2283
rect 514 2246 517 2313
rect 538 2273 541 2336
rect 546 2323 565 2326
rect 562 2303 565 2316
rect 570 2266 573 2336
rect 562 2263 573 2266
rect 506 2243 517 2246
rect 466 2136 469 2173
rect 466 2133 477 2136
rect 490 2126 493 2136
rect 498 2133 501 2206
rect 506 2203 509 2243
rect 482 2113 485 2126
rect 490 2123 501 2126
rect 442 2013 453 2016
rect 426 2003 437 2006
rect 442 2003 445 2013
rect 458 2006 461 2026
rect 450 2003 461 2006
rect 474 1986 477 2006
rect 498 2003 501 2016
rect 418 1983 429 1986
rect 426 1936 429 1983
rect 466 1983 477 1986
rect 386 1933 397 1936
rect 418 1933 429 1936
rect 386 1876 389 1933
rect 394 1886 397 1926
rect 418 1896 421 1933
rect 418 1893 429 1896
rect 394 1883 409 1886
rect 386 1873 397 1876
rect 330 1813 341 1816
rect 290 1783 301 1786
rect 290 1766 293 1783
rect 286 1763 293 1766
rect 286 1696 289 1763
rect 286 1693 293 1696
rect 290 1673 293 1693
rect 210 1653 229 1656
rect 274 1653 285 1656
rect 194 1643 205 1646
rect 178 1623 189 1626
rect 154 1603 165 1606
rect 130 1523 133 1546
rect 130 1486 133 1516
rect 122 1483 133 1486
rect 122 1436 125 1483
rect 122 1433 133 1436
rect 130 1413 133 1433
rect 90 1386 93 1406
rect 138 1396 141 1596
rect 74 1383 93 1386
rect 66 1293 77 1296
rect 74 1046 77 1293
rect 66 1043 77 1046
rect 66 753 69 1043
rect 74 976 77 1026
rect 90 976 93 1383
rect 134 1393 141 1396
rect 114 1023 117 1366
rect 122 1323 125 1346
rect 134 1286 137 1393
rect 162 1286 165 1603
rect 134 1283 141 1286
rect 138 1196 141 1283
rect 154 1283 165 1286
rect 130 1193 141 1196
rect 114 993 117 1016
rect 74 973 81 976
rect 90 973 125 976
rect 78 896 81 973
rect 98 923 101 936
rect 78 893 85 896
rect 82 836 85 893
rect 122 886 125 973
rect 118 883 125 886
rect 82 833 93 836
rect 90 656 93 833
rect 118 766 121 883
rect 130 776 133 1193
rect 146 1113 149 1226
rect 154 1103 157 1283
rect 162 1163 165 1216
rect 178 1183 181 1326
rect 170 1133 173 1156
rect 178 1123 181 1146
rect 146 923 149 946
rect 162 906 165 1076
rect 178 1013 181 1026
rect 170 1003 181 1006
rect 170 916 173 1003
rect 178 923 181 936
rect 170 913 181 916
rect 162 903 173 906
rect 170 876 173 903
rect 162 873 173 876
rect 138 793 141 816
rect 162 796 165 873
rect 178 803 181 913
rect 186 873 189 1623
rect 202 1593 205 1643
rect 226 1596 229 1653
rect 250 1613 253 1626
rect 218 1593 229 1596
rect 202 1523 205 1536
rect 210 1533 213 1556
rect 218 1523 221 1593
rect 282 1576 285 1653
rect 306 1626 309 1766
rect 274 1573 285 1576
rect 298 1623 309 1626
rect 226 1513 229 1536
rect 234 1516 237 1526
rect 250 1516 253 1536
rect 274 1523 277 1573
rect 298 1556 301 1623
rect 314 1563 317 1616
rect 330 1613 333 1806
rect 338 1706 341 1813
rect 346 1723 349 1806
rect 354 1793 357 1816
rect 378 1756 381 1846
rect 378 1753 389 1756
rect 386 1723 389 1753
rect 394 1733 397 1873
rect 406 1826 409 1883
rect 426 1846 429 1893
rect 418 1843 429 1846
rect 406 1823 413 1826
rect 410 1806 413 1823
rect 418 1813 421 1843
rect 410 1803 429 1806
rect 434 1756 437 1816
rect 442 1803 445 1926
rect 450 1883 453 1936
rect 466 1833 469 1983
rect 474 1923 477 1976
rect 498 1943 501 1996
rect 506 1936 509 2156
rect 514 2146 517 2216
rect 522 2203 525 2226
rect 530 2156 533 2216
rect 522 2153 533 2156
rect 538 2146 541 2206
rect 546 2153 549 2206
rect 514 2143 533 2146
rect 538 2143 549 2146
rect 554 2143 557 2246
rect 562 2193 565 2263
rect 578 2236 581 2386
rect 570 2233 581 2236
rect 570 2206 573 2233
rect 578 2213 581 2226
rect 570 2203 581 2206
rect 530 2136 533 2143
rect 514 2083 517 2136
rect 522 2056 525 2136
rect 530 2133 541 2136
rect 530 2113 533 2126
rect 518 2053 525 2056
rect 518 1986 521 2053
rect 518 1983 525 1986
rect 482 1933 493 1936
rect 498 1933 509 1936
rect 498 1853 501 1933
rect 434 1753 445 1756
rect 418 1706 421 1726
rect 338 1703 345 1706
rect 342 1606 345 1703
rect 410 1703 421 1706
rect 410 1626 413 1703
rect 434 1656 437 1736
rect 442 1723 445 1753
rect 466 1746 469 1826
rect 482 1803 485 1816
rect 466 1743 477 1746
rect 450 1726 453 1736
rect 458 1733 469 1736
rect 450 1723 461 1726
rect 466 1713 469 1733
rect 434 1653 461 1656
rect 282 1533 285 1556
rect 290 1553 301 1556
rect 234 1513 245 1516
rect 250 1513 261 1516
rect 242 1486 245 1506
rect 238 1483 245 1486
rect 194 1413 197 1426
rect 238 1416 241 1483
rect 258 1466 261 1513
rect 250 1463 261 1466
rect 250 1423 253 1463
rect 238 1413 245 1416
rect 258 1413 261 1446
rect 290 1436 293 1553
rect 298 1533 301 1546
rect 306 1533 317 1536
rect 322 1533 325 1606
rect 338 1603 345 1606
rect 354 1603 357 1626
rect 410 1623 421 1626
rect 362 1613 381 1616
rect 306 1513 309 1526
rect 306 1436 309 1456
rect 282 1433 293 1436
rect 302 1433 309 1436
rect 210 1363 213 1406
rect 194 1333 205 1336
rect 194 1246 197 1333
rect 202 1313 205 1326
rect 210 1253 213 1356
rect 242 1346 245 1413
rect 274 1376 277 1416
rect 266 1373 277 1376
rect 218 1333 221 1346
rect 242 1343 249 1346
rect 226 1246 229 1326
rect 234 1313 237 1336
rect 246 1296 249 1343
rect 266 1333 269 1373
rect 282 1363 285 1433
rect 246 1293 253 1296
rect 194 1243 205 1246
rect 194 1213 197 1226
rect 194 1106 197 1206
rect 202 1203 205 1243
rect 210 1243 229 1246
rect 202 1133 205 1166
rect 210 1123 213 1243
rect 226 1223 229 1243
rect 234 1206 237 1256
rect 250 1226 253 1293
rect 218 1153 221 1206
rect 230 1203 237 1206
rect 242 1223 253 1226
rect 218 1133 221 1146
rect 230 1116 233 1203
rect 230 1113 237 1116
rect 194 1103 213 1106
rect 186 813 189 826
rect 162 793 173 796
rect 130 773 149 776
rect 114 763 121 766
rect 114 706 117 763
rect 146 733 149 773
rect 170 746 173 793
rect 170 743 177 746
rect 114 703 125 706
rect 74 653 93 656
rect 74 636 77 653
rect 70 633 77 636
rect 70 586 73 633
rect 70 583 77 586
rect 74 506 77 583
rect 90 576 93 606
rect 122 576 125 703
rect 174 676 177 743
rect 170 673 177 676
rect 170 653 173 673
rect 138 593 141 616
rect 178 613 181 646
rect 186 623 189 726
rect 186 586 189 606
rect 90 573 125 576
rect 178 583 189 586
rect 98 533 101 573
rect 146 513 149 526
rect 74 503 101 506
rect 98 203 101 503
rect 178 446 181 583
rect 194 553 197 1096
rect 210 1036 213 1103
rect 234 1093 237 1113
rect 242 1106 245 1223
rect 250 1203 269 1206
rect 274 1196 277 1256
rect 258 1193 277 1196
rect 242 1103 249 1106
rect 246 1046 249 1103
rect 246 1043 253 1046
rect 202 1033 213 1036
rect 202 933 205 1033
rect 210 993 213 1006
rect 218 986 221 1016
rect 226 1013 237 1016
rect 226 1003 229 1013
rect 242 1006 245 1026
rect 234 1003 245 1006
rect 250 993 253 1043
rect 210 983 221 986
rect 202 913 205 926
rect 202 786 205 906
rect 210 876 213 983
rect 218 956 221 983
rect 258 973 261 1193
rect 218 953 261 956
rect 250 933 253 946
rect 242 896 245 926
rect 258 903 261 953
rect 266 896 269 1086
rect 274 983 277 1006
rect 282 1003 285 1216
rect 290 1086 293 1426
rect 302 1346 305 1433
rect 302 1343 309 1346
rect 298 1096 301 1326
rect 306 1213 309 1343
rect 314 1246 317 1466
rect 330 1366 333 1546
rect 338 1523 341 1603
rect 346 1446 349 1566
rect 362 1546 365 1613
rect 370 1563 373 1606
rect 362 1543 373 1546
rect 346 1443 357 1446
rect 362 1443 365 1536
rect 370 1513 373 1543
rect 378 1463 381 1536
rect 386 1533 389 1606
rect 418 1523 421 1623
rect 458 1613 461 1653
rect 434 1543 437 1606
rect 426 1456 429 1536
rect 434 1513 437 1526
rect 378 1453 429 1456
rect 330 1363 337 1366
rect 334 1276 337 1363
rect 330 1273 337 1276
rect 330 1253 333 1273
rect 314 1243 341 1246
rect 330 1213 333 1226
rect 322 1166 325 1206
rect 306 1163 325 1166
rect 306 1123 309 1163
rect 338 1146 341 1243
rect 330 1143 341 1146
rect 330 1096 333 1143
rect 298 1093 309 1096
rect 330 1093 341 1096
rect 290 1083 301 1086
rect 298 1013 301 1083
rect 338 1073 341 1093
rect 346 1066 349 1326
rect 354 1296 357 1443
rect 378 1413 381 1453
rect 442 1436 445 1536
rect 450 1533 453 1556
rect 466 1446 469 1536
rect 474 1523 477 1743
rect 482 1723 485 1736
rect 498 1723 501 1736
rect 506 1706 509 1926
rect 514 1896 517 1966
rect 522 1956 525 1983
rect 538 1963 541 2133
rect 546 2093 549 2143
rect 554 2103 557 2126
rect 546 2006 549 2066
rect 554 2013 557 2026
rect 546 2003 557 2006
rect 562 2003 565 2186
rect 570 2116 573 2166
rect 578 2123 581 2203
rect 586 2193 589 2466
rect 594 2406 597 2616
rect 602 2613 605 2693
rect 602 2573 605 2606
rect 610 2566 613 2656
rect 618 2576 621 2803
rect 650 2776 653 2806
rect 626 2773 653 2776
rect 626 2586 629 2773
rect 658 2756 661 2823
rect 666 2796 669 2806
rect 674 2803 677 2816
rect 682 2803 685 2823
rect 666 2793 693 2796
rect 674 2773 685 2776
rect 650 2753 661 2756
rect 642 2733 645 2746
rect 650 2736 653 2753
rect 658 2743 669 2746
rect 650 2733 661 2736
rect 642 2723 653 2726
rect 658 2716 661 2733
rect 658 2713 665 2716
rect 634 2613 637 2646
rect 650 2613 653 2686
rect 662 2626 665 2713
rect 658 2623 665 2626
rect 642 2596 645 2606
rect 658 2603 661 2623
rect 642 2593 669 2596
rect 674 2586 677 2766
rect 682 2743 685 2773
rect 690 2756 693 2776
rect 698 2763 701 2806
rect 690 2753 701 2756
rect 698 2736 701 2753
rect 706 2743 709 2806
rect 714 2766 717 2846
rect 722 2773 725 2826
rect 730 2823 749 2826
rect 730 2813 733 2823
rect 738 2793 741 2816
rect 746 2803 749 2823
rect 754 2813 757 2836
rect 754 2796 757 2806
rect 762 2803 765 2846
rect 770 2813 773 2913
rect 770 2796 773 2806
rect 754 2793 773 2796
rect 714 2763 725 2766
rect 682 2643 685 2736
rect 698 2733 709 2736
rect 690 2683 693 2726
rect 698 2703 701 2726
rect 682 2613 693 2616
rect 626 2583 661 2586
rect 618 2573 629 2576
rect 602 2546 605 2566
rect 610 2563 621 2566
rect 626 2556 629 2573
rect 610 2553 629 2556
rect 602 2543 621 2546
rect 602 2533 613 2536
rect 602 2473 605 2525
rect 610 2503 613 2533
rect 618 2523 621 2543
rect 634 2536 637 2556
rect 626 2533 637 2536
rect 610 2493 629 2496
rect 594 2403 605 2406
rect 610 2403 613 2466
rect 618 2413 621 2486
rect 594 2373 597 2396
rect 570 2113 581 2116
rect 586 2113 589 2186
rect 594 2183 597 2346
rect 602 2313 605 2403
rect 618 2373 621 2406
rect 602 2213 605 2276
rect 522 1953 533 1956
rect 530 1943 533 1953
rect 530 1923 533 1936
rect 554 1896 557 2003
rect 514 1893 525 1896
rect 554 1893 561 1896
rect 522 1836 525 1893
rect 502 1703 509 1706
rect 514 1833 525 1836
rect 502 1576 505 1703
rect 502 1573 509 1576
rect 506 1553 509 1573
rect 514 1536 517 1833
rect 522 1733 525 1816
rect 546 1766 549 1866
rect 542 1763 549 1766
rect 522 1613 525 1716
rect 530 1703 533 1726
rect 530 1603 533 1616
rect 542 1576 545 1763
rect 558 1756 561 1893
rect 570 1863 573 2106
rect 578 2003 581 2113
rect 594 2103 597 2126
rect 594 2046 597 2086
rect 602 2066 605 2136
rect 610 2116 613 2326
rect 618 2316 621 2336
rect 626 2333 629 2493
rect 634 2356 637 2526
rect 642 2513 645 2536
rect 650 2523 653 2566
rect 658 2533 661 2583
rect 666 2583 677 2586
rect 658 2503 661 2526
rect 666 2496 669 2583
rect 642 2493 669 2496
rect 642 2423 645 2493
rect 642 2393 645 2406
rect 650 2393 653 2466
rect 674 2453 677 2536
rect 666 2403 669 2416
rect 674 2403 677 2436
rect 634 2353 661 2356
rect 642 2333 645 2346
rect 618 2313 625 2316
rect 622 2246 625 2313
rect 622 2243 629 2246
rect 618 2213 621 2236
rect 618 2123 621 2196
rect 626 2163 629 2243
rect 626 2133 629 2146
rect 634 2116 637 2326
rect 650 2283 653 2326
rect 658 2303 661 2353
rect 666 2343 669 2396
rect 666 2283 669 2336
rect 650 2223 653 2276
rect 642 2166 645 2206
rect 650 2203 653 2216
rect 642 2163 653 2166
rect 642 2133 645 2156
rect 650 2136 653 2163
rect 658 2146 661 2226
rect 666 2213 669 2236
rect 674 2233 677 2396
rect 682 2233 685 2606
rect 690 2563 693 2613
rect 698 2593 701 2616
rect 690 2463 693 2536
rect 698 2523 701 2556
rect 706 2526 709 2733
rect 714 2683 717 2736
rect 722 2723 725 2763
rect 730 2716 733 2736
rect 738 2723 741 2736
rect 746 2723 749 2776
rect 770 2733 773 2746
rect 778 2733 781 2936
rect 786 2923 789 2963
rect 834 2946 837 3016
rect 866 2993 869 3006
rect 890 2976 893 3016
rect 794 2943 837 2946
rect 842 2973 893 2976
rect 794 2933 797 2943
rect 802 2933 813 2936
rect 842 2933 845 2973
rect 946 2946 949 3016
rect 978 2993 981 3053
rect 1018 3023 1021 3133
rect 1042 3063 1045 3153
rect 1066 3123 1069 3163
rect 1074 3086 1077 3213
rect 1082 3146 1085 3336
rect 1090 3323 1093 3403
rect 1106 3376 1109 3536
rect 1114 3533 1117 3573
rect 1138 3566 1141 3633
rect 1146 3583 1149 3643
rect 1130 3563 1141 3566
rect 1130 3533 1133 3563
rect 1138 3553 1141 3563
rect 1114 3513 1117 3526
rect 1122 3493 1125 3526
rect 1138 3523 1141 3536
rect 1146 3453 1149 3536
rect 1154 3533 1157 3596
rect 1170 3556 1173 3683
rect 1190 3656 1193 3723
rect 1202 3666 1205 3816
rect 1210 3783 1213 3806
rect 1226 3773 1229 3816
rect 1274 3813 1277 3833
rect 1282 3823 1293 3826
rect 1314 3823 1317 3833
rect 1234 3783 1237 3806
rect 1290 3756 1293 3816
rect 1298 3793 1301 3806
rect 1330 3786 1333 3816
rect 1346 3803 1349 3816
rect 1330 3783 1341 3786
rect 1258 3743 1261 3756
rect 1290 3753 1301 3756
rect 1210 3713 1213 3726
rect 1202 3663 1209 3666
rect 1190 3653 1197 3656
rect 1162 3546 1165 3556
rect 1170 3553 1189 3556
rect 1162 3543 1181 3546
rect 1178 3533 1181 3543
rect 1130 3413 1133 3446
rect 1154 3403 1157 3416
rect 1162 3396 1165 3526
rect 1178 3506 1181 3526
rect 1174 3503 1181 3506
rect 1174 3446 1177 3503
rect 1186 3463 1189 3553
rect 1194 3533 1197 3653
rect 1206 3606 1209 3663
rect 1242 3626 1245 3726
rect 1266 3706 1269 3736
rect 1290 3733 1293 3746
rect 1282 3713 1285 3726
rect 1266 3703 1293 3706
rect 1218 3613 1221 3626
rect 1242 3623 1253 3626
rect 1202 3603 1209 3606
rect 1202 3583 1205 3603
rect 1250 3566 1253 3623
rect 1274 3613 1277 3646
rect 1242 3563 1253 3566
rect 1242 3546 1245 3563
rect 1274 3553 1277 3606
rect 1282 3566 1285 3666
rect 1290 3603 1293 3703
rect 1298 3596 1301 3753
rect 1306 3733 1309 3776
rect 1306 3706 1309 3726
rect 1314 3723 1317 3746
rect 1338 3706 1341 3783
rect 1354 3733 1357 3756
rect 1354 3713 1357 3726
rect 1362 3713 1365 3776
rect 1394 3773 1397 3816
rect 1426 3813 1429 3913
rect 1482 3846 1485 3983
rect 1498 3943 1501 4016
rect 1534 3966 1537 4033
rect 1546 3993 1549 4016
rect 1578 4013 1581 4103
rect 1534 3963 1541 3966
rect 1538 3946 1541 3963
rect 1514 3933 1517 3946
rect 1538 3943 1549 3946
rect 1498 3903 1501 3926
rect 1546 3896 1549 3943
rect 1538 3893 1549 3896
rect 1482 3843 1493 3846
rect 1458 3803 1461 3816
rect 1490 3776 1493 3843
rect 1506 3793 1509 3816
rect 1482 3773 1493 3776
rect 1482 3756 1485 3773
rect 1466 3753 1485 3756
rect 1394 3743 1453 3746
rect 1306 3703 1317 3706
rect 1338 3703 1349 3706
rect 1314 3626 1317 3703
rect 1346 3666 1349 3703
rect 1346 3663 1353 3666
rect 1306 3623 1317 3626
rect 1306 3603 1309 3623
rect 1338 3613 1341 3636
rect 1350 3606 1353 3663
rect 1370 3626 1373 3726
rect 1402 3716 1405 3736
rect 1426 3733 1445 3736
rect 1450 3733 1453 3743
rect 1394 3713 1405 3716
rect 1394 3656 1397 3713
rect 1394 3653 1405 3656
rect 1402 3636 1405 3653
rect 1402 3633 1413 3636
rect 1370 3623 1405 3626
rect 1370 3613 1373 3623
rect 1410 3616 1413 3633
rect 1418 3623 1421 3726
rect 1426 3713 1429 3726
rect 1386 3613 1397 3616
rect 1402 3613 1413 3616
rect 1426 3613 1429 3666
rect 1314 3596 1317 3606
rect 1298 3593 1317 3596
rect 1346 3603 1353 3606
rect 1282 3563 1313 3566
rect 1242 3543 1253 3546
rect 1194 3446 1197 3526
rect 1218 3503 1221 3526
rect 1174 3443 1181 3446
rect 1194 3443 1205 3446
rect 1178 3403 1181 3443
rect 1154 3393 1165 3396
rect 1106 3373 1125 3376
rect 1090 3223 1093 3256
rect 1098 3243 1101 3336
rect 1106 3323 1109 3366
rect 1098 3163 1101 3236
rect 1082 3143 1093 3146
rect 1090 3086 1093 3143
rect 1106 3123 1109 3296
rect 1114 3223 1117 3336
rect 1122 3316 1125 3373
rect 1130 3323 1133 3346
rect 1154 3343 1157 3393
rect 1170 3333 1173 3386
rect 1122 3313 1141 3316
rect 1138 3266 1141 3313
rect 1130 3263 1141 3266
rect 1122 3186 1125 3246
rect 1114 3183 1125 3186
rect 1074 3083 1085 3086
rect 1090 3083 1097 3086
rect 786 2776 789 2846
rect 794 2803 797 2836
rect 802 2813 805 2926
rect 834 2876 837 2926
rect 834 2873 845 2876
rect 786 2773 797 2776
rect 754 2716 757 2726
rect 730 2713 757 2716
rect 754 2696 757 2713
rect 746 2693 757 2696
rect 714 2586 717 2656
rect 746 2636 749 2693
rect 762 2686 765 2726
rect 770 2696 773 2716
rect 778 2706 781 2726
rect 786 2723 789 2746
rect 794 2723 797 2773
rect 802 2756 805 2806
rect 810 2763 813 2806
rect 818 2793 821 2836
rect 834 2826 837 2836
rect 826 2823 837 2826
rect 802 2753 813 2756
rect 778 2703 789 2706
rect 770 2693 781 2696
rect 762 2683 773 2686
rect 762 2653 765 2676
rect 746 2633 757 2636
rect 722 2613 725 2626
rect 730 2593 733 2606
rect 738 2596 741 2616
rect 738 2593 749 2596
rect 714 2583 741 2586
rect 714 2533 717 2566
rect 706 2523 717 2526
rect 706 2436 709 2516
rect 714 2443 717 2523
rect 674 2173 677 2226
rect 682 2213 685 2226
rect 690 2213 693 2426
rect 698 2413 701 2436
rect 706 2433 717 2436
rect 714 2413 717 2433
rect 698 2403 709 2406
rect 722 2383 725 2526
rect 730 2393 733 2536
rect 738 2533 741 2583
rect 746 2573 749 2593
rect 754 2556 757 2633
rect 746 2553 757 2556
rect 738 2503 741 2516
rect 746 2496 749 2553
rect 762 2546 765 2646
rect 770 2596 773 2683
rect 778 2613 781 2693
rect 786 2683 789 2703
rect 794 2613 797 2656
rect 802 2626 805 2726
rect 810 2636 813 2753
rect 818 2733 821 2786
rect 818 2653 821 2726
rect 826 2643 829 2823
rect 834 2723 837 2776
rect 842 2763 845 2873
rect 850 2863 853 2946
rect 866 2943 949 2946
rect 858 2926 861 2936
rect 866 2933 869 2943
rect 954 2936 957 2976
rect 1002 2956 1005 3016
rect 1058 3006 1061 3016
rect 1042 3003 1061 3006
rect 1066 3003 1069 3076
rect 858 2923 869 2926
rect 858 2906 861 2923
rect 882 2913 885 2926
rect 858 2903 869 2906
rect 866 2856 869 2903
rect 882 2883 893 2886
rect 898 2883 901 2936
rect 914 2913 917 2936
rect 858 2853 869 2856
rect 858 2833 861 2853
rect 850 2806 853 2826
rect 858 2823 877 2826
rect 858 2813 861 2823
rect 850 2803 861 2806
rect 866 2803 869 2816
rect 874 2803 877 2823
rect 850 2736 853 2796
rect 858 2786 861 2803
rect 858 2783 877 2786
rect 882 2783 885 2816
rect 890 2786 893 2883
rect 898 2803 901 2816
rect 906 2803 909 2896
rect 922 2886 925 2936
rect 914 2883 925 2886
rect 914 2806 917 2883
rect 930 2826 933 2936
rect 922 2823 933 2826
rect 922 2813 925 2823
rect 938 2816 941 2936
rect 946 2933 957 2936
rect 962 2953 1005 2956
rect 962 2933 965 2953
rect 946 2836 949 2933
rect 954 2843 957 2926
rect 970 2906 973 2936
rect 970 2903 977 2906
rect 946 2833 957 2836
rect 930 2813 941 2816
rect 954 2813 957 2833
rect 914 2803 925 2806
rect 898 2793 909 2796
rect 890 2783 901 2786
rect 842 2733 853 2736
rect 842 2706 845 2733
rect 838 2703 845 2706
rect 810 2633 829 2636
rect 802 2623 821 2626
rect 802 2613 813 2616
rect 786 2603 797 2606
rect 802 2603 805 2613
rect 770 2593 789 2596
rect 738 2493 749 2496
rect 754 2543 765 2546
rect 738 2423 741 2493
rect 754 2476 757 2543
rect 762 2533 781 2536
rect 746 2473 757 2476
rect 762 2473 765 2526
rect 770 2493 773 2526
rect 738 2376 741 2416
rect 746 2396 749 2473
rect 754 2413 757 2456
rect 778 2423 781 2533
rect 786 2513 789 2593
rect 794 2533 797 2603
rect 810 2553 813 2606
rect 818 2573 821 2623
rect 826 2603 829 2633
rect 838 2586 841 2703
rect 850 2593 853 2726
rect 858 2713 861 2766
rect 866 2673 869 2736
rect 874 2733 877 2783
rect 874 2683 877 2726
rect 882 2723 885 2766
rect 890 2706 893 2736
rect 886 2703 893 2706
rect 886 2646 889 2703
rect 898 2673 901 2783
rect 906 2723 909 2793
rect 930 2786 933 2813
rect 962 2803 965 2886
rect 974 2836 977 2903
rect 970 2833 977 2836
rect 914 2783 933 2786
rect 866 2613 869 2646
rect 886 2643 893 2646
rect 890 2626 893 2643
rect 914 2636 917 2783
rect 970 2756 973 2833
rect 978 2793 981 2806
rect 986 2763 989 2936
rect 994 2783 997 2906
rect 1010 2893 1013 2966
rect 1034 2913 1037 2926
rect 1002 2793 1005 2806
rect 922 2723 925 2756
rect 930 2753 949 2756
rect 954 2753 973 2756
rect 930 2733 933 2753
rect 954 2746 957 2753
rect 938 2743 957 2746
rect 930 2646 933 2726
rect 938 2696 941 2743
rect 946 2726 949 2736
rect 954 2733 965 2736
rect 946 2723 957 2726
rect 946 2703 949 2723
rect 962 2703 965 2733
rect 978 2723 981 2736
rect 1002 2723 1005 2756
rect 938 2693 965 2696
rect 930 2643 941 2646
rect 914 2633 933 2636
rect 890 2623 909 2626
rect 906 2613 909 2623
rect 914 2613 917 2626
rect 834 2583 841 2586
rect 834 2546 837 2583
rect 842 2556 845 2576
rect 858 2573 861 2606
rect 866 2603 877 2606
rect 866 2563 869 2603
rect 842 2553 853 2556
rect 834 2543 845 2546
rect 754 2403 765 2406
rect 746 2393 765 2396
rect 698 2323 701 2346
rect 714 2333 717 2376
rect 722 2373 741 2376
rect 690 2153 693 2206
rect 658 2143 685 2146
rect 650 2133 661 2136
rect 610 2113 629 2116
rect 634 2113 641 2116
rect 650 2113 653 2126
rect 658 2123 661 2133
rect 602 2063 621 2066
rect 594 2043 605 2046
rect 586 1963 589 2016
rect 594 2003 597 2026
rect 602 1986 605 2043
rect 598 1983 605 1986
rect 578 1893 581 1926
rect 598 1876 601 1983
rect 594 1873 601 1876
rect 594 1826 597 1873
rect 554 1753 561 1756
rect 570 1823 597 1826
rect 554 1613 557 1753
rect 562 1603 565 1726
rect 570 1716 573 1823
rect 578 1733 581 1816
rect 586 1803 589 1816
rect 594 1723 597 1806
rect 570 1713 577 1716
rect 574 1626 577 1713
rect 570 1623 577 1626
rect 490 1476 493 1536
rect 510 1533 517 1536
rect 522 1573 545 1576
rect 498 1513 501 1526
rect 510 1486 513 1533
rect 522 1496 525 1573
rect 530 1506 533 1536
rect 546 1533 549 1546
rect 530 1503 541 1506
rect 522 1493 529 1496
rect 510 1483 517 1486
rect 482 1473 493 1476
rect 466 1443 473 1446
rect 426 1433 445 1436
rect 370 1323 373 1336
rect 394 1296 397 1386
rect 354 1293 365 1296
rect 362 1226 365 1293
rect 386 1293 397 1296
rect 354 1223 365 1226
rect 354 1106 357 1223
rect 378 1206 381 1286
rect 362 1123 365 1206
rect 370 1203 381 1206
rect 370 1133 373 1203
rect 386 1196 389 1293
rect 378 1193 389 1196
rect 354 1103 361 1106
rect 330 1063 349 1066
rect 290 1003 317 1006
rect 242 893 269 896
rect 210 873 221 876
rect 218 813 221 873
rect 210 793 213 806
rect 226 793 229 806
rect 234 803 237 826
rect 202 783 213 786
rect 210 766 213 783
rect 242 776 245 893
rect 274 856 277 976
rect 282 933 293 936
rect 266 853 277 856
rect 250 793 253 816
rect 266 776 269 853
rect 234 773 245 776
rect 250 773 269 776
rect 210 763 221 766
rect 218 686 221 763
rect 206 683 221 686
rect 234 686 237 773
rect 234 683 245 686
rect 206 626 209 683
rect 202 623 209 626
rect 178 443 189 446
rect 146 403 149 416
rect 170 413 181 416
rect 186 403 189 443
rect 154 333 181 336
rect 146 213 149 246
rect 178 213 181 333
rect 186 323 189 346
rect 194 213 197 536
rect 202 516 205 623
rect 210 593 213 606
rect 218 546 221 616
rect 234 603 237 616
rect 242 613 245 683
rect 218 543 229 546
rect 210 533 221 536
rect 202 513 209 516
rect 206 436 209 513
rect 218 503 221 526
rect 202 433 209 436
rect 202 323 205 433
rect 226 413 229 543
rect 234 523 237 556
rect 242 543 245 606
rect 250 596 253 773
rect 258 746 261 766
rect 258 743 265 746
rect 262 666 265 743
rect 274 676 277 726
rect 282 723 285 796
rect 290 726 293 886
rect 298 863 301 996
rect 314 993 317 1003
rect 306 856 309 986
rect 298 853 309 856
rect 298 733 301 853
rect 290 723 301 726
rect 282 676 285 686
rect 274 673 285 676
rect 262 663 277 666
rect 258 603 261 626
rect 250 593 261 596
rect 242 513 245 536
rect 250 486 253 566
rect 258 556 261 593
rect 266 563 269 616
rect 258 553 269 556
rect 258 503 261 536
rect 234 483 253 486
rect 210 403 221 406
rect 210 393 213 403
rect 234 396 237 483
rect 242 413 245 426
rect 218 393 237 396
rect 250 393 253 406
rect 258 403 261 436
rect 210 243 213 336
rect 218 306 221 393
rect 250 356 253 386
rect 242 353 253 356
rect 226 333 229 346
rect 242 306 245 353
rect 218 303 229 306
rect 242 303 253 306
rect 226 246 229 303
rect 218 243 229 246
rect 218 226 221 243
rect 210 223 221 226
rect 210 203 213 223
rect 218 203 221 223
rect 250 193 253 303
rect 266 273 269 553
rect 274 403 277 663
rect 282 603 285 673
rect 282 393 285 516
rect 290 433 293 716
rect 298 603 301 723
rect 306 633 309 846
rect 314 833 317 976
rect 322 953 325 1006
rect 330 993 333 1063
rect 358 1026 361 1103
rect 338 946 341 1016
rect 346 1003 349 1026
rect 354 1023 361 1026
rect 322 943 341 946
rect 322 876 325 943
rect 330 933 341 936
rect 338 906 341 926
rect 330 903 341 906
rect 330 893 333 903
rect 346 876 349 956
rect 354 893 357 1023
rect 370 1013 373 1126
rect 378 1106 381 1193
rect 386 1133 389 1146
rect 394 1123 397 1236
rect 402 1203 405 1406
rect 426 1366 429 1433
rect 426 1363 437 1366
rect 410 1146 413 1296
rect 418 1203 421 1326
rect 426 1213 429 1236
rect 410 1143 429 1146
rect 402 1126 405 1136
rect 410 1133 421 1136
rect 402 1123 413 1126
rect 426 1123 429 1143
rect 378 1103 405 1106
rect 322 873 333 876
rect 314 813 317 826
rect 314 733 325 736
rect 314 723 325 726
rect 314 653 317 723
rect 306 613 309 626
rect 306 603 317 606
rect 306 596 309 603
rect 322 596 325 716
rect 330 603 333 873
rect 338 873 349 876
rect 338 803 341 873
rect 338 733 341 746
rect 346 673 349 866
rect 354 813 357 836
rect 354 736 357 806
rect 362 803 365 1006
rect 370 743 373 1006
rect 378 1003 381 1096
rect 402 1046 405 1103
rect 394 1043 405 1046
rect 378 853 381 986
rect 386 976 389 1016
rect 394 983 397 1043
rect 402 1023 429 1026
rect 386 973 397 976
rect 386 933 389 956
rect 394 876 397 973
rect 402 933 405 1023
rect 410 993 413 1006
rect 418 1003 421 1016
rect 426 1013 429 1023
rect 434 1016 437 1363
rect 442 1156 445 1406
rect 470 1396 473 1443
rect 482 1413 485 1473
rect 466 1393 473 1396
rect 450 1333 461 1336
rect 450 1163 453 1333
rect 458 1203 461 1326
rect 466 1173 469 1393
rect 514 1356 517 1483
rect 474 1353 517 1356
rect 526 1356 529 1493
rect 538 1373 541 1503
rect 570 1436 573 1623
rect 586 1613 589 1706
rect 594 1696 597 1716
rect 594 1693 601 1696
rect 598 1606 601 1693
rect 578 1523 581 1606
rect 594 1603 601 1606
rect 594 1566 597 1603
rect 590 1563 597 1566
rect 610 1566 613 2056
rect 618 2013 621 2063
rect 626 2053 629 2113
rect 638 2026 641 2113
rect 634 2023 641 2026
rect 618 1903 621 1926
rect 626 1923 629 2006
rect 618 1803 621 1896
rect 618 1723 621 1736
rect 626 1663 629 1816
rect 634 1616 637 2023
rect 642 1933 645 2006
rect 650 1986 653 2056
rect 658 1993 661 2066
rect 666 2033 669 2126
rect 674 2053 677 2116
rect 682 2083 685 2143
rect 690 2103 693 2126
rect 698 2103 701 2236
rect 706 2096 709 2296
rect 714 2273 717 2326
rect 722 2236 725 2373
rect 738 2336 741 2346
rect 730 2333 741 2336
rect 738 2286 741 2326
rect 746 2293 749 2336
rect 666 2013 677 2016
rect 682 2013 685 2026
rect 690 2013 693 2096
rect 698 2093 709 2096
rect 714 2233 725 2236
rect 730 2283 741 2286
rect 666 1993 669 2006
rect 674 2003 693 2006
rect 650 1983 661 1986
rect 650 1933 653 1946
rect 642 1906 645 1926
rect 658 1923 661 1983
rect 666 1933 669 1976
rect 642 1903 653 1906
rect 650 1766 653 1903
rect 666 1803 669 1926
rect 642 1763 653 1766
rect 674 1763 677 1926
rect 682 1923 685 1996
rect 690 1893 693 2003
rect 698 1843 701 2093
rect 714 2086 717 2233
rect 722 2213 725 2226
rect 730 2156 733 2283
rect 738 2213 741 2276
rect 754 2263 757 2336
rect 762 2316 765 2393
rect 770 2323 773 2416
rect 762 2313 769 2316
rect 766 2256 769 2313
rect 766 2253 773 2256
rect 746 2223 749 2236
rect 738 2183 741 2206
rect 730 2153 741 2156
rect 722 2143 741 2146
rect 722 2123 725 2143
rect 730 2133 741 2136
rect 722 2093 725 2116
rect 706 2083 717 2086
rect 706 1926 709 2083
rect 714 2006 717 2066
rect 722 2056 725 2086
rect 730 2063 733 2133
rect 738 2113 741 2126
rect 746 2103 749 2196
rect 754 2076 757 2226
rect 762 2113 765 2236
rect 770 2233 773 2253
rect 770 2133 773 2226
rect 778 2116 781 2406
rect 786 2323 789 2496
rect 794 2393 797 2526
rect 810 2523 813 2536
rect 834 2523 837 2536
rect 842 2476 845 2543
rect 802 2363 805 2476
rect 834 2473 845 2476
rect 810 2313 813 2426
rect 818 2423 821 2436
rect 818 2403 821 2416
rect 826 2413 829 2446
rect 826 2373 829 2406
rect 834 2396 837 2473
rect 850 2443 853 2553
rect 842 2433 853 2436
rect 858 2426 861 2556
rect 866 2433 869 2466
rect 850 2416 853 2426
rect 858 2423 869 2426
rect 850 2413 861 2416
rect 842 2403 861 2406
rect 834 2393 845 2396
rect 826 2343 837 2346
rect 786 2133 789 2246
rect 794 2223 797 2266
rect 794 2193 797 2216
rect 802 2213 805 2256
rect 770 2083 773 2116
rect 778 2113 785 2116
rect 754 2073 773 2076
rect 722 2053 733 2056
rect 730 2013 733 2053
rect 714 2003 733 2006
rect 714 1933 725 1936
rect 706 1923 717 1926
rect 714 1906 717 1923
rect 682 1813 685 1826
rect 642 1683 645 1763
rect 634 1613 641 1616
rect 610 1563 617 1566
rect 590 1486 593 1563
rect 614 1486 617 1563
rect 626 1523 629 1606
rect 638 1516 641 1613
rect 650 1603 653 1736
rect 658 1693 661 1746
rect 666 1703 669 1736
rect 674 1663 677 1726
rect 706 1723 709 1906
rect 714 1903 721 1906
rect 718 1846 721 1903
rect 730 1856 733 2003
rect 738 1973 741 2006
rect 746 1966 749 2006
rect 738 1963 749 1966
rect 738 1933 741 1963
rect 738 1903 741 1926
rect 746 1863 749 1946
rect 754 1923 757 2016
rect 762 1883 765 2066
rect 770 1993 773 2073
rect 782 2046 785 2113
rect 794 2103 797 2126
rect 802 2123 805 2186
rect 778 2043 785 2046
rect 778 1986 781 2043
rect 786 2003 789 2026
rect 794 2013 797 2096
rect 802 2013 805 2116
rect 810 2043 813 2276
rect 818 2063 821 2286
rect 826 2233 829 2336
rect 834 2323 837 2343
rect 826 2213 829 2226
rect 834 2183 837 2266
rect 842 2216 845 2393
rect 850 2253 853 2336
rect 858 2323 861 2386
rect 850 2223 853 2236
rect 842 2213 853 2216
rect 794 2003 805 2006
rect 770 1983 781 1986
rect 770 1923 773 1983
rect 786 1923 789 1996
rect 794 1933 797 2003
rect 802 1963 805 1996
rect 802 1933 805 1946
rect 810 1856 813 2016
rect 818 1883 821 2056
rect 826 1983 829 2126
rect 834 2123 837 2176
rect 842 2133 845 2206
rect 834 1953 837 2116
rect 842 2103 845 2126
rect 850 2103 853 2213
rect 858 2163 861 2226
rect 866 2176 869 2423
rect 874 2313 877 2596
rect 882 2306 885 2606
rect 890 2573 893 2596
rect 914 2576 917 2606
rect 914 2573 925 2576
rect 890 2523 893 2536
rect 898 2523 901 2566
rect 914 2546 917 2566
rect 906 2543 917 2546
rect 890 2463 893 2486
rect 906 2476 909 2543
rect 898 2473 909 2476
rect 890 2423 893 2436
rect 906 2413 909 2446
rect 914 2406 917 2536
rect 898 2363 901 2406
rect 906 2403 917 2406
rect 922 2376 925 2573
rect 930 2526 933 2633
rect 938 2536 941 2643
rect 946 2546 949 2676
rect 962 2616 965 2693
rect 954 2563 957 2616
rect 962 2613 973 2616
rect 962 2553 965 2606
rect 946 2543 965 2546
rect 938 2533 949 2536
rect 930 2523 941 2526
rect 930 2483 933 2516
rect 930 2386 933 2426
rect 938 2403 941 2523
rect 946 2413 949 2533
rect 954 2513 957 2536
rect 962 2426 965 2543
rect 970 2496 973 2613
rect 978 2596 981 2716
rect 1010 2706 1013 2866
rect 1042 2846 1045 3003
rect 1050 2976 1053 2996
rect 1050 2973 1057 2976
rect 1054 2866 1057 2973
rect 1074 2966 1077 3046
rect 1094 3026 1097 3083
rect 1114 3043 1117 3183
rect 1122 3123 1125 3176
rect 1130 3143 1133 3263
rect 1202 3256 1205 3443
rect 1210 3383 1213 3466
rect 1218 3376 1221 3486
rect 1250 3456 1253 3543
rect 1258 3523 1261 3536
rect 1250 3453 1269 3456
rect 1226 3413 1229 3426
rect 1218 3373 1237 3376
rect 1218 3303 1221 3326
rect 1202 3253 1221 3256
rect 1146 3193 1149 3226
rect 1194 3203 1197 3216
rect 1162 3133 1165 3146
rect 1178 3133 1181 3156
rect 1154 3106 1157 3126
rect 1146 3103 1157 3106
rect 1146 3056 1149 3103
rect 1146 3053 1157 3056
rect 1154 3036 1157 3053
rect 1106 3033 1157 3036
rect 1094 3023 1101 3026
rect 1098 3003 1101 3023
rect 1106 3013 1109 3033
rect 1154 3023 1157 3033
rect 1162 3006 1165 3076
rect 1158 3003 1165 3006
rect 1074 2963 1081 2966
rect 1078 2886 1081 2963
rect 1098 2926 1101 2946
rect 1006 2703 1013 2706
rect 1018 2843 1045 2846
rect 1050 2863 1057 2866
rect 1074 2883 1081 2886
rect 1006 2636 1009 2703
rect 1018 2653 1021 2843
rect 1026 2803 1029 2816
rect 1034 2786 1037 2836
rect 1050 2793 1053 2863
rect 1026 2776 1029 2786
rect 1034 2783 1053 2786
rect 1026 2773 1045 2776
rect 1026 2643 1029 2766
rect 1042 2723 1045 2773
rect 1042 2676 1045 2706
rect 1038 2673 1045 2676
rect 994 2633 1009 2636
rect 986 2603 989 2626
rect 978 2593 989 2596
rect 978 2523 981 2566
rect 978 2503 981 2516
rect 986 2506 989 2593
rect 994 2576 997 2633
rect 1010 2593 1013 2606
rect 994 2573 1021 2576
rect 994 2526 997 2536
rect 1018 2533 1021 2573
rect 1038 2566 1041 2673
rect 1026 2563 1041 2566
rect 994 2523 1021 2526
rect 994 2513 1021 2516
rect 986 2503 1005 2506
rect 970 2493 977 2496
rect 974 2436 977 2493
rect 974 2433 981 2436
rect 954 2423 965 2426
rect 954 2403 957 2423
rect 962 2413 973 2416
rect 978 2413 981 2433
rect 962 2403 973 2406
rect 986 2403 989 2446
rect 994 2413 997 2476
rect 930 2383 949 2386
rect 922 2373 933 2376
rect 874 2303 885 2306
rect 874 2233 877 2303
rect 882 2226 885 2276
rect 874 2223 885 2226
rect 874 2183 877 2223
rect 890 2216 893 2336
rect 906 2333 909 2356
rect 930 2286 933 2373
rect 914 2283 933 2286
rect 898 2223 909 2226
rect 882 2213 893 2216
rect 866 2173 877 2176
rect 858 2136 861 2156
rect 858 2133 869 2136
rect 874 2126 877 2173
rect 866 2123 877 2126
rect 858 2103 861 2116
rect 866 2096 869 2123
rect 882 2116 885 2213
rect 890 2203 901 2206
rect 890 2123 893 2186
rect 858 2093 869 2096
rect 730 1853 749 1856
rect 714 1843 721 1846
rect 658 1613 661 1636
rect 690 1603 693 1626
rect 698 1613 701 1666
rect 590 1483 597 1486
rect 594 1446 597 1483
rect 610 1483 617 1486
rect 634 1513 641 1516
rect 594 1443 601 1446
rect 554 1433 573 1436
rect 554 1366 557 1433
rect 570 1393 573 1406
rect 598 1396 601 1443
rect 594 1393 601 1396
rect 554 1363 573 1366
rect 526 1353 533 1356
rect 474 1213 477 1353
rect 482 1306 485 1346
rect 490 1333 501 1336
rect 506 1326 509 1336
rect 514 1333 525 1336
rect 482 1303 489 1306
rect 486 1206 489 1303
rect 498 1233 501 1326
rect 506 1323 517 1326
rect 522 1283 525 1333
rect 530 1276 533 1353
rect 546 1313 549 1336
rect 514 1273 533 1276
rect 482 1203 489 1206
rect 442 1153 453 1156
rect 450 1086 453 1153
rect 474 1123 477 1146
rect 450 1083 469 1086
rect 482 1083 485 1203
rect 434 1013 453 1016
rect 426 993 429 1006
rect 410 933 413 946
rect 426 933 429 966
rect 386 873 397 876
rect 378 803 381 826
rect 386 803 389 873
rect 394 796 397 856
rect 410 853 413 926
rect 418 906 421 926
rect 442 923 445 1006
rect 450 986 453 1013
rect 466 1003 469 1083
rect 490 996 493 1176
rect 498 1076 501 1206
rect 514 1166 517 1273
rect 530 1213 533 1266
rect 522 1193 525 1206
rect 538 1203 541 1286
rect 546 1276 549 1306
rect 546 1273 557 1276
rect 554 1216 557 1273
rect 546 1213 557 1216
rect 570 1213 573 1363
rect 578 1323 581 1336
rect 586 1273 589 1316
rect 546 1196 549 1213
rect 530 1193 549 1196
rect 514 1163 521 1166
rect 518 1076 521 1163
rect 498 1073 505 1076
rect 502 1026 505 1073
rect 514 1073 521 1076
rect 514 1053 517 1073
rect 530 1056 533 1193
rect 538 1123 541 1136
rect 554 1106 557 1196
rect 586 1193 589 1216
rect 594 1203 597 1393
rect 602 1203 605 1236
rect 546 1103 557 1106
rect 530 1053 537 1056
rect 502 1023 509 1026
rect 482 993 493 996
rect 450 983 469 986
rect 450 906 453 936
rect 418 903 429 906
rect 426 856 429 903
rect 418 853 429 856
rect 442 903 453 906
rect 378 793 397 796
rect 354 733 365 736
rect 370 713 373 726
rect 378 693 381 793
rect 298 593 309 596
rect 314 593 325 596
rect 298 533 301 593
rect 314 533 317 593
rect 290 403 293 426
rect 298 386 301 456
rect 322 426 325 526
rect 338 503 341 636
rect 346 533 349 606
rect 354 533 357 606
rect 370 533 373 636
rect 378 563 381 616
rect 386 603 389 746
rect 394 733 397 786
rect 402 706 405 776
rect 410 723 413 806
rect 418 803 421 853
rect 442 836 445 903
rect 458 876 461 936
rect 466 896 469 983
rect 474 906 477 936
rect 482 913 485 993
rect 498 953 501 1016
rect 498 906 501 946
rect 506 943 509 1023
rect 534 976 537 1053
rect 546 1036 549 1103
rect 546 1033 557 1036
rect 546 993 549 1016
rect 530 973 537 976
rect 530 946 533 973
rect 554 946 557 1033
rect 562 953 565 1136
rect 570 1046 573 1176
rect 610 1173 613 1483
rect 618 1413 621 1426
rect 618 1303 621 1376
rect 626 1226 629 1326
rect 634 1233 637 1513
rect 642 1373 645 1396
rect 642 1313 645 1336
rect 650 1296 653 1536
rect 666 1533 669 1576
rect 706 1443 709 1526
rect 714 1436 717 1843
rect 722 1803 725 1826
rect 730 1813 741 1816
rect 722 1723 725 1736
rect 730 1706 733 1796
rect 726 1703 733 1706
rect 726 1656 729 1703
rect 738 1663 741 1813
rect 746 1793 749 1853
rect 770 1853 813 1856
rect 770 1803 773 1853
rect 826 1836 829 1926
rect 834 1843 837 1926
rect 802 1803 805 1836
rect 826 1833 837 1836
rect 826 1813 829 1826
rect 746 1706 749 1766
rect 746 1703 757 1706
rect 726 1653 733 1656
rect 730 1566 733 1653
rect 746 1603 749 1616
rect 730 1563 741 1566
rect 754 1563 757 1703
rect 762 1676 765 1776
rect 834 1753 837 1833
rect 842 1776 845 2066
rect 858 2036 861 2093
rect 874 2063 877 2116
rect 882 2113 893 2116
rect 850 2033 861 2036
rect 850 2003 853 2033
rect 858 1993 861 2016
rect 866 1983 869 2006
rect 874 1976 877 2016
rect 882 2003 885 2056
rect 850 1923 853 1956
rect 858 1933 861 1976
rect 866 1973 877 1976
rect 850 1783 853 1886
rect 866 1873 869 1973
rect 842 1773 861 1776
rect 850 1733 853 1756
rect 786 1703 789 1726
rect 834 1723 845 1726
rect 762 1673 773 1676
rect 770 1576 773 1673
rect 818 1613 821 1626
rect 762 1573 773 1576
rect 738 1506 741 1563
rect 762 1553 765 1573
rect 794 1556 797 1606
rect 786 1553 797 1556
rect 730 1503 741 1506
rect 682 1433 717 1436
rect 658 1303 661 1406
rect 674 1333 677 1416
rect 682 1366 685 1433
rect 690 1376 693 1416
rect 698 1383 701 1416
rect 706 1403 709 1426
rect 722 1416 725 1466
rect 714 1413 725 1416
rect 722 1376 725 1406
rect 690 1373 725 1376
rect 682 1363 717 1366
rect 674 1316 677 1326
rect 682 1323 685 1336
rect 690 1333 693 1346
rect 698 1323 701 1336
rect 706 1316 709 1336
rect 646 1293 653 1296
rect 646 1236 649 1293
rect 646 1233 653 1236
rect 618 1223 629 1226
rect 618 1213 621 1223
rect 634 1213 645 1216
rect 626 1193 629 1206
rect 578 1133 581 1146
rect 594 1133 597 1156
rect 586 1086 589 1126
rect 586 1083 597 1086
rect 570 1043 581 1046
rect 570 986 573 1036
rect 578 1013 581 1043
rect 594 1013 597 1083
rect 586 993 589 1006
rect 570 983 589 986
rect 586 953 589 983
rect 526 943 533 946
rect 474 903 501 906
rect 466 893 477 896
rect 458 873 469 876
rect 442 833 453 836
rect 450 816 453 833
rect 458 823 461 866
rect 466 843 469 873
rect 434 736 437 816
rect 418 716 421 736
rect 426 733 437 736
rect 442 736 445 816
rect 450 813 469 816
rect 450 803 461 806
rect 466 793 469 813
rect 466 773 469 786
rect 474 746 477 893
rect 482 813 485 856
rect 458 743 477 746
rect 442 733 453 736
rect 458 726 461 743
rect 426 723 461 726
rect 466 733 477 736
rect 418 713 445 716
rect 450 706 453 716
rect 402 703 417 706
rect 294 383 301 386
rect 306 423 325 426
rect 294 286 297 383
rect 306 343 309 423
rect 314 383 317 416
rect 338 413 341 436
rect 362 413 365 526
rect 378 453 381 536
rect 386 533 389 546
rect 394 516 397 626
rect 390 513 397 516
rect 370 406 373 416
rect 330 366 333 406
rect 362 403 373 406
rect 378 403 381 426
rect 362 376 365 403
rect 314 363 333 366
rect 354 373 365 376
rect 274 283 297 286
rect 258 166 261 206
rect 266 203 269 216
rect 218 163 261 166
rect 170 133 173 146
rect 218 123 221 163
rect 274 123 277 283
rect 290 256 293 276
rect 290 253 297 256
rect 282 203 285 226
rect 294 196 297 253
rect 290 193 297 196
rect 290 143 293 193
rect 306 123 309 326
rect 314 323 317 363
rect 330 286 333 346
rect 354 323 357 373
rect 390 366 393 513
rect 366 363 393 366
rect 366 316 369 363
rect 402 343 405 696
rect 414 626 417 703
rect 426 703 453 706
rect 414 623 421 626
rect 410 533 413 606
rect 418 603 421 623
rect 426 576 429 703
rect 418 573 429 576
rect 418 513 421 573
rect 418 413 421 436
rect 386 323 389 336
rect 410 323 413 406
rect 426 403 429 566
rect 434 523 437 666
rect 442 583 445 606
rect 450 593 453 606
rect 458 563 461 676
rect 466 556 469 733
rect 474 633 477 726
rect 474 596 477 616
rect 482 603 485 796
rect 490 733 493 806
rect 498 793 501 806
rect 506 786 509 816
rect 514 803 517 936
rect 526 816 529 943
rect 538 903 541 936
rect 538 826 541 896
rect 546 863 549 946
rect 554 943 589 946
rect 554 913 557 936
rect 562 923 573 926
rect 578 923 581 936
rect 538 823 549 826
rect 554 823 557 896
rect 586 893 589 943
rect 594 846 597 936
rect 602 916 605 1146
rect 610 1116 613 1136
rect 610 1113 617 1116
rect 614 1026 617 1113
rect 610 1023 617 1026
rect 610 1003 613 1023
rect 626 1003 629 1176
rect 634 1106 637 1206
rect 642 1156 645 1213
rect 650 1173 653 1233
rect 658 1166 661 1286
rect 666 1213 669 1316
rect 674 1313 709 1316
rect 666 1173 669 1206
rect 658 1163 669 1166
rect 642 1153 661 1156
rect 642 1123 645 1146
rect 634 1103 645 1106
rect 642 1036 645 1103
rect 634 1033 645 1036
rect 610 923 613 946
rect 602 913 613 916
rect 562 843 597 846
rect 526 813 533 816
rect 514 793 525 796
rect 530 786 533 813
rect 506 783 533 786
rect 506 736 509 783
rect 538 743 541 816
rect 506 733 517 736
rect 490 613 493 686
rect 506 613 509 726
rect 514 673 517 733
rect 522 703 525 726
rect 530 723 541 726
rect 546 696 549 823
rect 554 803 557 816
rect 522 693 549 696
rect 474 593 493 596
rect 450 553 469 556
rect 434 503 437 516
rect 442 433 445 536
rect 442 386 445 406
rect 450 386 453 553
rect 458 403 461 536
rect 474 533 477 546
rect 490 533 493 593
rect 498 573 501 606
rect 506 566 509 606
rect 498 563 509 566
rect 498 533 501 563
rect 466 443 469 526
rect 482 433 485 526
rect 498 453 501 526
rect 514 436 517 616
rect 522 603 525 693
rect 530 586 533 686
rect 526 583 533 586
rect 526 496 529 583
rect 538 573 541 636
rect 546 603 549 676
rect 538 503 541 566
rect 554 546 557 736
rect 562 683 565 843
rect 570 753 573 816
rect 586 813 589 836
rect 594 786 597 806
rect 590 783 597 786
rect 570 626 573 736
rect 590 726 593 783
rect 602 743 605 876
rect 610 733 613 913
rect 618 896 621 996
rect 626 913 629 926
rect 618 893 625 896
rect 622 826 625 893
rect 618 823 625 826
rect 618 746 621 823
rect 634 813 637 1033
rect 658 1023 661 1153
rect 666 1143 669 1163
rect 666 1123 669 1136
rect 674 1133 677 1196
rect 690 1193 693 1276
rect 690 1046 693 1126
rect 698 1123 701 1176
rect 706 1133 709 1156
rect 714 1116 717 1363
rect 722 1213 725 1346
rect 722 1123 725 1176
rect 730 1166 733 1503
rect 738 1423 741 1486
rect 762 1446 765 1536
rect 778 1476 781 1526
rect 786 1493 789 1553
rect 802 1533 805 1556
rect 826 1546 829 1666
rect 858 1606 861 1773
rect 866 1653 869 1826
rect 874 1773 877 1966
rect 874 1723 877 1756
rect 882 1706 885 1996
rect 890 1993 893 2113
rect 898 2096 901 2136
rect 906 2113 909 2206
rect 914 2133 917 2283
rect 922 2153 925 2206
rect 930 2203 933 2216
rect 938 2203 941 2366
rect 946 2196 949 2383
rect 962 2366 965 2403
rect 954 2363 965 2366
rect 954 2323 957 2363
rect 954 2203 957 2236
rect 962 2203 965 2246
rect 970 2203 973 2346
rect 986 2323 989 2366
rect 978 2213 981 2256
rect 994 2226 997 2406
rect 986 2223 997 2226
rect 1002 2306 1005 2503
rect 1010 2383 1013 2506
rect 1026 2496 1029 2563
rect 1050 2556 1053 2783
rect 1074 2766 1077 2883
rect 1090 2873 1093 2926
rect 1098 2923 1105 2926
rect 1102 2866 1105 2923
rect 1122 2913 1125 2936
rect 1146 2883 1149 2926
rect 1158 2906 1161 3003
rect 1158 2903 1165 2906
rect 1162 2883 1165 2903
rect 1098 2863 1105 2866
rect 1066 2763 1077 2766
rect 1058 2703 1061 2726
rect 1066 2673 1069 2763
rect 1082 2713 1085 2796
rect 1090 2766 1093 2826
rect 1098 2813 1101 2863
rect 1090 2763 1109 2766
rect 1082 2666 1085 2706
rect 1106 2673 1109 2763
rect 1082 2663 1109 2666
rect 1058 2566 1061 2616
rect 1058 2563 1069 2566
rect 1034 2553 1053 2556
rect 1066 2553 1069 2563
rect 1034 2513 1037 2553
rect 1050 2523 1053 2536
rect 1022 2493 1029 2496
rect 1022 2416 1025 2493
rect 1018 2413 1025 2416
rect 1018 2343 1021 2413
rect 1026 2376 1029 2406
rect 1034 2383 1037 2506
rect 1042 2423 1045 2476
rect 1042 2376 1045 2406
rect 1026 2373 1045 2376
rect 1050 2356 1053 2516
rect 1074 2503 1077 2646
rect 1082 2476 1085 2656
rect 1090 2573 1093 2616
rect 1098 2566 1101 2636
rect 1106 2593 1109 2663
rect 1066 2473 1085 2476
rect 1090 2563 1101 2566
rect 1090 2473 1093 2563
rect 1098 2523 1101 2536
rect 1066 2406 1069 2473
rect 1098 2466 1101 2516
rect 1074 2463 1101 2466
rect 1074 2413 1077 2463
rect 1106 2456 1109 2466
rect 1082 2453 1109 2456
rect 1082 2416 1085 2453
rect 1114 2446 1117 2866
rect 1122 2683 1125 2786
rect 1130 2763 1141 2766
rect 1130 2723 1133 2763
rect 1130 2686 1133 2716
rect 1130 2683 1141 2686
rect 1146 2676 1149 2806
rect 1138 2673 1149 2676
rect 1138 2626 1141 2673
rect 1154 2666 1157 2876
rect 1162 2813 1165 2826
rect 1162 2703 1165 2726
rect 1130 2623 1141 2626
rect 1146 2663 1157 2666
rect 1090 2423 1093 2446
rect 1098 2443 1117 2446
rect 1122 2446 1125 2606
rect 1130 2586 1133 2623
rect 1138 2606 1141 2616
rect 1146 2613 1149 2663
rect 1154 2613 1157 2656
rect 1162 2616 1165 2696
rect 1170 2626 1173 3006
rect 1178 2966 1181 3116
rect 1202 3096 1205 3176
rect 1194 3093 1205 3096
rect 1186 3013 1189 3046
rect 1178 2963 1189 2966
rect 1186 2933 1189 2963
rect 1194 2926 1197 3093
rect 1210 3026 1213 3246
rect 1218 3236 1221 3253
rect 1234 3243 1237 3373
rect 1218 3233 1225 3236
rect 1222 3176 1225 3233
rect 1218 3173 1225 3176
rect 1218 3053 1221 3173
rect 1226 3123 1229 3156
rect 1202 3016 1205 3026
rect 1210 3023 1221 3026
rect 1234 3023 1237 3076
rect 1202 3013 1213 3016
rect 1218 3006 1221 3023
rect 1210 2963 1213 3006
rect 1218 3003 1237 3006
rect 1242 2993 1245 3446
rect 1250 3323 1253 3416
rect 1258 3383 1261 3416
rect 1266 3333 1269 3453
rect 1274 3436 1277 3536
rect 1310 3506 1313 3563
rect 1322 3513 1325 3526
rect 1310 3503 1317 3506
rect 1274 3433 1293 3436
rect 1290 3403 1293 3433
rect 1314 3396 1317 3503
rect 1338 3436 1341 3556
rect 1346 3516 1349 3603
rect 1354 3523 1357 3576
rect 1346 3513 1353 3516
rect 1350 3466 1353 3513
rect 1350 3463 1357 3466
rect 1306 3393 1317 3396
rect 1330 3433 1341 3436
rect 1330 3396 1333 3433
rect 1338 3403 1341 3416
rect 1330 3393 1341 3396
rect 1282 3346 1285 3376
rect 1282 3343 1293 3346
rect 1250 3176 1253 3316
rect 1266 3263 1269 3326
rect 1274 3323 1293 3326
rect 1274 3223 1277 3323
rect 1298 3316 1301 3376
rect 1282 3313 1301 3316
rect 1306 3313 1309 3393
rect 1314 3333 1317 3366
rect 1258 3196 1261 3216
rect 1266 3213 1277 3216
rect 1282 3206 1285 3313
rect 1290 3213 1293 3296
rect 1298 3213 1301 3266
rect 1266 3203 1277 3206
rect 1282 3203 1301 3206
rect 1306 3196 1309 3286
rect 1314 3226 1317 3326
rect 1322 3283 1325 3326
rect 1330 3303 1333 3336
rect 1338 3323 1341 3393
rect 1354 3353 1357 3463
rect 1362 3426 1365 3606
rect 1370 3533 1373 3606
rect 1378 3436 1381 3536
rect 1386 3443 1389 3613
rect 1402 3603 1405 3613
rect 1410 3593 1413 3606
rect 1394 3493 1397 3516
rect 1402 3483 1405 3586
rect 1418 3583 1421 3606
rect 1410 3533 1421 3536
rect 1426 3513 1429 3526
rect 1378 3433 1389 3436
rect 1362 3423 1381 3426
rect 1370 3373 1373 3416
rect 1378 3363 1381 3423
rect 1362 3323 1365 3336
rect 1370 3303 1373 3326
rect 1378 3283 1381 3336
rect 1386 3326 1389 3433
rect 1418 3423 1421 3446
rect 1394 3366 1397 3416
rect 1402 3403 1413 3406
rect 1426 3376 1429 3426
rect 1434 3413 1437 3726
rect 1442 3673 1445 3733
rect 1442 3623 1445 3636
rect 1466 3626 1469 3753
rect 1522 3746 1525 3836
rect 1474 3743 1501 3746
rect 1482 3733 1493 3736
rect 1482 3723 1485 3733
rect 1466 3623 1477 3626
rect 1466 3593 1469 3606
rect 1474 3586 1477 3623
rect 1482 3593 1485 3626
rect 1490 3613 1493 3726
rect 1498 3723 1501 3743
rect 1514 3743 1525 3746
rect 1514 3733 1517 3743
rect 1538 3736 1541 3893
rect 1562 3883 1565 3926
rect 1546 3803 1549 3826
rect 1578 3806 1581 3946
rect 1602 3933 1605 4133
rect 1618 4096 1621 4146
rect 1614 4093 1621 4096
rect 1614 4036 1617 4093
rect 1650 4066 1653 4206
rect 1674 4193 1677 4216
rect 1666 4106 1669 4126
rect 1626 4063 1653 4066
rect 1614 4033 1621 4036
rect 1610 3996 1613 4016
rect 1618 4013 1621 4033
rect 1626 4003 1629 4063
rect 1634 4003 1637 4056
rect 1650 4053 1653 4063
rect 1662 4103 1669 4106
rect 1642 4003 1653 4006
rect 1610 3993 1637 3996
rect 1610 3853 1613 3926
rect 1618 3833 1621 3986
rect 1634 3923 1637 3993
rect 1586 3823 1613 3826
rect 1586 3813 1589 3823
rect 1554 3803 1581 3806
rect 1522 3733 1541 3736
rect 1554 3733 1557 3803
rect 1554 3716 1557 3726
rect 1562 3723 1565 3756
rect 1570 3733 1573 3796
rect 1594 3793 1597 3816
rect 1602 3813 1605 3823
rect 1610 3813 1613 3823
rect 1618 3813 1629 3816
rect 1602 3773 1605 3806
rect 1618 3803 1621 3813
rect 1634 3806 1637 3896
rect 1626 3803 1637 3806
rect 1642 3803 1645 4003
rect 1662 3966 1665 4103
rect 1682 4086 1685 4323
rect 1690 4216 1693 4236
rect 1690 4213 1697 4216
rect 1674 4083 1685 4086
rect 1674 3983 1677 4083
rect 1694 4066 1697 4213
rect 1714 4176 1717 4340
rect 1730 4326 1733 4340
rect 1786 4326 1789 4340
rect 1730 4323 1741 4326
rect 1738 4236 1741 4323
rect 1730 4233 1741 4236
rect 1762 4323 1789 4326
rect 1706 4173 1717 4176
rect 1706 4096 1709 4173
rect 1714 4123 1717 4136
rect 1722 4126 1725 4226
rect 1730 4213 1733 4233
rect 1738 4183 1741 4196
rect 1746 4193 1749 4206
rect 1754 4176 1757 4216
rect 1730 4173 1757 4176
rect 1730 4133 1733 4173
rect 1762 4146 1765 4323
rect 1786 4223 1789 4256
rect 1770 4213 1789 4216
rect 1746 4133 1749 4146
rect 1762 4143 1773 4146
rect 1722 4123 1733 4126
rect 1730 4113 1733 4123
rect 1706 4093 1717 4096
rect 1690 4063 1697 4066
rect 1690 4043 1693 4063
rect 1682 4023 1709 4026
rect 1682 4013 1685 4023
rect 1690 3983 1693 4016
rect 1698 3993 1701 4006
rect 1662 3963 1669 3966
rect 1666 3946 1669 3963
rect 1706 3953 1709 4023
rect 1714 3993 1717 4093
rect 1762 4023 1765 4066
rect 1730 4013 1757 4016
rect 1666 3943 1725 3946
rect 1650 3933 1661 3936
rect 1674 3926 1677 3936
rect 1682 3933 1693 3936
rect 1650 3923 1661 3926
rect 1666 3903 1669 3926
rect 1674 3923 1685 3926
rect 1626 3793 1629 3803
rect 1594 3736 1597 3756
rect 1586 3726 1589 3736
rect 1594 3733 1605 3736
rect 1578 3716 1581 3726
rect 1586 3723 1597 3726
rect 1554 3713 1581 3716
rect 1442 3533 1445 3556
rect 1442 3403 1445 3436
rect 1426 3373 1437 3376
rect 1394 3363 1405 3366
rect 1394 3343 1397 3356
rect 1386 3323 1393 3326
rect 1390 3276 1393 3323
rect 1402 3296 1405 3363
rect 1426 3326 1429 3356
rect 1434 3333 1437 3373
rect 1418 3303 1421 3326
rect 1426 3323 1437 3326
rect 1442 3323 1445 3336
rect 1434 3313 1437 3323
rect 1402 3293 1437 3296
rect 1386 3273 1393 3276
rect 1314 3223 1341 3226
rect 1258 3193 1293 3196
rect 1250 3173 1257 3176
rect 1254 3056 1257 3173
rect 1266 3103 1269 3166
rect 1290 3146 1293 3193
rect 1298 3193 1309 3196
rect 1298 3153 1301 3193
rect 1314 3146 1317 3196
rect 1338 3163 1341 3223
rect 1290 3143 1317 3146
rect 1250 3053 1257 3056
rect 1250 2973 1253 3053
rect 1242 2943 1253 2946
rect 1258 2943 1261 3036
rect 1274 3033 1277 3126
rect 1266 3003 1277 3006
rect 1282 2966 1285 3016
rect 1290 3006 1293 3143
rect 1298 3073 1301 3136
rect 1306 3116 1309 3126
rect 1314 3123 1317 3143
rect 1322 3133 1325 3156
rect 1330 3153 1341 3156
rect 1330 3116 1333 3153
rect 1306 3113 1333 3116
rect 1306 3023 1309 3086
rect 1338 3036 1341 3136
rect 1346 3123 1349 3266
rect 1354 3223 1381 3226
rect 1354 3213 1357 3223
rect 1354 3173 1357 3206
rect 1362 3176 1365 3216
rect 1378 3193 1381 3206
rect 1362 3173 1373 3176
rect 1354 3133 1357 3156
rect 1386 3133 1389 3273
rect 1394 3146 1397 3166
rect 1402 3156 1405 3226
rect 1426 3203 1429 3216
rect 1434 3183 1437 3293
rect 1450 3256 1453 3586
rect 1474 3583 1485 3586
rect 1458 3533 1469 3536
rect 1474 3493 1477 3526
rect 1466 3423 1477 3426
rect 1458 3403 1461 3416
rect 1474 3373 1477 3406
rect 1482 3336 1485 3583
rect 1490 3553 1493 3606
rect 1490 3523 1493 3536
rect 1498 3533 1501 3686
rect 1506 3613 1509 3626
rect 1522 3613 1525 3656
rect 1530 3643 1541 3646
rect 1554 3643 1573 3646
rect 1530 3613 1533 3643
rect 1554 3636 1557 3643
rect 1538 3633 1557 3636
rect 1506 3603 1517 3606
rect 1490 3506 1493 3516
rect 1506 3513 1509 3526
rect 1514 3506 1517 3536
rect 1490 3503 1517 3506
rect 1490 3343 1493 3503
rect 1498 3403 1501 3416
rect 1514 3413 1517 3466
rect 1506 3373 1509 3406
rect 1522 3363 1525 3606
rect 1538 3603 1541 3633
rect 1482 3333 1501 3336
rect 1458 3296 1461 3326
rect 1482 3303 1485 3326
rect 1490 3313 1493 3326
rect 1490 3296 1493 3306
rect 1458 3293 1493 3296
rect 1446 3253 1453 3256
rect 1446 3186 1449 3253
rect 1446 3183 1453 3186
rect 1402 3153 1413 3156
rect 1394 3143 1405 3146
rect 1402 3116 1405 3143
rect 1394 3113 1405 3116
rect 1394 3066 1397 3113
rect 1394 3063 1405 3066
rect 1330 3033 1341 3036
rect 1290 3003 1301 3006
rect 1330 3003 1333 3033
rect 1354 3013 1357 3046
rect 1402 3043 1405 3063
rect 1270 2963 1285 2966
rect 1186 2923 1197 2926
rect 1178 2793 1181 2846
rect 1186 2803 1189 2923
rect 1202 2833 1205 2926
rect 1210 2886 1213 2936
rect 1226 2903 1229 2936
rect 1210 2883 1221 2886
rect 1194 2746 1197 2816
rect 1202 2793 1205 2826
rect 1210 2783 1213 2816
rect 1218 2766 1221 2883
rect 1186 2743 1197 2746
rect 1210 2763 1221 2766
rect 1178 2643 1181 2726
rect 1186 2716 1189 2743
rect 1194 2723 1197 2736
rect 1186 2713 1197 2716
rect 1202 2703 1205 2726
rect 1210 2696 1213 2763
rect 1218 2733 1221 2756
rect 1218 2713 1221 2726
rect 1226 2706 1229 2816
rect 1234 2803 1237 2826
rect 1234 2735 1237 2766
rect 1242 2736 1245 2886
rect 1250 2803 1253 2943
rect 1258 2763 1261 2926
rect 1270 2896 1273 2963
rect 1266 2893 1273 2896
rect 1266 2816 1269 2893
rect 1314 2876 1317 2926
rect 1322 2886 1325 2976
rect 1338 2903 1341 2936
rect 1322 2883 1349 2886
rect 1362 2883 1365 2936
rect 1274 2873 1301 2876
rect 1314 2873 1325 2876
rect 1274 2843 1277 2873
rect 1274 2823 1277 2836
rect 1266 2813 1277 2816
rect 1266 2793 1269 2806
rect 1274 2803 1277 2813
rect 1282 2776 1285 2816
rect 1290 2803 1293 2846
rect 1306 2803 1309 2826
rect 1314 2813 1317 2836
rect 1274 2773 1285 2776
rect 1242 2733 1253 2736
rect 1234 2723 1245 2726
rect 1226 2703 1233 2706
rect 1210 2693 1221 2696
rect 1170 2623 1189 2626
rect 1162 2613 1173 2616
rect 1138 2603 1165 2606
rect 1130 2583 1137 2586
rect 1134 2526 1137 2583
rect 1130 2523 1137 2526
rect 1130 2473 1133 2523
rect 1146 2516 1149 2576
rect 1154 2533 1157 2596
rect 1178 2593 1181 2606
rect 1186 2586 1189 2606
rect 1170 2583 1189 2586
rect 1146 2513 1153 2516
rect 1122 2443 1133 2446
rect 1082 2413 1093 2416
rect 1098 2413 1101 2443
rect 1106 2433 1125 2436
rect 1046 2353 1053 2356
rect 1018 2306 1021 2336
rect 1002 2303 1021 2306
rect 986 2206 989 2223
rect 978 2203 989 2206
rect 930 2193 949 2196
rect 898 2093 905 2096
rect 902 2016 905 2093
rect 902 2013 909 2016
rect 898 1936 901 2006
rect 906 1966 909 2013
rect 914 1983 917 2016
rect 906 1963 917 1966
rect 890 1933 901 1936
rect 906 1933 909 1946
rect 890 1903 893 1933
rect 878 1703 885 1706
rect 878 1636 881 1703
rect 878 1633 885 1636
rect 866 1613 877 1616
rect 858 1603 869 1606
rect 866 1566 869 1603
rect 866 1563 873 1566
rect 826 1543 837 1546
rect 834 1496 837 1543
rect 826 1493 837 1496
rect 778 1473 789 1476
rect 754 1443 765 1446
rect 738 1403 741 1416
rect 754 1396 757 1443
rect 770 1403 773 1436
rect 754 1393 765 1396
rect 762 1346 765 1393
rect 762 1343 773 1346
rect 746 1323 749 1336
rect 770 1316 773 1343
rect 778 1333 781 1466
rect 786 1403 789 1473
rect 786 1323 789 1346
rect 770 1313 789 1316
rect 738 1173 741 1306
rect 770 1213 773 1236
rect 778 1213 781 1256
rect 786 1206 789 1313
rect 778 1203 789 1206
rect 730 1163 737 1166
rect 714 1113 725 1116
rect 666 1043 693 1046
rect 650 993 653 1016
rect 642 923 645 936
rect 650 906 653 926
rect 646 903 653 906
rect 646 826 649 903
rect 658 843 661 936
rect 666 916 669 1043
rect 682 1026 685 1036
rect 682 1023 701 1026
rect 706 1023 709 1046
rect 674 1013 693 1016
rect 666 913 673 916
rect 670 856 673 913
rect 682 906 685 936
rect 690 923 693 1013
rect 698 963 701 1023
rect 706 973 709 1006
rect 722 983 725 1113
rect 734 1036 737 1163
rect 746 1133 749 1146
rect 734 1033 741 1036
rect 738 1013 741 1033
rect 730 993 733 1006
rect 746 1003 749 1116
rect 754 1106 757 1126
rect 762 1123 765 1136
rect 778 1123 781 1203
rect 786 1113 789 1126
rect 794 1116 797 1466
rect 802 1406 805 1416
rect 810 1413 813 1446
rect 802 1403 821 1406
rect 818 1383 821 1403
rect 810 1346 813 1366
rect 810 1343 817 1346
rect 814 1286 817 1343
rect 810 1283 817 1286
rect 826 1283 829 1493
rect 834 1396 837 1436
rect 842 1403 845 1416
rect 850 1403 853 1526
rect 870 1486 873 1563
rect 866 1483 873 1486
rect 866 1456 869 1483
rect 866 1453 873 1456
rect 834 1393 853 1396
rect 834 1333 837 1386
rect 802 1133 805 1206
rect 794 1113 801 1116
rect 754 1103 761 1106
rect 758 996 761 1103
rect 754 993 761 996
rect 714 933 717 966
rect 754 956 757 993
rect 682 903 697 906
rect 706 903 717 906
rect 670 853 677 856
rect 646 823 653 826
rect 658 823 661 836
rect 650 806 653 823
rect 666 813 669 836
rect 674 823 677 853
rect 682 816 685 896
rect 694 836 697 903
rect 694 833 701 836
rect 698 816 701 833
rect 706 823 709 896
rect 674 813 685 816
rect 626 803 653 806
rect 674 803 677 813
rect 650 756 653 803
rect 650 753 657 756
rect 618 743 645 746
rect 618 726 621 736
rect 642 733 645 743
rect 578 713 581 726
rect 586 723 593 726
rect 586 696 589 723
rect 594 703 597 716
rect 602 713 605 726
rect 578 693 589 696
rect 578 663 581 693
rect 562 623 573 626
rect 562 566 565 623
rect 570 613 581 616
rect 586 613 589 686
rect 610 626 613 726
rect 618 723 645 726
rect 642 683 645 716
rect 654 666 657 753
rect 650 663 657 666
rect 666 663 669 746
rect 650 636 653 663
rect 634 633 653 636
rect 594 603 597 626
rect 610 623 629 626
rect 610 613 613 623
rect 562 563 605 566
rect 546 543 557 546
rect 546 533 549 543
rect 526 493 533 496
rect 530 446 533 493
rect 530 443 549 446
rect 442 383 469 386
rect 322 283 333 286
rect 362 313 369 316
rect 322 203 325 283
rect 362 216 365 313
rect 330 213 341 216
rect 346 213 365 216
rect 330 123 333 206
rect 346 203 349 213
rect 354 196 357 206
rect 370 203 373 226
rect 394 213 397 246
rect 402 203 405 226
rect 410 213 421 216
rect 442 203 445 236
rect 458 203 461 326
rect 466 323 469 383
rect 474 366 477 416
rect 498 413 501 436
rect 506 433 517 436
rect 506 416 509 433
rect 506 413 517 416
rect 490 383 493 406
rect 474 363 485 366
rect 482 316 485 363
rect 530 343 533 406
rect 506 323 509 336
rect 538 323 541 386
rect 474 313 485 316
rect 474 243 477 313
rect 546 306 549 443
rect 538 303 549 306
rect 538 256 541 303
rect 538 253 549 256
rect 546 233 549 253
rect 482 213 485 226
rect 354 193 389 196
rect 386 123 389 193
rect 426 133 429 146
rect 474 123 477 146
rect 530 133 533 166
rect 530 116 533 126
rect 538 123 541 196
rect 546 133 549 146
rect 554 123 557 536
rect 570 403 573 536
rect 594 523 597 546
rect 586 323 589 396
rect 602 316 605 563
rect 610 536 613 606
rect 618 593 621 616
rect 626 563 629 623
rect 634 576 637 633
rect 650 593 653 606
rect 634 573 641 576
rect 610 533 621 536
rect 638 516 641 573
rect 650 523 653 536
rect 638 513 645 516
rect 642 436 645 513
rect 642 433 653 436
rect 618 383 621 416
rect 650 413 653 433
rect 578 313 605 316
rect 578 236 581 313
rect 610 243 613 326
rect 618 306 621 346
rect 658 343 661 536
rect 666 523 669 556
rect 674 506 677 726
rect 682 696 685 736
rect 690 723 693 816
rect 698 813 709 816
rect 698 723 701 736
rect 706 696 709 813
rect 714 803 717 836
rect 714 723 717 746
rect 682 693 709 696
rect 714 693 717 716
rect 670 503 677 506
rect 670 416 673 503
rect 682 423 685 666
rect 690 533 693 616
rect 706 533 709 576
rect 698 503 701 526
rect 714 473 717 616
rect 722 593 725 956
rect 730 953 757 956
rect 730 823 733 953
rect 738 913 741 946
rect 746 843 749 926
rect 738 756 741 816
rect 754 803 757 936
rect 762 816 765 976
rect 770 943 773 1106
rect 770 913 773 936
rect 770 823 773 876
rect 762 813 773 816
rect 778 813 781 996
rect 786 986 789 1086
rect 798 1056 801 1113
rect 810 1093 813 1283
rect 818 1103 821 1216
rect 834 1213 837 1326
rect 842 1293 845 1326
rect 826 1106 829 1126
rect 834 1123 837 1206
rect 842 1203 845 1226
rect 826 1103 833 1106
rect 794 1053 801 1056
rect 794 1003 797 1053
rect 802 1033 813 1036
rect 802 1023 805 1033
rect 818 1023 821 1066
rect 802 993 805 1016
rect 786 983 813 986
rect 786 906 789 936
rect 794 923 797 946
rect 802 906 805 966
rect 810 933 813 983
rect 810 913 813 926
rect 786 903 793 906
rect 802 903 813 906
rect 818 903 821 1016
rect 830 956 833 1103
rect 842 1013 845 1136
rect 850 1123 853 1393
rect 858 1326 861 1446
rect 870 1386 873 1453
rect 866 1383 873 1386
rect 866 1363 869 1383
rect 866 1333 869 1346
rect 874 1326 877 1336
rect 858 1323 877 1326
rect 874 1246 877 1266
rect 866 1243 877 1246
rect 866 1156 869 1243
rect 866 1153 877 1156
rect 850 1023 853 1106
rect 826 953 833 956
rect 842 953 845 1006
rect 790 836 793 903
rect 786 833 793 836
rect 730 753 741 756
rect 730 716 733 753
rect 762 746 765 806
rect 746 743 765 746
rect 746 733 749 743
rect 746 723 757 726
rect 762 723 765 736
rect 746 716 749 723
rect 770 716 773 813
rect 730 713 749 716
rect 762 713 773 716
rect 738 613 741 626
rect 754 623 757 656
rect 746 573 749 616
rect 730 463 733 536
rect 754 446 757 616
rect 762 533 765 713
rect 770 613 773 686
rect 778 653 781 756
rect 786 646 789 833
rect 802 813 805 846
rect 810 766 813 903
rect 794 763 813 766
rect 794 733 797 763
rect 802 733 805 756
rect 802 703 805 726
rect 810 713 813 726
rect 778 643 789 646
rect 778 613 781 643
rect 786 613 789 636
rect 778 523 781 546
rect 670 413 677 416
rect 698 413 701 436
rect 706 413 709 446
rect 746 443 757 446
rect 794 446 797 656
rect 802 613 805 676
rect 802 586 805 606
rect 810 603 813 696
rect 802 583 809 586
rect 806 516 809 583
rect 802 513 809 516
rect 802 493 805 513
rect 794 443 801 446
rect 634 333 653 336
rect 618 303 629 306
rect 642 303 645 326
rect 562 213 565 236
rect 574 233 581 236
rect 574 186 577 233
rect 594 203 597 216
rect 574 183 581 186
rect 578 136 581 183
rect 562 126 565 136
rect 570 133 581 136
rect 562 123 573 126
rect 578 116 581 133
rect 530 113 581 116
rect 610 103 613 136
rect 626 133 629 303
rect 650 256 653 333
rect 666 323 669 336
rect 674 316 677 413
rect 698 356 701 406
rect 706 403 717 406
rect 706 383 709 403
rect 722 366 725 416
rect 730 403 733 436
rect 746 426 749 443
rect 742 423 749 426
rect 722 363 733 366
rect 670 313 677 316
rect 682 353 701 356
rect 642 253 653 256
rect 642 213 645 253
rect 626 113 629 126
rect 634 123 637 206
rect 658 176 661 306
rect 670 236 673 313
rect 650 173 661 176
rect 666 233 673 236
rect 642 133 645 146
rect 650 123 653 173
rect 658 113 661 136
rect 666 103 669 233
rect 674 156 677 216
rect 682 163 685 353
rect 722 336 725 356
rect 690 323 693 336
rect 714 333 725 336
rect 730 326 733 363
rect 742 346 745 423
rect 742 343 749 346
rect 698 306 701 326
rect 722 323 733 326
rect 746 323 749 343
rect 754 333 757 406
rect 770 383 773 406
rect 798 396 801 443
rect 794 393 801 396
rect 778 336 781 376
rect 770 333 781 336
rect 690 203 693 306
rect 698 303 709 306
rect 722 303 725 323
rect 778 303 781 333
rect 794 313 797 393
rect 810 353 813 416
rect 818 373 821 846
rect 826 823 829 953
rect 834 906 837 936
rect 842 923 845 946
rect 858 933 861 1136
rect 874 1106 877 1153
rect 882 1116 885 1633
rect 890 1236 893 1876
rect 898 1723 901 1926
rect 906 1883 909 1926
rect 914 1876 917 1963
rect 922 1923 925 2066
rect 930 2013 933 2193
rect 970 2186 973 2196
rect 938 2183 949 2186
rect 938 2143 941 2183
rect 938 2023 941 2136
rect 946 2063 949 2166
rect 954 2123 957 2186
rect 962 2183 973 2186
rect 954 2056 957 2076
rect 962 2063 965 2183
rect 946 2046 949 2056
rect 954 2053 965 2056
rect 946 2043 957 2046
rect 930 1993 933 2006
rect 938 1983 941 2016
rect 954 2013 957 2043
rect 946 2003 957 2006
rect 962 2003 965 2053
rect 970 2003 973 2096
rect 978 2023 981 2166
rect 994 2146 997 2216
rect 1002 2163 1005 2303
rect 1010 2233 1013 2266
rect 1046 2236 1049 2353
rect 1058 2343 1061 2406
rect 1066 2403 1085 2406
rect 1046 2233 1053 2236
rect 1010 2203 1013 2216
rect 1026 2213 1045 2216
rect 1002 2153 1013 2156
rect 994 2143 1005 2146
rect 1002 2086 1005 2143
rect 1010 2096 1013 2153
rect 1018 2133 1021 2206
rect 1026 2183 1029 2213
rect 1034 2166 1037 2206
rect 1026 2163 1037 2166
rect 1018 2103 1021 2126
rect 1010 2093 1021 2096
rect 1002 2083 1013 2086
rect 986 2016 989 2046
rect 978 2013 989 2016
rect 994 2016 997 2056
rect 994 2013 1005 2016
rect 930 1933 933 1976
rect 938 1923 941 1936
rect 906 1873 917 1876
rect 906 1633 909 1873
rect 914 1813 917 1866
rect 922 1823 925 1886
rect 922 1753 925 1816
rect 938 1766 941 1826
rect 930 1763 941 1766
rect 914 1733 917 1746
rect 914 1616 917 1706
rect 930 1696 933 1763
rect 938 1743 941 1756
rect 930 1693 941 1696
rect 910 1613 917 1616
rect 898 1563 901 1606
rect 898 1403 901 1556
rect 910 1546 913 1613
rect 922 1546 925 1656
rect 938 1623 941 1693
rect 938 1583 941 1606
rect 910 1543 917 1546
rect 922 1543 941 1546
rect 906 1503 909 1526
rect 906 1396 909 1446
rect 898 1393 909 1396
rect 898 1303 901 1393
rect 914 1376 917 1543
rect 922 1493 925 1536
rect 930 1513 933 1536
rect 938 1506 941 1543
rect 930 1503 941 1506
rect 930 1413 933 1503
rect 946 1426 949 1996
rect 954 1793 957 2003
rect 978 1983 981 2013
rect 1010 2006 1013 2083
rect 970 1946 973 1966
rect 970 1943 977 1946
rect 962 1826 965 1926
rect 974 1856 977 1943
rect 986 1883 989 1926
rect 970 1853 977 1856
rect 970 1833 973 1853
rect 962 1823 973 1826
rect 962 1803 965 1816
rect 970 1806 973 1823
rect 978 1813 981 1826
rect 970 1803 981 1806
rect 986 1803 989 1866
rect 954 1723 957 1746
rect 954 1593 957 1636
rect 962 1586 965 1796
rect 970 1596 973 1736
rect 978 1716 981 1803
rect 994 1753 997 2006
rect 1002 2003 1013 2006
rect 978 1713 985 1716
rect 982 1646 985 1713
rect 978 1643 985 1646
rect 978 1613 981 1643
rect 994 1633 997 1726
rect 986 1603 989 1626
rect 994 1596 997 1606
rect 970 1593 997 1596
rect 954 1583 965 1586
rect 954 1493 957 1583
rect 978 1526 981 1546
rect 978 1523 985 1526
rect 970 1446 973 1516
rect 962 1443 973 1446
rect 946 1423 953 1426
rect 910 1373 917 1376
rect 910 1276 913 1373
rect 910 1273 917 1276
rect 890 1233 901 1236
rect 890 1203 893 1226
rect 890 1133 893 1146
rect 898 1123 901 1233
rect 906 1203 909 1256
rect 906 1133 909 1186
rect 914 1153 917 1273
rect 922 1233 925 1406
rect 930 1323 933 1356
rect 922 1203 925 1226
rect 930 1203 933 1276
rect 938 1223 941 1416
rect 950 1366 953 1423
rect 962 1413 965 1443
rect 982 1436 985 1523
rect 994 1513 997 1536
rect 978 1433 985 1436
rect 962 1383 965 1406
rect 946 1363 953 1366
rect 946 1316 949 1363
rect 954 1333 957 1346
rect 962 1323 965 1336
rect 946 1313 953 1316
rect 950 1236 953 1313
rect 962 1253 965 1286
rect 946 1233 953 1236
rect 914 1133 917 1146
rect 906 1123 917 1126
rect 906 1116 909 1123
rect 882 1113 909 1116
rect 914 1106 917 1116
rect 866 1103 877 1106
rect 906 1103 917 1106
rect 866 1003 869 1103
rect 874 1093 885 1096
rect 882 1016 885 1093
rect 874 1013 885 1016
rect 890 1013 893 1096
rect 882 993 885 1006
rect 850 913 861 916
rect 866 906 869 926
rect 874 923 877 986
rect 834 903 869 906
rect 842 846 845 903
rect 882 886 885 916
rect 874 883 885 886
rect 842 843 849 846
rect 826 733 829 816
rect 834 783 837 836
rect 834 723 837 776
rect 846 756 849 843
rect 858 813 861 836
rect 874 806 877 883
rect 874 803 885 806
rect 858 786 861 796
rect 858 783 869 786
rect 842 753 849 756
rect 826 633 829 716
rect 826 623 837 626
rect 842 623 845 753
rect 850 733 869 736
rect 850 693 853 733
rect 850 633 853 686
rect 866 683 869 716
rect 874 713 877 766
rect 826 613 829 623
rect 826 556 829 596
rect 834 583 837 616
rect 842 586 845 606
rect 858 586 861 606
rect 842 583 861 586
rect 826 553 877 556
rect 826 523 829 553
rect 834 346 837 536
rect 850 533 853 546
rect 866 526 869 536
rect 874 533 877 553
rect 842 443 845 526
rect 858 506 861 526
rect 866 523 877 526
rect 882 523 885 803
rect 890 783 893 986
rect 898 973 901 1006
rect 906 933 909 1103
rect 922 1083 925 1196
rect 930 1153 941 1156
rect 930 1123 933 1136
rect 938 1133 941 1153
rect 930 1083 941 1086
rect 914 983 917 1016
rect 898 903 901 926
rect 854 503 861 506
rect 854 436 857 503
rect 854 433 861 436
rect 842 413 853 416
rect 842 403 845 413
rect 858 406 861 433
rect 850 403 861 406
rect 802 323 805 346
rect 810 343 837 346
rect 706 246 709 303
rect 802 286 805 306
rect 794 283 805 286
rect 698 243 709 246
rect 698 196 701 243
rect 722 203 725 216
rect 762 213 765 246
rect 794 236 797 283
rect 794 233 805 236
rect 802 213 805 233
rect 810 226 813 343
rect 818 293 821 326
rect 826 243 829 336
rect 842 333 845 346
rect 850 326 853 403
rect 866 386 869 486
rect 890 466 893 756
rect 898 723 901 856
rect 914 826 917 926
rect 922 913 925 1026
rect 930 973 933 1083
rect 946 1076 949 1233
rect 954 1203 957 1216
rect 954 1153 957 1196
rect 954 1123 957 1146
rect 962 1123 965 1236
rect 954 1113 965 1116
rect 938 1073 949 1076
rect 938 1006 941 1073
rect 946 1013 949 1026
rect 954 1023 957 1056
rect 962 1023 965 1113
rect 970 1016 973 1396
rect 978 1126 981 1433
rect 986 1383 989 1416
rect 994 1413 997 1496
rect 994 1393 997 1406
rect 1002 1356 1005 2003
rect 1010 1863 1013 1996
rect 1018 1943 1021 2093
rect 1026 1916 1029 2163
rect 1042 2133 1045 2206
rect 1034 2043 1037 2066
rect 1034 2003 1037 2036
rect 1042 1943 1045 2126
rect 1050 2073 1053 2233
rect 1058 2203 1061 2326
rect 1066 2136 1069 2376
rect 1082 2286 1085 2403
rect 1078 2283 1085 2286
rect 1090 2283 1093 2413
rect 1098 2313 1101 2406
rect 1106 2303 1109 2366
rect 1078 2226 1081 2283
rect 1098 2243 1109 2246
rect 1114 2236 1117 2426
rect 1122 2403 1125 2433
rect 1130 2403 1133 2443
rect 1138 2393 1141 2506
rect 1150 2436 1153 2513
rect 1146 2433 1153 2436
rect 1122 2333 1125 2386
rect 1138 2333 1141 2386
rect 1146 2363 1149 2433
rect 1154 2383 1157 2416
rect 1162 2356 1165 2526
rect 1146 2353 1165 2356
rect 1098 2233 1117 2236
rect 1074 2223 1081 2226
rect 1074 2203 1077 2223
rect 1090 2213 1093 2226
rect 1098 2196 1101 2233
rect 1122 2226 1125 2326
rect 1130 2306 1133 2326
rect 1146 2323 1149 2353
rect 1130 2303 1137 2306
rect 1074 2193 1101 2196
rect 1098 2156 1101 2186
rect 1106 2163 1109 2226
rect 1114 2223 1125 2226
rect 1066 2133 1073 2136
rect 1082 2133 1085 2156
rect 1098 2153 1109 2156
rect 1058 2066 1061 2126
rect 1070 2086 1073 2133
rect 1090 2123 1093 2136
rect 1098 2106 1101 2136
rect 1094 2103 1101 2106
rect 1070 2083 1085 2086
rect 1050 2063 1061 2066
rect 1050 2013 1053 2063
rect 1066 2013 1069 2036
rect 1034 1926 1037 1936
rect 1034 1923 1053 1926
rect 1010 1793 1013 1846
rect 1018 1786 1021 1916
rect 1026 1913 1037 1916
rect 1026 1823 1029 1876
rect 1026 1793 1029 1816
rect 1010 1783 1021 1786
rect 1010 1713 1013 1783
rect 1018 1693 1021 1746
rect 1010 1533 1013 1656
rect 1026 1626 1029 1786
rect 1034 1743 1037 1913
rect 1058 1906 1061 2006
rect 1074 2003 1077 2076
rect 1082 1996 1085 2083
rect 1094 2036 1097 2103
rect 1106 2053 1109 2153
rect 1114 2133 1117 2223
rect 1134 2176 1137 2303
rect 1154 2293 1157 2336
rect 1162 2236 1165 2326
rect 1146 2233 1165 2236
rect 1146 2183 1149 2233
rect 1170 2226 1173 2583
rect 1194 2576 1197 2676
rect 1210 2603 1213 2686
rect 1218 2673 1221 2693
rect 1230 2646 1233 2703
rect 1230 2643 1237 2646
rect 1242 2643 1245 2706
rect 1194 2573 1221 2576
rect 1178 2533 1181 2556
rect 1186 2533 1197 2536
rect 1178 2413 1181 2476
rect 1186 2463 1189 2526
rect 1202 2506 1205 2526
rect 1210 2513 1213 2536
rect 1218 2523 1221 2573
rect 1226 2566 1229 2596
rect 1234 2573 1237 2643
rect 1242 2586 1245 2616
rect 1250 2593 1253 2733
rect 1242 2583 1253 2586
rect 1226 2563 1237 2566
rect 1226 2533 1229 2556
rect 1226 2506 1229 2516
rect 1202 2503 1229 2506
rect 1194 2413 1197 2446
rect 1178 2396 1181 2406
rect 1186 2403 1197 2406
rect 1202 2403 1205 2476
rect 1210 2403 1213 2446
rect 1218 2396 1221 2466
rect 1234 2446 1237 2563
rect 1250 2533 1253 2583
rect 1258 2573 1261 2736
rect 1266 2733 1269 2756
rect 1274 2646 1277 2773
rect 1282 2733 1285 2766
rect 1298 2726 1301 2736
rect 1306 2733 1309 2796
rect 1282 2723 1293 2726
rect 1298 2723 1309 2726
rect 1290 2696 1293 2723
rect 1282 2693 1293 2696
rect 1282 2673 1285 2693
rect 1290 2656 1293 2686
rect 1290 2653 1301 2656
rect 1274 2643 1293 2646
rect 1298 2643 1301 2653
rect 1290 2626 1293 2643
rect 1290 2623 1301 2626
rect 1274 2613 1293 2616
rect 1266 2526 1269 2536
rect 1274 2533 1277 2613
rect 1258 2513 1261 2526
rect 1266 2523 1277 2526
rect 1242 2456 1245 2506
rect 1266 2486 1269 2523
rect 1258 2483 1269 2486
rect 1258 2463 1261 2483
rect 1282 2476 1285 2576
rect 1290 2533 1293 2556
rect 1266 2473 1285 2476
rect 1242 2453 1261 2456
rect 1234 2443 1253 2446
rect 1178 2393 1197 2396
rect 1178 2333 1181 2376
rect 1154 2223 1173 2226
rect 1134 2173 1157 2176
rect 1122 2086 1125 2166
rect 1130 2133 1133 2156
rect 1138 2123 1141 2166
rect 1146 2123 1149 2156
rect 1154 2116 1157 2173
rect 1150 2113 1157 2116
rect 1122 2083 1141 2086
rect 1050 1903 1061 1906
rect 1066 1993 1085 1996
rect 1090 2033 1097 2036
rect 1090 1993 1093 2033
rect 1106 2003 1109 2026
rect 1042 1813 1045 1826
rect 1042 1753 1045 1796
rect 1050 1793 1053 1903
rect 1058 1803 1061 1816
rect 1042 1733 1061 1736
rect 1058 1723 1061 1733
rect 1066 1716 1069 1993
rect 1074 1833 1077 1946
rect 1082 1883 1085 1936
rect 1074 1813 1085 1816
rect 1074 1763 1077 1806
rect 1042 1713 1069 1716
rect 1042 1646 1045 1713
rect 1042 1643 1053 1646
rect 1026 1623 1037 1626
rect 1018 1583 1021 1616
rect 1018 1533 1021 1556
rect 1034 1546 1037 1623
rect 1050 1603 1053 1643
rect 1058 1613 1061 1686
rect 1066 1586 1069 1606
rect 1026 1543 1037 1546
rect 1058 1583 1069 1586
rect 1026 1526 1029 1543
rect 1018 1513 1021 1526
rect 1026 1523 1037 1526
rect 1034 1513 1037 1523
rect 1058 1496 1061 1583
rect 1058 1493 1069 1496
rect 1010 1393 1013 1456
rect 1042 1413 1045 1476
rect 1050 1393 1053 1406
rect 1058 1376 1061 1396
rect 1054 1373 1061 1376
rect 998 1353 1005 1356
rect 986 1283 989 1336
rect 998 1236 1001 1353
rect 1018 1333 1021 1366
rect 1042 1323 1045 1346
rect 998 1233 1005 1236
rect 986 1183 989 1206
rect 986 1153 989 1176
rect 986 1133 989 1146
rect 978 1123 989 1126
rect 978 1083 981 1116
rect 954 1013 973 1016
rect 938 1003 949 1006
rect 922 853 925 906
rect 930 903 933 946
rect 906 803 909 826
rect 914 823 925 826
rect 914 753 917 816
rect 898 483 901 706
rect 906 693 909 736
rect 914 653 917 726
rect 922 663 925 823
rect 930 813 933 836
rect 938 803 941 966
rect 946 906 949 1003
rect 954 993 957 1013
rect 962 986 965 1006
rect 954 983 965 986
rect 970 983 973 1006
rect 978 993 981 1016
rect 954 926 957 983
rect 962 933 965 956
rect 954 923 965 926
rect 970 923 973 946
rect 946 903 953 906
rect 950 836 953 903
rect 946 833 953 836
rect 930 733 933 756
rect 930 713 941 716
rect 946 693 949 833
rect 954 686 957 816
rect 962 803 965 923
rect 978 883 981 936
rect 962 703 965 736
rect 938 683 957 686
rect 906 556 909 616
rect 930 603 933 676
rect 906 553 925 556
rect 906 523 909 536
rect 914 523 917 546
rect 922 533 925 553
rect 922 523 933 526
rect 874 463 893 466
rect 874 413 877 463
rect 866 383 885 386
rect 890 383 893 406
rect 914 396 917 416
rect 906 393 917 396
rect 834 323 853 326
rect 858 333 877 336
rect 858 323 861 333
rect 810 223 821 226
rect 690 193 701 196
rect 810 193 813 216
rect 818 203 821 223
rect 850 213 853 323
rect 858 213 869 216
rect 690 156 693 193
rect 674 153 693 156
rect 690 123 693 136
rect 714 123 717 146
rect 810 133 813 156
rect 770 103 773 126
rect 842 123 845 206
rect 858 203 861 213
rect 866 196 869 206
rect 882 196 885 383
rect 890 316 893 326
rect 898 323 901 336
rect 906 333 909 393
rect 922 326 925 523
rect 938 456 941 683
rect 946 553 949 666
rect 970 653 973 866
rect 978 783 981 806
rect 978 646 981 746
rect 986 736 989 1123
rect 994 1063 997 1216
rect 1002 1173 1005 1233
rect 1010 1213 1013 1286
rect 1018 1206 1021 1306
rect 1054 1276 1057 1373
rect 1054 1273 1061 1276
rect 1010 1203 1021 1206
rect 1026 1203 1029 1236
rect 1034 1223 1037 1266
rect 1034 1213 1045 1216
rect 1002 1123 1005 1166
rect 994 783 997 1006
rect 1002 916 1005 1086
rect 1010 1063 1013 1203
rect 1018 1096 1021 1166
rect 1026 1143 1029 1196
rect 1034 1183 1037 1213
rect 1026 1113 1029 1136
rect 1034 1116 1037 1176
rect 1042 1143 1045 1206
rect 1050 1203 1053 1256
rect 1050 1136 1053 1156
rect 1042 1133 1053 1136
rect 1042 1123 1053 1126
rect 1034 1113 1053 1116
rect 1018 1093 1045 1096
rect 1018 1023 1021 1086
rect 1026 1016 1029 1066
rect 1010 923 1013 1016
rect 1018 1013 1029 1016
rect 1034 1013 1037 1056
rect 1018 996 1021 1013
rect 1026 1003 1037 1006
rect 1018 993 1029 996
rect 1026 933 1029 993
rect 1034 973 1037 1003
rect 1042 983 1045 1093
rect 1050 1003 1053 1113
rect 1058 986 1061 1273
rect 1066 1003 1069 1493
rect 1074 1473 1077 1516
rect 1082 1493 1085 1796
rect 1090 1716 1093 1986
rect 1098 1933 1101 1976
rect 1106 1923 1109 1996
rect 1122 1926 1125 1976
rect 1114 1923 1125 1926
rect 1098 1733 1101 1906
rect 1106 1793 1109 1866
rect 1114 1823 1117 1923
rect 1130 1916 1133 2066
rect 1126 1913 1133 1916
rect 1126 1856 1129 1913
rect 1122 1853 1129 1856
rect 1114 1786 1117 1816
rect 1106 1783 1117 1786
rect 1106 1723 1109 1783
rect 1122 1776 1125 1853
rect 1114 1773 1125 1776
rect 1090 1713 1097 1716
rect 1094 1636 1097 1713
rect 1114 1676 1117 1773
rect 1130 1766 1133 1836
rect 1090 1633 1097 1636
rect 1106 1673 1117 1676
rect 1122 1763 1133 1766
rect 1090 1516 1093 1633
rect 1098 1563 1101 1616
rect 1106 1556 1109 1673
rect 1122 1603 1125 1763
rect 1138 1756 1141 2083
rect 1150 2036 1153 2113
rect 1162 2063 1165 2216
rect 1170 2196 1173 2223
rect 1178 2203 1181 2306
rect 1186 2203 1189 2386
rect 1170 2193 1189 2196
rect 1170 2073 1173 2186
rect 1186 2183 1189 2193
rect 1178 2063 1181 2136
rect 1146 2033 1153 2036
rect 1146 1906 1149 2033
rect 1154 1953 1157 2016
rect 1178 1993 1181 2036
rect 1186 1966 1189 2126
rect 1162 1963 1189 1966
rect 1194 1966 1197 2393
rect 1210 2393 1221 2396
rect 1226 2423 1245 2426
rect 1202 2303 1205 2336
rect 1210 2323 1213 2393
rect 1202 2123 1205 2286
rect 1218 2283 1221 2346
rect 1226 2276 1229 2423
rect 1234 2383 1237 2416
rect 1242 2413 1245 2423
rect 1242 2376 1245 2406
rect 1250 2396 1253 2443
rect 1258 2403 1261 2453
rect 1266 2413 1269 2473
rect 1274 2406 1277 2466
rect 1266 2403 1277 2406
rect 1250 2393 1261 2396
rect 1242 2373 1253 2376
rect 1234 2293 1237 2336
rect 1242 2326 1245 2366
rect 1250 2333 1253 2373
rect 1258 2363 1261 2393
rect 1266 2343 1269 2403
rect 1242 2323 1249 2326
rect 1210 2273 1229 2276
rect 1210 2163 1213 2273
rect 1218 2213 1221 2226
rect 1226 2213 1229 2266
rect 1246 2236 1249 2323
rect 1258 2263 1261 2326
rect 1266 2316 1269 2336
rect 1274 2323 1277 2386
rect 1282 2333 1285 2406
rect 1290 2383 1293 2526
rect 1290 2316 1293 2346
rect 1266 2313 1293 2316
rect 1298 2296 1301 2623
rect 1306 2593 1309 2686
rect 1306 2403 1309 2536
rect 1314 2413 1317 2806
rect 1322 2733 1325 2873
rect 1330 2813 1333 2856
rect 1338 2793 1341 2806
rect 1346 2803 1349 2883
rect 1370 2823 1373 2926
rect 1354 2803 1357 2816
rect 1362 2813 1373 2816
rect 1378 2806 1381 2906
rect 1386 2886 1389 2996
rect 1394 2966 1397 3006
rect 1410 3003 1413 3153
rect 1418 3133 1421 3166
rect 1418 3116 1421 3126
rect 1426 3123 1429 3176
rect 1450 3163 1453 3183
rect 1418 3113 1445 3116
rect 1450 3013 1453 3136
rect 1466 3133 1469 3226
rect 1482 3213 1485 3293
rect 1490 3283 1493 3293
rect 1394 2963 1409 2966
rect 1406 2906 1409 2963
rect 1406 2903 1413 2906
rect 1418 2903 1421 2926
rect 1434 2923 1437 2996
rect 1386 2883 1405 2886
rect 1362 2793 1365 2806
rect 1370 2803 1381 2806
rect 1370 2786 1373 2803
rect 1386 2793 1389 2816
rect 1402 2813 1405 2883
rect 1346 2783 1373 2786
rect 1322 2533 1325 2726
rect 1330 2633 1333 2726
rect 1330 2606 1333 2616
rect 1338 2613 1341 2716
rect 1346 2676 1349 2783
rect 1394 2776 1397 2806
rect 1354 2773 1397 2776
rect 1354 2713 1357 2773
rect 1362 2713 1365 2766
rect 1378 2723 1381 2736
rect 1410 2733 1413 2903
rect 1442 2836 1445 2936
rect 1450 2863 1453 2926
rect 1426 2833 1445 2836
rect 1362 2683 1365 2706
rect 1346 2673 1381 2676
rect 1346 2613 1349 2626
rect 1370 2616 1373 2636
rect 1378 2623 1381 2673
rect 1330 2603 1357 2606
rect 1330 2576 1333 2596
rect 1362 2583 1365 2616
rect 1370 2613 1389 2616
rect 1370 2593 1373 2606
rect 1330 2573 1357 2576
rect 1330 2533 1341 2536
rect 1322 2516 1325 2526
rect 1322 2513 1333 2516
rect 1338 2513 1341 2526
rect 1314 2396 1317 2406
rect 1306 2393 1317 2396
rect 1322 2396 1325 2506
rect 1330 2416 1333 2513
rect 1346 2506 1349 2566
rect 1342 2503 1349 2506
rect 1354 2503 1357 2573
rect 1342 2446 1345 2503
rect 1362 2486 1365 2576
rect 1378 2563 1381 2606
rect 1386 2596 1389 2613
rect 1394 2603 1397 2686
rect 1386 2593 1397 2596
rect 1386 2556 1389 2586
rect 1394 2573 1397 2593
rect 1402 2566 1405 2726
rect 1410 2593 1413 2726
rect 1370 2553 1389 2556
rect 1370 2533 1373 2553
rect 1338 2443 1345 2446
rect 1354 2483 1365 2486
rect 1338 2423 1341 2443
rect 1330 2413 1349 2416
rect 1330 2403 1341 2406
rect 1322 2393 1333 2396
rect 1306 2343 1309 2393
rect 1294 2293 1301 2296
rect 1246 2233 1253 2236
rect 1218 2196 1221 2206
rect 1226 2203 1237 2206
rect 1242 2203 1245 2216
rect 1218 2193 1245 2196
rect 1210 2103 1213 2136
rect 1226 2133 1229 2166
rect 1234 2133 1237 2186
rect 1242 2163 1245 2193
rect 1250 2183 1253 2233
rect 1258 2203 1261 2226
rect 1266 2196 1269 2286
rect 1258 2193 1269 2196
rect 1218 2116 1221 2126
rect 1218 2113 1237 2116
rect 1202 2023 1205 2056
rect 1210 2003 1213 2066
rect 1202 1973 1205 1986
rect 1194 1963 1205 1966
rect 1154 1923 1157 1936
rect 1146 1903 1157 1906
rect 1162 1836 1165 1963
rect 1170 1933 1173 1956
rect 1178 1923 1181 1946
rect 1202 1936 1205 1963
rect 1210 1953 1213 1996
rect 1218 1946 1221 2056
rect 1234 2046 1237 2113
rect 1242 2053 1245 2156
rect 1234 2043 1245 2046
rect 1186 1903 1189 1936
rect 1194 1933 1205 1936
rect 1210 1943 1221 1946
rect 1146 1833 1165 1836
rect 1146 1803 1149 1826
rect 1154 1823 1165 1826
rect 1154 1813 1157 1823
rect 1130 1753 1141 1756
rect 1130 1603 1133 1753
rect 1138 1643 1141 1726
rect 1146 1723 1149 1796
rect 1162 1793 1165 1816
rect 1154 1676 1157 1736
rect 1170 1726 1173 1876
rect 1178 1803 1181 1826
rect 1186 1803 1189 1826
rect 1194 1796 1197 1933
rect 1202 1896 1205 1926
rect 1210 1903 1213 1943
rect 1218 1923 1221 1936
rect 1226 1923 1229 2016
rect 1234 2003 1237 2026
rect 1242 2013 1245 2043
rect 1250 1973 1253 2126
rect 1258 2086 1261 2193
rect 1266 2113 1269 2186
rect 1274 2163 1277 2206
rect 1282 2153 1285 2246
rect 1294 2236 1297 2293
rect 1306 2243 1309 2336
rect 1314 2333 1317 2386
rect 1322 2333 1325 2376
rect 1322 2303 1325 2326
rect 1330 2286 1333 2393
rect 1338 2293 1341 2396
rect 1346 2286 1349 2413
rect 1354 2296 1357 2483
rect 1362 2403 1365 2416
rect 1370 2403 1373 2476
rect 1378 2443 1381 2536
rect 1386 2466 1389 2553
rect 1394 2563 1405 2566
rect 1394 2533 1397 2563
rect 1402 2513 1405 2536
rect 1410 2523 1413 2556
rect 1386 2463 1405 2466
rect 1386 2436 1389 2456
rect 1378 2433 1389 2436
rect 1362 2303 1365 2336
rect 1370 2323 1373 2366
rect 1378 2346 1381 2433
rect 1386 2403 1389 2426
rect 1386 2363 1389 2396
rect 1378 2343 1389 2346
rect 1378 2313 1381 2343
rect 1354 2293 1373 2296
rect 1326 2283 1333 2286
rect 1294 2233 1301 2236
rect 1298 2216 1301 2233
rect 1290 2213 1301 2216
rect 1290 2183 1293 2213
rect 1298 2146 1301 2206
rect 1306 2203 1309 2216
rect 1298 2143 1309 2146
rect 1282 2103 1285 2136
rect 1306 2123 1309 2143
rect 1258 2083 1269 2086
rect 1202 1893 1213 1896
rect 1178 1793 1197 1796
rect 1202 1793 1205 1886
rect 1178 1733 1181 1793
rect 1194 1783 1205 1786
rect 1170 1723 1189 1726
rect 1194 1703 1197 1736
rect 1202 1733 1205 1783
rect 1154 1673 1181 1676
rect 1146 1613 1149 1636
rect 1162 1613 1173 1616
rect 1098 1533 1101 1556
rect 1106 1553 1117 1556
rect 1090 1513 1097 1516
rect 1074 1393 1077 1416
rect 1082 1413 1085 1446
rect 1094 1436 1097 1513
rect 1090 1433 1097 1436
rect 1090 1336 1093 1433
rect 1098 1403 1101 1416
rect 1086 1333 1093 1336
rect 1086 1286 1089 1333
rect 1086 1283 1093 1286
rect 1098 1283 1101 1326
rect 1074 1213 1077 1226
rect 1074 1163 1077 1196
rect 1054 983 1061 986
rect 1018 923 1029 926
rect 1034 923 1037 946
rect 1002 913 1017 916
rect 1002 843 1005 906
rect 1014 836 1017 913
rect 1026 853 1029 923
rect 1042 896 1045 936
rect 1054 916 1057 983
rect 1054 913 1061 916
rect 1042 893 1053 896
rect 1014 833 1021 836
rect 1002 753 1005 816
rect 1010 793 1013 816
rect 1018 803 1021 833
rect 1026 813 1029 836
rect 1034 773 1037 806
rect 1042 803 1045 866
rect 1042 756 1045 786
rect 1034 753 1045 756
rect 986 733 997 736
rect 986 673 989 726
rect 1002 703 1005 726
rect 962 586 965 646
rect 978 643 993 646
rect 954 583 965 586
rect 954 516 957 583
rect 962 533 965 556
rect 978 533 981 596
rect 990 516 993 643
rect 1002 573 1005 616
rect 1002 523 1005 556
rect 954 513 965 516
rect 934 453 941 456
rect 934 396 937 453
rect 962 436 965 513
rect 958 433 965 436
rect 986 513 993 516
rect 986 436 989 513
rect 986 433 997 436
rect 934 393 941 396
rect 938 333 941 393
rect 958 376 961 433
rect 954 373 961 376
rect 970 373 973 416
rect 994 386 997 433
rect 1010 413 1013 736
rect 1018 733 1021 746
rect 1018 673 1021 726
rect 1034 636 1037 753
rect 1034 633 1045 636
rect 1042 593 1045 633
rect 1018 503 1021 536
rect 1034 533 1037 576
rect 1026 493 1029 526
rect 1034 523 1045 526
rect 1034 433 1037 523
rect 994 383 1005 386
rect 914 323 925 326
rect 914 316 917 323
rect 890 313 917 316
rect 890 203 893 216
rect 898 203 901 236
rect 914 213 917 313
rect 954 223 957 373
rect 978 333 981 356
rect 922 213 933 216
rect 906 196 909 206
rect 922 203 925 213
rect 930 203 941 206
rect 978 203 981 226
rect 866 193 893 196
rect 906 193 949 196
rect 890 123 893 193
rect 922 123 925 136
rect 946 123 949 193
rect 1002 123 1005 383
rect 1010 353 1013 406
rect 1050 393 1053 893
rect 1058 733 1061 913
rect 1066 886 1069 996
rect 1074 956 1077 1136
rect 1082 1076 1085 1236
rect 1090 1213 1093 1283
rect 1106 1236 1109 1546
rect 1114 1516 1117 1553
rect 1122 1523 1125 1556
rect 1114 1513 1125 1516
rect 1114 1413 1117 1496
rect 1122 1406 1125 1513
rect 1130 1486 1133 1596
rect 1138 1533 1141 1566
rect 1146 1553 1149 1586
rect 1154 1563 1157 1606
rect 1146 1526 1149 1546
rect 1146 1523 1153 1526
rect 1130 1483 1141 1486
rect 1130 1423 1133 1476
rect 1114 1403 1125 1406
rect 1114 1323 1117 1403
rect 1138 1366 1141 1483
rect 1150 1426 1153 1523
rect 1162 1443 1165 1606
rect 1170 1533 1173 1606
rect 1178 1516 1181 1673
rect 1194 1626 1197 1646
rect 1194 1623 1201 1626
rect 1174 1513 1181 1516
rect 1174 1436 1177 1513
rect 1174 1433 1181 1436
rect 1122 1363 1141 1366
rect 1146 1423 1153 1426
rect 1122 1236 1125 1363
rect 1130 1333 1133 1356
rect 1146 1346 1149 1423
rect 1170 1406 1173 1416
rect 1154 1403 1173 1406
rect 1138 1343 1149 1346
rect 1106 1233 1113 1236
rect 1122 1233 1133 1236
rect 1090 1126 1093 1206
rect 1098 1183 1101 1226
rect 1110 1176 1113 1233
rect 1122 1203 1125 1226
rect 1110 1173 1125 1176
rect 1122 1156 1125 1173
rect 1114 1153 1125 1156
rect 1106 1136 1109 1146
rect 1098 1133 1109 1136
rect 1090 1123 1107 1126
rect 1114 1083 1117 1153
rect 1082 1073 1093 1076
rect 1082 973 1085 1016
rect 1090 1013 1093 1073
rect 1122 1036 1125 1146
rect 1098 1033 1125 1036
rect 1090 963 1093 1006
rect 1074 953 1093 956
rect 1074 923 1077 936
rect 1082 903 1085 926
rect 1066 883 1077 886
rect 1066 763 1069 816
rect 1074 806 1077 883
rect 1074 803 1085 806
rect 1066 733 1077 736
rect 1066 703 1069 726
rect 1082 706 1085 726
rect 1078 703 1085 706
rect 1078 636 1081 703
rect 1058 613 1061 636
rect 1078 633 1085 636
rect 1082 616 1085 633
rect 1090 626 1093 953
rect 1098 933 1101 1033
rect 1114 1006 1117 1026
rect 1114 1003 1125 1006
rect 1106 923 1109 986
rect 1122 973 1125 996
rect 1114 933 1117 946
rect 1130 933 1133 1233
rect 1138 1116 1141 1343
rect 1146 1283 1149 1336
rect 1154 1303 1157 1396
rect 1162 1323 1165 1396
rect 1178 1386 1181 1433
rect 1186 1413 1189 1616
rect 1198 1566 1201 1623
rect 1194 1563 1201 1566
rect 1174 1383 1181 1386
rect 1174 1326 1177 1383
rect 1186 1363 1189 1406
rect 1194 1403 1197 1563
rect 1210 1546 1213 1893
rect 1218 1813 1221 1826
rect 1218 1733 1221 1806
rect 1234 1803 1237 1966
rect 1242 1856 1245 1936
rect 1250 1923 1253 1946
rect 1258 1933 1261 2076
rect 1242 1853 1261 1856
rect 1258 1813 1261 1853
rect 1226 1706 1229 1726
rect 1222 1703 1229 1706
rect 1222 1636 1225 1703
rect 1222 1633 1229 1636
rect 1218 1603 1221 1616
rect 1202 1543 1213 1546
rect 1186 1333 1189 1346
rect 1170 1323 1177 1326
rect 1146 1213 1149 1226
rect 1146 1133 1149 1156
rect 1138 1113 1145 1116
rect 1142 1036 1145 1113
rect 1138 1033 1145 1036
rect 1138 926 1141 1033
rect 1098 896 1101 916
rect 1122 903 1125 926
rect 1130 923 1141 926
rect 1098 893 1105 896
rect 1102 836 1105 893
rect 1102 833 1109 836
rect 1098 723 1101 826
rect 1106 766 1109 833
rect 1114 803 1117 886
rect 1122 793 1125 846
rect 1130 803 1133 923
rect 1138 813 1141 856
rect 1106 763 1141 766
rect 1106 636 1109 656
rect 1114 643 1117 756
rect 1138 696 1141 763
rect 1130 693 1141 696
rect 1106 633 1117 636
rect 1090 623 1109 626
rect 1074 613 1085 616
rect 1058 533 1061 556
rect 1066 536 1069 606
rect 1082 583 1085 606
rect 1090 603 1093 616
rect 1066 533 1077 536
rect 1042 366 1045 386
rect 1058 383 1061 416
rect 1074 366 1077 533
rect 1082 526 1085 576
rect 1090 533 1093 596
rect 1082 523 1093 526
rect 1042 363 1053 366
rect 1026 323 1029 346
rect 1050 306 1053 363
rect 1042 303 1053 306
rect 1066 363 1077 366
rect 1066 306 1069 363
rect 1066 303 1077 306
rect 1042 283 1045 303
rect 1026 203 1029 216
rect 1074 213 1077 303
rect 1082 213 1085 496
rect 1090 413 1093 523
rect 1098 506 1101 606
rect 1106 573 1109 623
rect 1106 533 1109 556
rect 1114 546 1117 633
rect 1130 613 1133 693
rect 1114 543 1125 546
rect 1114 523 1117 536
rect 1122 516 1125 543
rect 1130 533 1133 576
rect 1138 533 1141 606
rect 1122 513 1133 516
rect 1098 503 1109 506
rect 1106 406 1109 503
rect 1098 403 1109 406
rect 1122 403 1125 506
rect 1130 423 1133 513
rect 1138 413 1141 526
rect 1098 323 1101 403
rect 1146 376 1149 1016
rect 1154 953 1157 1266
rect 1170 1246 1173 1323
rect 1178 1303 1181 1316
rect 1186 1263 1189 1326
rect 1170 1243 1177 1246
rect 1162 1203 1165 1236
rect 1162 1183 1165 1196
rect 1174 1186 1177 1243
rect 1194 1206 1197 1396
rect 1190 1203 1197 1206
rect 1174 1183 1181 1186
rect 1162 1123 1165 1146
rect 1170 1103 1173 1146
rect 1178 1133 1181 1183
rect 1190 1146 1193 1203
rect 1186 1143 1193 1146
rect 1186 1126 1189 1143
rect 1202 1126 1205 1543
rect 1210 1523 1213 1536
rect 1218 1533 1221 1556
rect 1226 1526 1229 1633
rect 1234 1603 1237 1796
rect 1242 1703 1245 1736
rect 1250 1723 1253 1756
rect 1258 1706 1261 1796
rect 1254 1703 1261 1706
rect 1242 1603 1245 1636
rect 1254 1616 1257 1703
rect 1254 1613 1261 1616
rect 1258 1593 1261 1613
rect 1234 1533 1245 1536
rect 1218 1513 1221 1526
rect 1226 1523 1233 1526
rect 1210 1303 1213 1476
rect 1218 1393 1221 1496
rect 1230 1476 1233 1523
rect 1230 1473 1237 1476
rect 1242 1473 1245 1516
rect 1234 1456 1237 1473
rect 1234 1453 1241 1456
rect 1218 1323 1221 1346
rect 1218 1266 1221 1316
rect 1178 1123 1189 1126
rect 1194 1123 1205 1126
rect 1210 1263 1221 1266
rect 1178 1096 1181 1123
rect 1170 1093 1181 1096
rect 1162 946 1165 1016
rect 1170 1003 1173 1093
rect 1194 1076 1197 1123
rect 1210 1116 1213 1263
rect 1218 1213 1221 1256
rect 1218 1153 1221 1196
rect 1226 1136 1229 1446
rect 1238 1356 1241 1453
rect 1250 1413 1253 1446
rect 1258 1413 1261 1516
rect 1250 1393 1253 1406
rect 1234 1353 1241 1356
rect 1234 1333 1237 1353
rect 1266 1346 1269 2083
rect 1274 1933 1277 2006
rect 1274 1823 1277 1926
rect 1282 1923 1285 2076
rect 1290 2013 1293 2056
rect 1290 1956 1293 2006
rect 1306 1966 1309 2106
rect 1314 2053 1317 2266
rect 1326 2206 1329 2283
rect 1338 2276 1341 2286
rect 1346 2283 1365 2286
rect 1338 2273 1357 2276
rect 1326 2203 1333 2206
rect 1322 2073 1325 2186
rect 1330 2006 1333 2203
rect 1338 2183 1341 2266
rect 1346 2103 1349 2226
rect 1338 2013 1341 2026
rect 1330 2003 1341 2006
rect 1346 2003 1349 2076
rect 1354 2063 1357 2273
rect 1362 2223 1365 2283
rect 1370 2256 1373 2293
rect 1386 2283 1389 2336
rect 1394 2263 1397 2416
rect 1402 2413 1405 2463
rect 1410 2453 1413 2516
rect 1418 2486 1421 2806
rect 1426 2803 1429 2833
rect 1434 2803 1437 2816
rect 1426 2633 1429 2796
rect 1442 2783 1445 2826
rect 1450 2763 1453 2816
rect 1458 2813 1461 2936
rect 1466 2923 1469 2976
rect 1474 2906 1477 3046
rect 1470 2903 1477 2906
rect 1470 2816 1473 2903
rect 1466 2813 1473 2816
rect 1466 2783 1469 2813
rect 1482 2806 1485 3076
rect 1490 3013 1493 3256
rect 1498 3223 1501 3333
rect 1506 3326 1509 3356
rect 1506 3323 1525 3326
rect 1498 2996 1501 3206
rect 1490 2993 1501 2996
rect 1506 2976 1509 3316
rect 1522 3276 1525 3323
rect 1530 3313 1533 3526
rect 1538 3463 1541 3526
rect 1538 3413 1541 3426
rect 1538 3336 1541 3406
rect 1546 3346 1549 3626
rect 1554 3613 1557 3626
rect 1554 3533 1557 3556
rect 1562 3546 1565 3636
rect 1570 3553 1573 3643
rect 1562 3543 1573 3546
rect 1554 3403 1557 3526
rect 1562 3413 1565 3446
rect 1546 3343 1557 3346
rect 1538 3333 1549 3336
rect 1538 3313 1541 3326
rect 1530 3283 1533 3306
rect 1522 3273 1533 3276
rect 1514 3226 1517 3246
rect 1530 3226 1533 3273
rect 1538 3233 1541 3306
rect 1514 3223 1525 3226
rect 1530 3223 1541 3226
rect 1514 3183 1517 3223
rect 1530 3203 1533 3216
rect 1514 3113 1517 3126
rect 1530 3116 1533 3166
rect 1538 3126 1541 3223
rect 1546 3136 1549 3333
rect 1554 3253 1557 3343
rect 1562 3313 1565 3406
rect 1570 3353 1573 3543
rect 1578 3523 1581 3706
rect 1586 3623 1589 3666
rect 1602 3653 1605 3733
rect 1610 3723 1613 3746
rect 1650 3736 1653 3876
rect 1658 3773 1661 3846
rect 1594 3546 1597 3626
rect 1602 3583 1605 3636
rect 1610 3623 1613 3676
rect 1594 3543 1605 3546
rect 1586 3483 1589 3516
rect 1578 3413 1581 3466
rect 1586 3413 1589 3426
rect 1578 3373 1581 3406
rect 1594 3396 1597 3536
rect 1602 3496 1605 3543
rect 1610 3523 1613 3566
rect 1618 3516 1621 3646
rect 1626 3623 1629 3736
rect 1634 3733 1653 3736
rect 1634 3633 1637 3733
rect 1642 3723 1661 3726
rect 1642 3616 1645 3723
rect 1626 3603 1629 3616
rect 1634 3613 1645 3616
rect 1650 3613 1653 3716
rect 1658 3713 1661 3723
rect 1658 3663 1661 3706
rect 1626 3523 1629 3596
rect 1634 3583 1637 3613
rect 1658 3606 1661 3636
rect 1642 3573 1645 3606
rect 1650 3603 1661 3606
rect 1634 3516 1637 3536
rect 1642 3523 1645 3536
rect 1618 3513 1637 3516
rect 1602 3493 1613 3496
rect 1610 3436 1613 3493
rect 1634 3483 1637 3513
rect 1650 3503 1653 3603
rect 1586 3393 1597 3396
rect 1602 3433 1613 3436
rect 1570 3333 1573 3346
rect 1562 3213 1565 3226
rect 1546 3133 1557 3136
rect 1538 3123 1549 3126
rect 1530 3113 1549 3116
rect 1514 3013 1517 3076
rect 1530 3003 1533 3106
rect 1538 3013 1541 3026
rect 1546 3013 1549 3113
rect 1562 3103 1565 3176
rect 1570 3083 1573 3326
rect 1578 3203 1581 3286
rect 1586 3143 1589 3393
rect 1594 3303 1597 3386
rect 1594 3225 1597 3266
rect 1602 3236 1605 3433
rect 1610 3403 1613 3416
rect 1610 3276 1613 3376
rect 1626 3373 1629 3416
rect 1642 3413 1645 3446
rect 1634 3336 1637 3406
rect 1650 3396 1653 3426
rect 1658 3403 1661 3586
rect 1666 3463 1669 3816
rect 1674 3803 1677 3886
rect 1682 3766 1685 3856
rect 1690 3823 1693 3933
rect 1698 3913 1701 3936
rect 1714 3923 1717 3936
rect 1722 3933 1725 3943
rect 1690 3813 1701 3816
rect 1690 3803 1693 3813
rect 1698 3793 1701 3806
rect 1682 3763 1693 3766
rect 1682 3713 1685 3756
rect 1690 3733 1693 3763
rect 1698 3723 1701 3786
rect 1706 3753 1709 3856
rect 1714 3833 1717 3906
rect 1714 3736 1717 3826
rect 1722 3783 1725 3816
rect 1730 3796 1733 4013
rect 1738 3983 1741 4006
rect 1754 3993 1757 4006
rect 1770 4003 1773 4143
rect 1778 4073 1781 4213
rect 1786 4153 1789 4206
rect 1794 4136 1797 4266
rect 1850 4263 1853 4340
rect 1802 4166 1805 4246
rect 1818 4223 1829 4226
rect 1850 4223 1853 4236
rect 1810 4213 1821 4216
rect 1826 4213 1829 4223
rect 1810 4193 1813 4213
rect 1818 4186 1821 4206
rect 1810 4183 1821 4186
rect 1826 4183 1829 4206
rect 1834 4203 1853 4206
rect 1802 4163 1813 4166
rect 1810 4146 1813 4163
rect 1810 4143 1817 4146
rect 1786 4133 1797 4136
rect 1778 3996 1781 4026
rect 1770 3993 1781 3996
rect 1786 3993 1789 4133
rect 1738 3926 1741 3936
rect 1746 3933 1757 3936
rect 1738 3923 1749 3926
rect 1754 3826 1757 3933
rect 1762 3913 1765 3976
rect 1770 3843 1773 3993
rect 1738 3813 1741 3826
rect 1754 3823 1765 3826
rect 1746 3803 1749 3816
rect 1730 3793 1741 3796
rect 1706 3733 1717 3736
rect 1674 3703 1701 3706
rect 1674 3623 1677 3666
rect 1682 3573 1685 3626
rect 1690 3613 1693 3636
rect 1698 3613 1701 3703
rect 1706 3616 1709 3733
rect 1714 3663 1717 3726
rect 1722 3713 1725 3736
rect 1730 3676 1733 3776
rect 1754 3756 1757 3816
rect 1746 3753 1757 3756
rect 1722 3673 1733 3676
rect 1714 3623 1717 3646
rect 1722 3623 1725 3673
rect 1738 3643 1741 3736
rect 1746 3723 1749 3753
rect 1754 3723 1757 3736
rect 1730 3623 1733 3636
rect 1706 3613 1717 3616
rect 1714 3583 1717 3613
rect 1738 3596 1741 3616
rect 1722 3593 1741 3596
rect 1722 3576 1725 3593
rect 1706 3573 1725 3576
rect 1674 3466 1677 3526
rect 1682 3486 1685 3536
rect 1690 3493 1693 3566
rect 1706 3526 1709 3573
rect 1698 3523 1709 3526
rect 1698 3513 1701 3523
rect 1714 3516 1717 3526
rect 1706 3513 1717 3516
rect 1730 3513 1733 3586
rect 1746 3556 1749 3636
rect 1754 3623 1757 3636
rect 1762 3576 1765 3823
rect 1770 3783 1773 3836
rect 1778 3753 1781 3986
rect 1786 3903 1789 3966
rect 1794 3933 1797 4126
rect 1814 4086 1817 4143
rect 1834 4133 1837 4203
rect 1858 4193 1861 4286
rect 1938 4283 1941 4340
rect 1946 4337 1981 4340
rect 1866 4183 1869 4206
rect 1874 4173 1877 4216
rect 1882 4166 1885 4206
rect 1890 4196 1893 4216
rect 1906 4213 1909 4276
rect 1922 4213 1925 4276
rect 1938 4223 1941 4266
rect 1930 4213 1941 4216
rect 1930 4206 1933 4213
rect 1914 4203 1933 4206
rect 1938 4196 1941 4206
rect 1890 4193 1941 4196
rect 1882 4163 1893 4166
rect 1826 4113 1829 4126
rect 1842 4123 1845 4136
rect 1866 4133 1869 4146
rect 1898 4143 1901 4186
rect 1882 4133 1893 4136
rect 1906 4133 1909 4146
rect 1858 4093 1861 4126
rect 1866 4113 1869 4126
rect 1914 4123 1917 4176
rect 1930 4133 1933 4156
rect 1946 4143 1949 4337
rect 1994 4316 1997 4340
rect 2010 4326 2013 4340
rect 2058 4337 2085 4340
rect 2098 4337 2117 4340
rect 2010 4323 2021 4326
rect 1970 4313 2005 4316
rect 1810 4083 1817 4086
rect 1802 3826 1805 4016
rect 1810 4003 1813 4083
rect 1850 4026 1853 4046
rect 1850 4023 1861 4026
rect 1826 4003 1829 4016
rect 1810 3926 1813 3936
rect 1818 3933 1821 3966
rect 1810 3923 1821 3926
rect 1826 3916 1829 3956
rect 1842 3933 1845 3996
rect 1858 3956 1861 4023
rect 1850 3953 1861 3956
rect 1818 3913 1829 3916
rect 1834 3916 1837 3926
rect 1834 3913 1845 3916
rect 1786 3823 1805 3826
rect 1786 3803 1789 3823
rect 1794 3783 1797 3816
rect 1810 3773 1813 3836
rect 1818 3803 1821 3913
rect 1826 3813 1829 3866
rect 1834 3803 1837 3913
rect 1850 3896 1853 3953
rect 1858 3923 1861 3936
rect 1874 3933 1877 4016
rect 1890 4003 1893 4116
rect 1954 4086 1957 4286
rect 1962 4173 1965 4216
rect 1970 4193 1973 4313
rect 1986 4173 1989 4246
rect 1962 4126 1965 4146
rect 1994 4133 1997 4216
rect 1962 4123 1969 4126
rect 1938 4083 1957 4086
rect 1906 3963 1909 4016
rect 1890 3933 1893 3956
rect 1866 3906 1869 3926
rect 1882 3913 1885 3926
rect 1898 3906 1901 3936
rect 1906 3923 1909 3956
rect 1914 3953 1917 4016
rect 1938 4003 1941 4083
rect 1966 4066 1969 4123
rect 1962 4063 1969 4066
rect 1962 4046 1965 4063
rect 1954 4043 1965 4046
rect 1922 3946 1925 3996
rect 1914 3943 1925 3946
rect 1914 3916 1917 3943
rect 1930 3936 1933 3956
rect 1922 3933 1933 3936
rect 1938 3933 1941 3986
rect 1922 3923 1925 3933
rect 1930 3923 1941 3926
rect 1914 3913 1929 3916
rect 1866 3903 1901 3906
rect 1906 3903 1917 3906
rect 1850 3893 1869 3896
rect 1842 3813 1845 3846
rect 1858 3813 1861 3836
rect 1834 3786 1837 3796
rect 1858 3786 1861 3806
rect 1834 3783 1861 3786
rect 1786 3736 1789 3746
rect 1770 3733 1789 3736
rect 1770 3603 1773 3726
rect 1786 3713 1789 3726
rect 1778 3593 1781 3676
rect 1794 3646 1797 3736
rect 1802 3693 1805 3726
rect 1810 3723 1813 3736
rect 1818 3683 1821 3736
rect 1826 3723 1829 3776
rect 1834 3713 1837 3736
rect 1790 3643 1797 3646
rect 1762 3573 1773 3576
rect 1738 3553 1749 3556
rect 1698 3486 1701 3506
rect 1706 3493 1717 3496
rect 1682 3483 1701 3486
rect 1674 3463 1681 3466
rect 1666 3423 1669 3436
rect 1618 3333 1637 3336
rect 1642 3393 1653 3396
rect 1618 3323 1621 3333
rect 1626 3323 1637 3326
rect 1618 3283 1621 3316
rect 1626 3293 1629 3323
rect 1634 3276 1637 3316
rect 1642 3303 1645 3393
rect 1666 3383 1669 3416
rect 1678 3366 1681 3463
rect 1690 3413 1693 3426
rect 1706 3406 1709 3426
rect 1702 3403 1709 3406
rect 1690 3373 1693 3396
rect 1650 3313 1653 3356
rect 1658 3293 1661 3316
rect 1666 3313 1669 3366
rect 1674 3363 1681 3366
rect 1610 3273 1629 3276
rect 1634 3273 1653 3276
rect 1602 3233 1621 3236
rect 1594 3222 1605 3225
rect 1610 3183 1613 3206
rect 1618 3176 1621 3233
rect 1626 3213 1629 3273
rect 1634 3213 1637 3266
rect 1642 3206 1645 3226
rect 1650 3223 1653 3273
rect 1658 3213 1661 3256
rect 1578 3113 1581 3136
rect 1602 3133 1605 3176
rect 1610 3173 1621 3176
rect 1634 3203 1645 3206
rect 1610 3133 1613 3173
rect 1634 3163 1637 3203
rect 1642 3173 1661 3176
rect 1666 3173 1669 3306
rect 1586 3116 1589 3126
rect 1586 3113 1597 3116
rect 1602 3103 1605 3126
rect 1626 3093 1629 3136
rect 1634 3113 1637 3156
rect 1642 3133 1645 3173
rect 1658 3166 1661 3173
rect 1674 3166 1677 3363
rect 1682 3306 1685 3346
rect 1690 3313 1693 3356
rect 1702 3336 1705 3403
rect 1702 3333 1709 3336
rect 1714 3333 1717 3493
rect 1698 3306 1701 3316
rect 1682 3303 1701 3306
rect 1682 3293 1693 3296
rect 1682 3233 1685 3256
rect 1690 3226 1693 3293
rect 1698 3233 1701 3296
rect 1706 3263 1709 3333
rect 1650 3123 1653 3166
rect 1658 3163 1677 3166
rect 1682 3153 1685 3226
rect 1690 3223 1701 3226
rect 1698 3213 1701 3223
rect 1706 3206 1709 3246
rect 1690 3203 1709 3206
rect 1554 3003 1557 3046
rect 1578 3013 1581 3046
rect 1586 3023 1589 3056
rect 1522 2993 1533 2996
rect 1490 2973 1509 2976
rect 1490 2923 1493 2973
rect 1498 2883 1501 2936
rect 1490 2813 1493 2866
rect 1474 2776 1477 2806
rect 1482 2803 1493 2806
rect 1498 2803 1501 2876
rect 1458 2773 1477 2776
rect 1442 2686 1445 2736
rect 1434 2683 1445 2686
rect 1426 2496 1429 2606
rect 1434 2546 1437 2683
rect 1442 2603 1445 2636
rect 1442 2556 1445 2596
rect 1450 2563 1453 2756
rect 1442 2553 1453 2556
rect 1434 2543 1445 2546
rect 1434 2503 1437 2526
rect 1426 2493 1437 2496
rect 1418 2483 1429 2486
rect 1402 2353 1405 2406
rect 1410 2376 1413 2446
rect 1418 2383 1421 2436
rect 1426 2413 1429 2483
rect 1434 2406 1437 2493
rect 1426 2403 1437 2406
rect 1410 2373 1421 2376
rect 1402 2316 1405 2346
rect 1410 2343 1413 2366
rect 1418 2343 1421 2373
rect 1426 2336 1429 2403
rect 1442 2396 1445 2543
rect 1450 2533 1453 2553
rect 1458 2516 1461 2773
rect 1466 2733 1469 2766
rect 1490 2756 1493 2796
rect 1506 2766 1509 2926
rect 1514 2913 1517 2936
rect 1522 2886 1525 2926
rect 1514 2883 1525 2886
rect 1514 2793 1517 2883
rect 1546 2876 1549 2936
rect 1570 2933 1573 3006
rect 1594 2996 1597 3016
rect 1586 2993 1597 2996
rect 1602 2993 1605 3036
rect 1522 2873 1549 2876
rect 1474 2753 1493 2756
rect 1498 2763 1509 2766
rect 1466 2683 1469 2726
rect 1466 2553 1469 2656
rect 1474 2593 1477 2753
rect 1498 2746 1501 2763
rect 1514 2756 1517 2786
rect 1506 2753 1517 2756
rect 1498 2743 1509 2746
rect 1482 2703 1485 2736
rect 1498 2723 1501 2734
rect 1490 2613 1493 2696
rect 1482 2576 1485 2606
rect 1498 2603 1501 2686
rect 1506 2596 1509 2743
rect 1514 2603 1517 2706
rect 1474 2573 1485 2576
rect 1474 2533 1477 2573
rect 1482 2523 1485 2566
rect 1490 2543 1493 2596
rect 1498 2593 1509 2596
rect 1450 2473 1453 2516
rect 1458 2513 1465 2516
rect 1462 2446 1465 2513
rect 1490 2503 1493 2516
rect 1498 2496 1501 2593
rect 1482 2493 1501 2496
rect 1458 2443 1465 2446
rect 1450 2403 1453 2436
rect 1418 2333 1429 2336
rect 1434 2393 1445 2396
rect 1402 2313 1413 2316
rect 1402 2266 1405 2306
rect 1410 2303 1413 2313
rect 1418 2306 1421 2333
rect 1426 2313 1429 2326
rect 1418 2303 1429 2306
rect 1402 2263 1413 2266
rect 1370 2253 1397 2256
rect 1362 2196 1365 2216
rect 1362 2193 1373 2196
rect 1362 2056 1365 2186
rect 1370 2126 1373 2193
rect 1378 2186 1381 2206
rect 1386 2203 1389 2246
rect 1394 2193 1397 2253
rect 1402 2226 1405 2263
rect 1418 2233 1421 2286
rect 1402 2223 1413 2226
rect 1402 2186 1405 2223
rect 1418 2216 1421 2226
rect 1378 2183 1405 2186
rect 1410 2213 1421 2216
rect 1410 2143 1413 2213
rect 1370 2123 1381 2126
rect 1370 2073 1373 2123
rect 1378 2096 1381 2106
rect 1394 2103 1397 2136
rect 1378 2093 1393 2096
rect 1354 2053 1365 2056
rect 1314 1973 1325 1976
rect 1298 1963 1309 1966
rect 1314 1956 1317 1966
rect 1290 1953 1301 1956
rect 1290 1856 1293 1946
rect 1282 1853 1293 1856
rect 1282 1776 1285 1853
rect 1282 1773 1293 1776
rect 1274 1613 1277 1736
rect 1282 1713 1285 1726
rect 1282 1656 1285 1696
rect 1290 1666 1293 1773
rect 1298 1693 1301 1953
rect 1306 1953 1317 1956
rect 1306 1933 1309 1953
rect 1322 1946 1325 1973
rect 1314 1943 1325 1946
rect 1306 1676 1309 1926
rect 1314 1823 1317 1943
rect 1314 1803 1317 1816
rect 1322 1793 1325 1936
rect 1330 1923 1333 1996
rect 1338 1936 1341 2003
rect 1346 1943 1349 1956
rect 1338 1933 1349 1936
rect 1354 1933 1357 2053
rect 1378 2023 1381 2056
rect 1390 2036 1393 2093
rect 1390 2033 1397 2036
rect 1386 1973 1389 2016
rect 1394 1966 1397 2033
rect 1362 1963 1397 1966
rect 1338 1843 1341 1926
rect 1346 1836 1349 1933
rect 1362 1926 1365 1963
rect 1330 1833 1349 1836
rect 1354 1923 1365 1926
rect 1314 1783 1325 1786
rect 1314 1703 1317 1783
rect 1330 1776 1333 1833
rect 1338 1803 1341 1826
rect 1346 1796 1349 1826
rect 1354 1813 1357 1923
rect 1362 1906 1365 1916
rect 1362 1903 1369 1906
rect 1366 1836 1369 1903
rect 1366 1833 1373 1836
rect 1370 1813 1373 1833
rect 1362 1803 1373 1806
rect 1322 1773 1333 1776
rect 1306 1673 1317 1676
rect 1290 1663 1309 1666
rect 1282 1653 1301 1656
rect 1282 1633 1293 1636
rect 1282 1526 1285 1633
rect 1274 1523 1285 1526
rect 1290 1506 1293 1536
rect 1298 1523 1301 1653
rect 1290 1503 1297 1506
rect 1282 1456 1285 1496
rect 1274 1453 1285 1456
rect 1274 1423 1277 1453
rect 1282 1403 1285 1446
rect 1294 1436 1297 1503
rect 1290 1433 1297 1436
rect 1290 1413 1293 1433
rect 1306 1413 1309 1663
rect 1314 1603 1317 1673
rect 1314 1513 1317 1596
rect 1322 1563 1325 1773
rect 1330 1613 1333 1696
rect 1338 1676 1341 1796
rect 1346 1793 1365 1796
rect 1338 1673 1349 1676
rect 1322 1523 1325 1536
rect 1330 1496 1333 1606
rect 1338 1563 1341 1606
rect 1322 1493 1333 1496
rect 1322 1436 1325 1493
rect 1322 1433 1333 1436
rect 1330 1413 1333 1433
rect 1290 1403 1325 1406
rect 1250 1343 1269 1346
rect 1234 1213 1237 1306
rect 1242 1143 1245 1336
rect 1250 1253 1253 1343
rect 1250 1173 1253 1216
rect 1258 1203 1261 1336
rect 1266 1186 1269 1326
rect 1274 1276 1277 1326
rect 1282 1323 1285 1396
rect 1290 1386 1293 1403
rect 1290 1383 1297 1386
rect 1294 1316 1297 1383
rect 1290 1313 1297 1316
rect 1290 1293 1293 1313
rect 1298 1293 1309 1296
rect 1274 1273 1289 1276
rect 1262 1183 1269 1186
rect 1218 1133 1229 1136
rect 1178 1073 1197 1076
rect 1202 1113 1213 1116
rect 1218 1123 1237 1126
rect 1154 943 1165 946
rect 1154 913 1157 943
rect 1170 923 1173 976
rect 1178 943 1181 1073
rect 1202 1053 1205 1113
rect 1194 983 1197 1016
rect 1162 903 1165 916
rect 1170 913 1189 916
rect 1170 903 1173 913
rect 1178 836 1181 906
rect 1194 863 1197 926
rect 1202 856 1205 966
rect 1210 916 1213 1106
rect 1218 1076 1221 1123
rect 1226 1096 1229 1116
rect 1234 1113 1253 1116
rect 1234 1103 1237 1113
rect 1242 1103 1253 1106
rect 1262 1096 1265 1183
rect 1226 1093 1265 1096
rect 1274 1086 1277 1226
rect 1286 1206 1289 1273
rect 1306 1266 1309 1293
rect 1314 1276 1317 1346
rect 1314 1273 1333 1276
rect 1306 1263 1325 1266
rect 1298 1213 1301 1226
rect 1286 1203 1293 1206
rect 1306 1203 1309 1263
rect 1282 1153 1285 1186
rect 1258 1083 1277 1086
rect 1218 1073 1237 1076
rect 1218 933 1221 1006
rect 1226 933 1229 1066
rect 1234 1013 1237 1073
rect 1234 923 1237 976
rect 1242 933 1245 1006
rect 1250 973 1253 1026
rect 1210 913 1217 916
rect 1162 833 1181 836
rect 1186 853 1205 856
rect 1154 773 1157 816
rect 1154 723 1157 746
rect 1162 706 1165 833
rect 1170 783 1173 806
rect 1158 703 1165 706
rect 1158 626 1161 703
rect 1178 686 1181 776
rect 1170 683 1181 686
rect 1158 623 1165 626
rect 1162 603 1165 623
rect 1170 613 1173 683
rect 1186 626 1189 853
rect 1214 836 1217 913
rect 1210 833 1217 836
rect 1210 786 1213 833
rect 1218 803 1221 816
rect 1194 703 1197 776
rect 1202 733 1205 786
rect 1210 783 1217 786
rect 1214 726 1217 783
rect 1210 723 1217 726
rect 1186 623 1205 626
rect 1154 553 1157 596
rect 1106 373 1149 376
rect 1106 286 1109 373
rect 1154 366 1157 546
rect 1162 503 1165 596
rect 1178 593 1189 596
rect 1194 593 1197 616
rect 1178 533 1181 593
rect 1194 533 1197 576
rect 1202 546 1205 623
rect 1210 603 1213 723
rect 1202 543 1213 546
rect 1170 523 1181 526
rect 1186 523 1197 526
rect 1170 413 1173 436
rect 1162 383 1165 406
rect 1178 403 1181 523
rect 1194 476 1197 496
rect 1190 473 1197 476
rect 1190 386 1193 473
rect 1202 413 1205 536
rect 1210 493 1213 543
rect 1210 453 1213 486
rect 1190 383 1197 386
rect 1210 383 1213 406
rect 1122 363 1157 366
rect 1122 323 1125 363
rect 1130 333 1133 346
rect 1154 333 1157 356
rect 1194 333 1197 383
rect 1098 283 1109 286
rect 1098 196 1101 283
rect 1138 266 1141 326
rect 1122 263 1181 266
rect 1122 213 1125 263
rect 1106 203 1117 206
rect 1130 203 1133 226
rect 1138 213 1141 236
rect 1178 213 1181 263
rect 1138 196 1141 206
rect 1098 193 1141 196
rect 1034 123 1037 136
rect 1082 123 1085 166
rect 1170 163 1173 206
rect 1186 166 1189 306
rect 1178 163 1189 166
rect 1178 156 1181 163
rect 1162 153 1181 156
rect 1162 123 1165 153
rect 1178 133 1181 146
rect 1194 143 1197 216
rect 1218 213 1221 586
rect 1226 376 1229 866
rect 1234 753 1237 916
rect 1250 883 1253 926
rect 1258 903 1261 1083
rect 1290 1056 1293 1203
rect 1282 1053 1293 1056
rect 1266 966 1269 1026
rect 1282 1023 1285 1053
rect 1282 976 1285 1006
rect 1306 976 1309 1086
rect 1282 973 1309 976
rect 1266 963 1285 966
rect 1290 963 1293 973
rect 1266 896 1269 936
rect 1282 913 1285 963
rect 1314 956 1317 1256
rect 1322 1223 1325 1263
rect 1322 1173 1325 1206
rect 1310 953 1317 956
rect 1266 893 1273 896
rect 1242 703 1245 736
rect 1234 453 1237 636
rect 1242 613 1245 626
rect 1250 613 1253 756
rect 1258 706 1261 866
rect 1270 836 1273 893
rect 1310 876 1313 953
rect 1310 873 1317 876
rect 1314 856 1317 873
rect 1322 863 1325 1156
rect 1330 1083 1333 1273
rect 1338 1213 1341 1556
rect 1346 1516 1349 1673
rect 1346 1513 1353 1516
rect 1350 1446 1353 1513
rect 1346 1443 1353 1446
rect 1346 1423 1349 1443
rect 1346 1313 1349 1326
rect 1354 1323 1357 1406
rect 1346 1163 1349 1296
rect 1362 1276 1365 1793
rect 1370 1723 1373 1803
rect 1378 1793 1381 1936
rect 1402 1836 1405 2136
rect 1410 1916 1413 2066
rect 1418 2033 1421 2206
rect 1418 2003 1421 2026
rect 1418 1973 1421 1996
rect 1418 1923 1421 1966
rect 1410 1913 1417 1916
rect 1414 1856 1417 1913
rect 1426 1866 1429 2303
rect 1434 2133 1437 2393
rect 1442 2333 1445 2346
rect 1442 2116 1445 2326
rect 1450 2316 1453 2396
rect 1458 2383 1461 2443
rect 1466 2403 1469 2426
rect 1474 2396 1477 2446
rect 1482 2413 1485 2493
rect 1490 2423 1501 2426
rect 1466 2393 1477 2396
rect 1458 2333 1461 2366
rect 1466 2323 1469 2393
rect 1450 2313 1457 2316
rect 1454 2246 1457 2313
rect 1474 2266 1477 2336
rect 1482 2333 1485 2386
rect 1450 2243 1457 2246
rect 1450 2223 1453 2243
rect 1466 2223 1469 2266
rect 1474 2263 1485 2266
rect 1474 2243 1477 2263
rect 1474 2216 1477 2226
rect 1450 2193 1453 2216
rect 1466 2213 1477 2216
rect 1466 2163 1469 2213
rect 1450 2123 1453 2136
rect 1466 2126 1469 2136
rect 1474 2133 1477 2206
rect 1482 2156 1485 2216
rect 1490 2193 1493 2423
rect 1506 2383 1509 2546
rect 1514 2416 1517 2526
rect 1522 2423 1525 2873
rect 1530 2783 1533 2816
rect 1546 2736 1549 2826
rect 1546 2733 1557 2736
rect 1530 2613 1533 2636
rect 1538 2616 1541 2696
rect 1546 2676 1549 2726
rect 1554 2683 1557 2733
rect 1562 2686 1565 2836
rect 1570 2806 1573 2866
rect 1586 2826 1589 2993
rect 1618 2986 1621 3046
rect 1626 3023 1629 3056
rect 1634 3003 1637 3076
rect 1658 3033 1661 3136
rect 1666 3043 1669 3146
rect 1690 3126 1693 3203
rect 1674 3123 1693 3126
rect 1698 3136 1701 3196
rect 1714 3173 1717 3326
rect 1722 3223 1725 3496
rect 1730 3383 1733 3506
rect 1738 3423 1741 3553
rect 1746 3513 1749 3546
rect 1762 3543 1765 3566
rect 1770 3536 1773 3573
rect 1754 3506 1757 3536
rect 1762 3533 1773 3536
rect 1762 3513 1765 3533
rect 1770 3523 1781 3526
rect 1746 3496 1749 3506
rect 1754 3503 1773 3506
rect 1746 3493 1765 3496
rect 1746 3416 1749 3486
rect 1738 3413 1749 3416
rect 1730 3296 1733 3376
rect 1738 3303 1741 3406
rect 1754 3403 1757 3426
rect 1746 3313 1749 3336
rect 1730 3293 1749 3296
rect 1730 3233 1733 3256
rect 1738 3223 1741 3286
rect 1746 3223 1749 3293
rect 1754 3283 1757 3346
rect 1762 3333 1765 3493
rect 1778 3413 1781 3516
rect 1790 3506 1793 3643
rect 1802 3623 1805 3636
rect 1802 3593 1805 3616
rect 1810 3566 1813 3626
rect 1826 3606 1829 3616
rect 1826 3603 1837 3606
rect 1842 3603 1845 3746
rect 1850 3693 1853 3716
rect 1858 3703 1861 3746
rect 1866 3733 1869 3893
rect 1866 3686 1869 3716
rect 1858 3683 1869 3686
rect 1850 3613 1853 3626
rect 1826 3576 1829 3596
rect 1834 3586 1837 3603
rect 1834 3583 1845 3586
rect 1802 3563 1813 3566
rect 1822 3573 1829 3576
rect 1790 3503 1797 3506
rect 1786 3423 1789 3486
rect 1770 3356 1773 3406
rect 1770 3353 1789 3356
rect 1770 3296 1773 3336
rect 1778 3323 1781 3346
rect 1762 3293 1773 3296
rect 1762 3276 1765 3293
rect 1754 3273 1765 3276
rect 1754 3223 1757 3273
rect 1762 3233 1765 3266
rect 1778 3263 1781 3316
rect 1770 3223 1773 3256
rect 1730 3213 1781 3216
rect 1698 3133 1717 3136
rect 1674 3113 1677 3123
rect 1682 3083 1685 3116
rect 1698 3103 1701 3133
rect 1706 3103 1709 3116
rect 1714 3113 1717 3133
rect 1706 3023 1709 3086
rect 1722 3046 1725 3206
rect 1730 3133 1733 3213
rect 1738 3186 1741 3206
rect 1738 3183 1745 3186
rect 1742 3126 1745 3183
rect 1786 3156 1789 3353
rect 1794 3223 1797 3503
rect 1802 3413 1805 3563
rect 1822 3516 1825 3573
rect 1834 3526 1837 3576
rect 1842 3566 1845 3583
rect 1858 3573 1861 3683
rect 1874 3676 1877 3866
rect 1882 3773 1885 3816
rect 1890 3746 1893 3903
rect 1906 3746 1909 3903
rect 1926 3856 1929 3913
rect 1926 3853 1933 3856
rect 1882 3743 1893 3746
rect 1898 3733 1901 3746
rect 1906 3743 1917 3746
rect 1898 3693 1901 3726
rect 1906 3703 1909 3736
rect 1866 3673 1877 3676
rect 1866 3603 1869 3673
rect 1882 3666 1885 3676
rect 1874 3663 1885 3666
rect 1874 3613 1877 3663
rect 1842 3563 1861 3566
rect 1834 3523 1845 3526
rect 1858 3523 1861 3563
rect 1810 3503 1813 3516
rect 1822 3513 1829 3516
rect 1818 3436 1821 3486
rect 1826 3456 1829 3513
rect 1842 3513 1853 3516
rect 1826 3453 1837 3456
rect 1810 3423 1813 3436
rect 1818 3433 1829 3436
rect 1802 3323 1805 3406
rect 1738 3123 1745 3126
rect 1754 3153 1789 3156
rect 1794 3153 1797 3206
rect 1802 3203 1805 3296
rect 1810 3213 1813 3366
rect 1738 3073 1741 3123
rect 1754 3076 1757 3153
rect 1810 3143 1813 3156
rect 1778 3083 1781 3126
rect 1754 3073 1789 3076
rect 1722 3043 1733 3046
rect 1714 3033 1725 3036
rect 1618 2983 1661 2986
rect 1594 2886 1597 2926
rect 1594 2883 1605 2886
rect 1578 2813 1581 2826
rect 1586 2823 1597 2826
rect 1570 2803 1581 2806
rect 1578 2783 1581 2803
rect 1586 2766 1589 2816
rect 1570 2763 1589 2766
rect 1570 2693 1573 2763
rect 1594 2706 1597 2823
rect 1602 2803 1605 2883
rect 1610 2836 1613 2846
rect 1610 2833 1629 2836
rect 1634 2833 1637 2926
rect 1642 2923 1645 2936
rect 1642 2866 1645 2886
rect 1650 2873 1653 2936
rect 1642 2863 1653 2866
rect 1610 2813 1613 2833
rect 1618 2803 1621 2826
rect 1642 2823 1645 2856
rect 1634 2783 1637 2806
rect 1650 2766 1653 2863
rect 1658 2836 1661 2983
rect 1682 2936 1685 3006
rect 1722 2963 1725 3026
rect 1674 2933 1685 2936
rect 1666 2883 1669 2926
rect 1658 2833 1669 2836
rect 1658 2813 1661 2826
rect 1666 2803 1669 2833
rect 1674 2826 1677 2933
rect 1682 2886 1685 2926
rect 1690 2913 1693 2936
rect 1706 2886 1709 2936
rect 1730 2933 1733 3043
rect 1738 2976 1741 3006
rect 1786 3003 1789 3073
rect 1794 3013 1797 3076
rect 1738 2973 1745 2976
rect 1742 2926 1745 2973
rect 1794 2963 1797 2996
rect 1738 2923 1745 2926
rect 1682 2883 1701 2886
rect 1706 2883 1725 2886
rect 1698 2846 1701 2883
rect 1698 2843 1709 2846
rect 1674 2823 1685 2826
rect 1698 2823 1701 2836
rect 1674 2786 1677 2816
rect 1586 2703 1597 2706
rect 1602 2703 1605 2766
rect 1610 2763 1653 2766
rect 1658 2783 1677 2786
rect 1610 2726 1613 2763
rect 1658 2756 1661 2783
rect 1682 2776 1685 2823
rect 1690 2813 1701 2816
rect 1698 2783 1701 2813
rect 1674 2773 1685 2776
rect 1634 2753 1661 2756
rect 1618 2733 1629 2736
rect 1610 2723 1621 2726
rect 1626 2723 1629 2733
rect 1562 2683 1581 2686
rect 1546 2673 1557 2676
rect 1538 2613 1549 2616
rect 1538 2563 1541 2606
rect 1530 2533 1541 2536
rect 1514 2413 1525 2416
rect 1530 2413 1533 2526
rect 1538 2513 1541 2526
rect 1546 2496 1549 2613
rect 1554 2603 1557 2673
rect 1562 2613 1565 2676
rect 1570 2586 1573 2636
rect 1542 2493 1549 2496
rect 1554 2583 1573 2586
rect 1542 2426 1545 2493
rect 1554 2443 1557 2583
rect 1578 2576 1581 2683
rect 1562 2573 1581 2576
rect 1562 2523 1565 2573
rect 1570 2533 1573 2566
rect 1538 2423 1545 2426
rect 1522 2406 1525 2413
rect 1538 2406 1541 2423
rect 1546 2413 1557 2416
rect 1514 2366 1517 2406
rect 1522 2403 1533 2406
rect 1538 2403 1549 2406
rect 1554 2403 1557 2413
rect 1506 2363 1517 2366
rect 1498 2313 1501 2346
rect 1482 2153 1493 2156
rect 1434 2083 1437 2116
rect 1442 2113 1449 2116
rect 1446 2056 1449 2113
rect 1446 2053 1453 2056
rect 1442 2013 1445 2036
rect 1450 2016 1453 2053
rect 1458 2023 1461 2126
rect 1466 2123 1477 2126
rect 1466 2103 1469 2116
rect 1474 2096 1477 2123
rect 1466 2093 1477 2096
rect 1450 2013 1461 2016
rect 1434 1963 1437 2006
rect 1450 2003 1453 2013
rect 1426 1863 1433 1866
rect 1414 1853 1421 1856
rect 1394 1793 1397 1836
rect 1402 1833 1413 1836
rect 1418 1813 1421 1853
rect 1402 1786 1405 1806
rect 1410 1803 1421 1806
rect 1402 1783 1409 1786
rect 1378 1623 1381 1726
rect 1386 1593 1389 1736
rect 1406 1686 1409 1783
rect 1402 1683 1409 1686
rect 1402 1643 1405 1683
rect 1418 1626 1421 1803
rect 1430 1786 1433 1863
rect 1426 1783 1433 1786
rect 1426 1706 1429 1783
rect 1434 1723 1437 1766
rect 1426 1703 1433 1706
rect 1430 1636 1433 1703
rect 1394 1623 1421 1626
rect 1426 1633 1433 1636
rect 1442 1636 1445 1996
rect 1450 1913 1453 1966
rect 1458 1856 1461 2006
rect 1450 1853 1461 1856
rect 1450 1803 1453 1853
rect 1466 1826 1469 2093
rect 1474 2003 1477 2026
rect 1482 1946 1485 2116
rect 1474 1943 1485 1946
rect 1474 1916 1477 1943
rect 1490 1936 1493 2153
rect 1498 1996 1501 2306
rect 1506 2303 1509 2363
rect 1506 2183 1509 2206
rect 1506 2083 1509 2106
rect 1506 2003 1509 2016
rect 1498 1993 1509 1996
rect 1482 1933 1493 1936
rect 1506 1936 1509 1993
rect 1514 1946 1517 2346
rect 1522 2196 1525 2396
rect 1530 2203 1533 2403
rect 1538 2343 1541 2386
rect 1546 2336 1549 2403
rect 1562 2346 1565 2416
rect 1570 2403 1573 2476
rect 1554 2343 1565 2346
rect 1538 2303 1541 2336
rect 1546 2333 1557 2336
rect 1570 2333 1573 2346
rect 1538 2213 1541 2246
rect 1546 2203 1549 2326
rect 1522 2193 1541 2196
rect 1522 2133 1525 2186
rect 1522 2113 1525 2126
rect 1522 2063 1525 2106
rect 1530 2053 1533 2186
rect 1538 2156 1541 2193
rect 1554 2183 1557 2333
rect 1562 2256 1565 2326
rect 1578 2323 1581 2526
rect 1562 2253 1581 2256
rect 1570 2226 1573 2246
rect 1578 2236 1581 2253
rect 1586 2243 1589 2703
rect 1610 2696 1613 2716
rect 1594 2613 1597 2696
rect 1602 2693 1613 2696
rect 1594 2566 1597 2606
rect 1602 2573 1605 2693
rect 1618 2646 1621 2723
rect 1634 2716 1637 2753
rect 1666 2736 1669 2756
rect 1642 2733 1653 2736
rect 1658 2733 1669 2736
rect 1642 2723 1645 2733
rect 1634 2713 1645 2716
rect 1650 2703 1653 2726
rect 1610 2643 1621 2646
rect 1626 2693 1637 2696
rect 1610 2596 1613 2643
rect 1618 2613 1621 2636
rect 1626 2613 1629 2693
rect 1634 2613 1637 2626
rect 1618 2603 1637 2606
rect 1642 2603 1645 2636
rect 1658 2616 1661 2733
rect 1666 2703 1669 2726
rect 1674 2636 1677 2773
rect 1706 2766 1709 2843
rect 1714 2803 1717 2816
rect 1682 2686 1685 2766
rect 1698 2763 1709 2766
rect 1690 2735 1693 2756
rect 1698 2731 1701 2763
rect 1690 2728 1701 2731
rect 1690 2693 1693 2728
rect 1698 2696 1701 2724
rect 1706 2703 1709 2736
rect 1698 2693 1717 2696
rect 1682 2683 1701 2686
rect 1674 2633 1685 2636
rect 1690 2633 1693 2676
rect 1610 2593 1629 2596
rect 1594 2563 1605 2566
rect 1602 2496 1605 2563
rect 1594 2493 1605 2496
rect 1594 2443 1597 2493
rect 1626 2486 1629 2593
rect 1602 2483 1629 2486
rect 1594 2403 1597 2426
rect 1602 2413 1605 2483
rect 1610 2453 1629 2456
rect 1610 2443 1613 2453
rect 1610 2386 1613 2436
rect 1594 2383 1613 2386
rect 1594 2343 1597 2383
rect 1618 2376 1621 2426
rect 1602 2373 1621 2376
rect 1626 2373 1629 2446
rect 1594 2283 1597 2336
rect 1602 2326 1605 2373
rect 1610 2343 1613 2366
rect 1602 2323 1609 2326
rect 1606 2276 1609 2323
rect 1602 2273 1609 2276
rect 1578 2233 1589 2236
rect 1570 2223 1581 2226
rect 1562 2156 1565 2206
rect 1570 2203 1573 2216
rect 1578 2203 1581 2223
rect 1538 2153 1549 2156
rect 1562 2153 1573 2156
rect 1546 2076 1549 2153
rect 1570 2123 1573 2153
rect 1578 2143 1581 2186
rect 1538 2073 1549 2076
rect 1530 2006 1533 2016
rect 1522 2003 1533 2006
rect 1514 1943 1525 1946
rect 1530 1943 1533 2003
rect 1538 1993 1541 2073
rect 1546 2003 1549 2066
rect 1554 2003 1557 2026
rect 1562 1966 1565 2056
rect 1538 1963 1565 1966
rect 1506 1933 1517 1936
rect 1474 1913 1481 1916
rect 1490 1913 1493 1926
rect 1478 1836 1481 1913
rect 1498 1846 1501 1926
rect 1498 1843 1509 1846
rect 1478 1833 1485 1836
rect 1490 1833 1501 1836
rect 1506 1833 1509 1843
rect 1458 1823 1469 1826
rect 1458 1813 1461 1823
rect 1458 1802 1468 1805
rect 1474 1803 1477 1816
rect 1450 1733 1453 1796
rect 1458 1733 1461 1802
rect 1458 1643 1461 1726
rect 1442 1633 1461 1636
rect 1394 1586 1397 1623
rect 1402 1613 1421 1616
rect 1402 1603 1405 1613
rect 1370 1583 1397 1586
rect 1370 1563 1373 1583
rect 1410 1576 1413 1606
rect 1378 1573 1413 1576
rect 1378 1523 1381 1573
rect 1386 1533 1389 1566
rect 1426 1563 1429 1633
rect 1434 1603 1437 1616
rect 1458 1603 1461 1633
rect 1466 1586 1469 1796
rect 1462 1583 1469 1586
rect 1394 1523 1397 1556
rect 1378 1343 1381 1406
rect 1386 1276 1389 1376
rect 1394 1323 1397 1336
rect 1362 1273 1369 1276
rect 1338 1123 1341 1156
rect 1354 1103 1357 1266
rect 1366 1196 1369 1273
rect 1378 1273 1389 1276
rect 1402 1273 1405 1536
rect 1450 1526 1453 1546
rect 1378 1253 1381 1273
rect 1410 1266 1413 1416
rect 1418 1363 1421 1526
rect 1442 1523 1453 1526
rect 1462 1526 1465 1583
rect 1474 1533 1477 1726
rect 1482 1593 1485 1833
rect 1490 1793 1493 1826
rect 1490 1723 1493 1756
rect 1462 1523 1469 1526
rect 1442 1466 1445 1523
rect 1466 1476 1469 1523
rect 1482 1513 1485 1586
rect 1490 1576 1493 1626
rect 1498 1613 1501 1833
rect 1514 1806 1517 1916
rect 1522 1813 1525 1943
rect 1530 1906 1533 1936
rect 1538 1923 1541 1936
rect 1546 1913 1549 1946
rect 1562 1913 1565 1963
rect 1570 1943 1573 2066
rect 1578 1973 1581 2126
rect 1530 1903 1537 1906
rect 1534 1846 1537 1903
rect 1530 1843 1537 1846
rect 1530 1813 1533 1843
rect 1570 1813 1573 1936
rect 1578 1923 1581 1956
rect 1586 1933 1589 2233
rect 1594 2123 1597 2206
rect 1602 2193 1605 2273
rect 1618 2246 1621 2356
rect 1626 2323 1629 2346
rect 1634 2306 1637 2603
rect 1650 2583 1653 2616
rect 1658 2613 1669 2616
rect 1658 2563 1661 2606
rect 1674 2583 1677 2606
rect 1682 2576 1685 2633
rect 1690 2603 1693 2626
rect 1674 2573 1685 2576
rect 1642 2523 1645 2536
rect 1614 2243 1621 2246
rect 1630 2303 1637 2306
rect 1614 2156 1617 2243
rect 1630 2236 1633 2303
rect 1626 2233 1633 2236
rect 1626 2206 1629 2233
rect 1634 2213 1637 2226
rect 1626 2203 1637 2206
rect 1626 2183 1629 2196
rect 1610 2153 1617 2156
rect 1594 2083 1597 2106
rect 1602 2013 1605 2056
rect 1610 2006 1613 2153
rect 1618 2013 1621 2126
rect 1626 2123 1629 2166
rect 1594 1986 1597 2006
rect 1610 2003 1621 2006
rect 1594 1983 1613 1986
rect 1514 1803 1533 1806
rect 1514 1793 1525 1796
rect 1506 1593 1509 1736
rect 1514 1733 1517 1793
rect 1514 1686 1517 1726
rect 1522 1703 1525 1766
rect 1514 1683 1521 1686
rect 1518 1616 1521 1683
rect 1514 1613 1521 1616
rect 1490 1573 1501 1576
rect 1490 1523 1493 1566
rect 1466 1473 1477 1476
rect 1442 1463 1449 1466
rect 1426 1366 1429 1416
rect 1446 1396 1449 1463
rect 1446 1393 1453 1396
rect 1458 1393 1461 1416
rect 1450 1376 1453 1393
rect 1450 1373 1461 1376
rect 1426 1363 1453 1366
rect 1458 1346 1461 1373
rect 1474 1356 1477 1473
rect 1498 1436 1501 1573
rect 1506 1523 1509 1536
rect 1514 1473 1517 1613
rect 1530 1603 1533 1803
rect 1546 1733 1549 1806
rect 1578 1796 1581 1836
rect 1562 1793 1581 1796
rect 1538 1713 1541 1726
rect 1442 1343 1461 1346
rect 1466 1353 1477 1356
rect 1490 1433 1501 1436
rect 1490 1356 1493 1433
rect 1506 1413 1509 1426
rect 1490 1353 1501 1356
rect 1418 1323 1421 1336
rect 1386 1263 1413 1266
rect 1362 1193 1369 1196
rect 1330 963 1333 1016
rect 1346 966 1349 986
rect 1346 963 1353 966
rect 1330 903 1333 926
rect 1350 906 1353 963
rect 1346 903 1353 906
rect 1346 886 1349 903
rect 1338 883 1349 886
rect 1314 853 1325 856
rect 1266 833 1273 836
rect 1266 786 1269 833
rect 1290 803 1293 816
rect 1266 783 1293 786
rect 1266 733 1269 746
rect 1274 723 1277 736
rect 1282 733 1285 756
rect 1290 733 1293 783
rect 1322 753 1325 853
rect 1330 783 1333 816
rect 1258 703 1269 706
rect 1266 626 1269 703
rect 1266 623 1277 626
rect 1242 573 1245 606
rect 1258 593 1261 606
rect 1266 583 1269 616
rect 1242 553 1269 556
rect 1242 523 1245 553
rect 1258 526 1261 536
rect 1250 523 1261 526
rect 1250 456 1253 523
rect 1258 493 1261 516
rect 1266 503 1269 536
rect 1274 496 1277 623
rect 1282 553 1285 666
rect 1290 576 1293 616
rect 1298 593 1301 606
rect 1290 573 1297 576
rect 1306 573 1309 636
rect 1314 613 1317 746
rect 1338 736 1341 883
rect 1362 813 1365 1193
rect 1370 1123 1373 1176
rect 1378 1143 1381 1186
rect 1378 1106 1381 1136
rect 1374 1103 1381 1106
rect 1374 1026 1377 1103
rect 1374 1023 1381 1026
rect 1370 973 1373 1006
rect 1378 953 1381 1023
rect 1370 883 1373 926
rect 1322 703 1325 736
rect 1334 733 1341 736
rect 1354 733 1357 806
rect 1370 773 1373 806
rect 1334 636 1337 733
rect 1346 636 1349 726
rect 1362 723 1365 736
rect 1370 733 1373 746
rect 1378 703 1381 736
rect 1386 706 1389 1263
rect 1426 1256 1429 1336
rect 1402 1253 1429 1256
rect 1394 1183 1397 1216
rect 1402 1173 1405 1253
rect 1434 1246 1437 1286
rect 1426 1243 1437 1246
rect 1394 1023 1397 1146
rect 1402 1126 1405 1166
rect 1410 1136 1413 1216
rect 1426 1213 1429 1243
rect 1418 1153 1421 1206
rect 1434 1183 1437 1206
rect 1410 1133 1421 1136
rect 1402 1123 1413 1126
rect 1418 1116 1421 1133
rect 1410 1113 1421 1116
rect 1442 1116 1445 1343
rect 1450 1263 1453 1326
rect 1450 1203 1453 1236
rect 1458 1133 1461 1256
rect 1442 1113 1453 1116
rect 1394 933 1397 1006
rect 1402 973 1405 1016
rect 1402 913 1405 926
rect 1410 923 1413 1113
rect 1418 1086 1421 1106
rect 1418 1083 1429 1086
rect 1426 1036 1429 1083
rect 1418 1033 1429 1036
rect 1418 1013 1421 1033
rect 1426 966 1429 1006
rect 1418 963 1429 966
rect 1426 903 1429 936
rect 1434 923 1437 1016
rect 1442 973 1445 1006
rect 1442 913 1445 936
rect 1450 896 1453 1113
rect 1458 913 1461 1066
rect 1446 893 1453 896
rect 1394 803 1397 836
rect 1402 823 1437 826
rect 1402 743 1405 823
rect 1410 813 1421 816
rect 1386 703 1393 706
rect 1362 683 1381 686
rect 1362 673 1365 683
rect 1334 633 1341 636
rect 1346 633 1357 636
rect 1322 603 1325 626
rect 1266 493 1277 496
rect 1242 453 1253 456
rect 1242 433 1245 453
rect 1226 373 1233 376
rect 1218 183 1221 206
rect 1230 196 1233 373
rect 1242 363 1245 406
rect 1266 386 1269 493
rect 1262 383 1269 386
rect 1242 323 1245 346
rect 1262 316 1265 383
rect 1274 323 1277 386
rect 1262 313 1269 316
rect 1266 293 1269 313
rect 1250 203 1253 216
rect 1230 193 1237 196
rect 1234 176 1237 193
rect 1234 173 1261 176
rect 1218 123 1221 146
rect 1258 123 1261 173
rect 1282 83 1285 526
rect 1294 496 1297 573
rect 1290 493 1297 496
rect 1306 513 1317 516
rect 1306 493 1309 513
rect 1322 496 1325 536
rect 1314 493 1325 496
rect 1290 473 1293 493
rect 1290 383 1293 416
rect 1290 326 1293 376
rect 1306 373 1309 406
rect 1314 376 1317 493
rect 1330 476 1333 616
rect 1326 473 1333 476
rect 1326 406 1329 473
rect 1326 403 1333 406
rect 1338 403 1341 633
rect 1346 593 1349 626
rect 1354 543 1357 633
rect 1362 613 1373 616
rect 1378 613 1381 676
rect 1390 636 1393 703
rect 1410 686 1413 813
rect 1418 796 1421 806
rect 1426 803 1429 816
rect 1434 803 1437 823
rect 1446 796 1449 893
rect 1418 793 1449 796
rect 1426 733 1429 786
rect 1458 776 1461 906
rect 1466 863 1469 1353
rect 1474 1313 1477 1336
rect 1482 1333 1493 1336
rect 1498 1326 1501 1353
rect 1506 1333 1509 1406
rect 1514 1353 1517 1416
rect 1482 1283 1485 1326
rect 1498 1323 1517 1326
rect 1498 1253 1501 1316
rect 1506 1233 1509 1316
rect 1474 1223 1493 1226
rect 1474 1156 1477 1223
rect 1490 1216 1493 1223
rect 1482 1183 1485 1216
rect 1490 1213 1501 1216
rect 1506 1203 1509 1226
rect 1474 1153 1485 1156
rect 1474 1003 1477 1136
rect 1482 996 1485 1153
rect 1490 1106 1493 1156
rect 1498 1123 1501 1176
rect 1490 1103 1497 1106
rect 1494 1036 1497 1103
rect 1474 993 1485 996
rect 1490 1033 1497 1036
rect 1474 913 1477 993
rect 1490 973 1493 1033
rect 1498 983 1501 1016
rect 1454 773 1461 776
rect 1434 723 1437 736
rect 1442 716 1445 736
rect 1454 726 1457 773
rect 1466 766 1469 816
rect 1474 803 1477 906
rect 1482 813 1485 926
rect 1490 803 1493 956
rect 1498 893 1501 936
rect 1498 813 1501 836
rect 1506 786 1509 1146
rect 1514 933 1517 1323
rect 1522 1133 1525 1596
rect 1530 1533 1533 1566
rect 1546 1523 1549 1626
rect 1554 1613 1557 1726
rect 1530 1493 1533 1516
rect 1538 1413 1541 1426
rect 1530 1363 1533 1406
rect 1546 1403 1549 1416
rect 1554 1396 1557 1536
rect 1562 1506 1565 1793
rect 1578 1743 1581 1756
rect 1570 1703 1573 1736
rect 1586 1723 1589 1826
rect 1570 1603 1573 1616
rect 1578 1603 1581 1666
rect 1594 1663 1597 1976
rect 1610 1973 1613 1983
rect 1610 1846 1613 1946
rect 1618 1923 1621 2003
rect 1610 1843 1621 1846
rect 1602 1703 1605 1726
rect 1610 1723 1613 1836
rect 1618 1753 1621 1843
rect 1586 1613 1589 1656
rect 1618 1613 1621 1656
rect 1626 1596 1629 2116
rect 1634 2063 1637 2203
rect 1642 2156 1645 2456
rect 1650 2413 1653 2526
rect 1666 2486 1669 2536
rect 1658 2483 1669 2486
rect 1658 2386 1661 2483
rect 1666 2403 1669 2416
rect 1674 2396 1677 2573
rect 1682 2523 1685 2566
rect 1690 2503 1693 2536
rect 1698 2506 1701 2683
rect 1714 2623 1717 2693
rect 1722 2656 1725 2883
rect 1738 2876 1741 2923
rect 1738 2873 1745 2876
rect 1730 2803 1733 2866
rect 1742 2826 1745 2873
rect 1742 2823 1749 2826
rect 1738 2763 1741 2816
rect 1746 2766 1749 2823
rect 1754 2803 1757 2926
rect 1762 2813 1765 2846
rect 1770 2803 1773 2836
rect 1778 2766 1781 2896
rect 1746 2763 1757 2766
rect 1746 2723 1749 2756
rect 1754 2706 1757 2763
rect 1770 2763 1781 2766
rect 1770 2753 1773 2763
rect 1750 2703 1757 2706
rect 1722 2653 1741 2656
rect 1738 2626 1741 2653
rect 1750 2646 1753 2703
rect 1750 2643 1757 2646
rect 1738 2623 1749 2626
rect 1714 2563 1717 2606
rect 1738 2576 1741 2616
rect 1746 2583 1749 2623
rect 1722 2573 1741 2576
rect 1706 2523 1709 2546
rect 1722 2533 1725 2573
rect 1730 2513 1733 2526
rect 1698 2503 1709 2506
rect 1746 2503 1749 2526
rect 1682 2403 1685 2476
rect 1706 2446 1709 2503
rect 1698 2443 1709 2446
rect 1674 2393 1685 2396
rect 1658 2383 1677 2386
rect 1650 2313 1653 2376
rect 1666 2333 1669 2366
rect 1658 2226 1661 2326
rect 1674 2323 1677 2383
rect 1682 2306 1685 2393
rect 1690 2313 1693 2416
rect 1674 2303 1685 2306
rect 1674 2246 1677 2303
rect 1690 2263 1693 2306
rect 1674 2243 1685 2246
rect 1658 2223 1677 2226
rect 1650 2203 1653 2216
rect 1658 2166 1661 2206
rect 1666 2183 1669 2216
rect 1658 2163 1669 2166
rect 1642 2153 1653 2156
rect 1650 2063 1653 2153
rect 1666 2143 1669 2163
rect 1674 2123 1677 2223
rect 1682 2076 1685 2243
rect 1690 2203 1693 2226
rect 1698 2176 1701 2443
rect 1706 2303 1709 2386
rect 1722 2356 1725 2406
rect 1746 2403 1749 2476
rect 1714 2353 1725 2356
rect 1722 2333 1725 2346
rect 1714 2226 1717 2326
rect 1730 2323 1733 2356
rect 1746 2336 1749 2376
rect 1738 2333 1749 2336
rect 1722 2236 1725 2316
rect 1738 2306 1741 2333
rect 1730 2303 1741 2306
rect 1730 2283 1733 2303
rect 1746 2296 1749 2326
rect 1738 2293 1749 2296
rect 1722 2233 1733 2236
rect 1714 2223 1725 2226
rect 1690 2173 1701 2176
rect 1690 2163 1693 2173
rect 1706 2166 1709 2206
rect 1714 2203 1717 2216
rect 1698 2163 1709 2166
rect 1698 2156 1701 2163
rect 1690 2153 1701 2156
rect 1690 2123 1693 2153
rect 1658 2073 1685 2076
rect 1634 2033 1645 2036
rect 1634 1933 1637 2033
rect 1658 1986 1661 2073
rect 1658 1983 1669 1986
rect 1634 1916 1637 1926
rect 1642 1923 1645 1936
rect 1650 1933 1653 1946
rect 1634 1913 1653 1916
rect 1634 1843 1637 1856
rect 1634 1793 1637 1816
rect 1642 1813 1645 1886
rect 1650 1853 1653 1913
rect 1658 1883 1661 1966
rect 1666 1943 1669 1983
rect 1674 1936 1677 2066
rect 1698 2026 1701 2146
rect 1698 2023 1709 2026
rect 1698 1973 1701 2016
rect 1706 1953 1709 2023
rect 1714 1946 1717 2166
rect 1722 1966 1725 2223
rect 1730 2213 1733 2233
rect 1730 2183 1733 2206
rect 1730 2123 1733 2166
rect 1738 2156 1741 2293
rect 1746 2193 1749 2286
rect 1746 2163 1749 2186
rect 1738 2153 1749 2156
rect 1738 2073 1741 2086
rect 1738 1976 1741 2066
rect 1730 1973 1741 1976
rect 1746 1973 1749 2153
rect 1722 1963 1749 1966
rect 1670 1933 1677 1936
rect 1670 1856 1673 1933
rect 1666 1853 1673 1856
rect 1650 1803 1653 1846
rect 1666 1836 1669 1853
rect 1658 1833 1669 1836
rect 1618 1593 1629 1596
rect 1578 1533 1581 1566
rect 1562 1503 1581 1506
rect 1546 1393 1557 1396
rect 1530 1273 1533 1356
rect 1546 1326 1549 1393
rect 1538 1323 1549 1326
rect 1554 1323 1557 1336
rect 1538 1306 1541 1323
rect 1538 1303 1549 1306
rect 1530 1223 1533 1266
rect 1546 1236 1549 1303
rect 1538 1233 1549 1236
rect 1538 1213 1541 1233
rect 1562 1216 1565 1346
rect 1570 1323 1573 1416
rect 1578 1323 1581 1503
rect 1602 1416 1605 1526
rect 1618 1486 1621 1593
rect 1634 1566 1637 1736
rect 1642 1723 1645 1756
rect 1658 1733 1661 1833
rect 1682 1826 1685 1946
rect 1698 1943 1717 1946
rect 1666 1823 1685 1826
rect 1650 1636 1653 1656
rect 1642 1603 1645 1636
rect 1650 1633 1661 1636
rect 1650 1613 1653 1633
rect 1666 1626 1669 1823
rect 1690 1816 1693 1936
rect 1674 1793 1677 1816
rect 1682 1813 1693 1816
rect 1682 1763 1685 1813
rect 1658 1623 1669 1626
rect 1674 1623 1677 1706
rect 1682 1663 1685 1726
rect 1690 1716 1693 1806
rect 1698 1733 1701 1943
rect 1706 1896 1709 1916
rect 1714 1906 1717 1936
rect 1722 1923 1725 1946
rect 1730 1913 1733 1936
rect 1738 1923 1741 1956
rect 1746 1923 1749 1963
rect 1754 1943 1757 2643
rect 1762 2543 1765 2706
rect 1786 2636 1789 2926
rect 1794 2893 1797 2926
rect 1794 2843 1797 2866
rect 1778 2633 1789 2636
rect 1778 2576 1781 2633
rect 1794 2616 1797 2836
rect 1770 2573 1781 2576
rect 1790 2613 1797 2616
rect 1762 2503 1765 2536
rect 1770 2523 1773 2573
rect 1790 2556 1793 2613
rect 1790 2553 1797 2556
rect 1778 2466 1781 2526
rect 1762 2463 1781 2466
rect 1762 2286 1765 2463
rect 1786 2456 1789 2536
rect 1794 2533 1797 2553
rect 1794 2513 1797 2526
rect 1770 2453 1789 2456
rect 1770 2413 1773 2453
rect 1794 2436 1797 2506
rect 1790 2433 1797 2436
rect 1770 2353 1773 2386
rect 1790 2356 1793 2433
rect 1790 2353 1797 2356
rect 1770 2303 1773 2336
rect 1786 2303 1789 2336
rect 1794 2323 1797 2353
rect 1802 2316 1805 3136
rect 1818 3086 1821 3433
rect 1826 3363 1829 3426
rect 1826 3333 1829 3346
rect 1826 3133 1829 3306
rect 1834 3213 1837 3453
rect 1842 3373 1845 3513
rect 1866 3506 1869 3566
rect 1850 3433 1853 3506
rect 1862 3503 1869 3506
rect 1862 3426 1865 3503
rect 1874 3493 1877 3596
rect 1882 3483 1885 3646
rect 1890 3506 1893 3686
rect 1898 3586 1901 3616
rect 1914 3603 1917 3743
rect 1922 3683 1925 3756
rect 1930 3723 1933 3853
rect 1938 3746 1941 3906
rect 1946 3863 1949 4016
rect 1954 3976 1957 4043
rect 1978 4036 1981 4126
rect 1962 4033 1981 4036
rect 1962 3983 1965 4033
rect 1978 4003 1981 4016
rect 1954 3973 1989 3976
rect 1954 3943 1973 3946
rect 1954 3933 1957 3943
rect 1962 3856 1965 3936
rect 1970 3923 1973 3943
rect 1978 3906 1981 3936
rect 1954 3853 1965 3856
rect 1974 3903 1981 3906
rect 1946 3793 1949 3816
rect 1938 3743 1949 3746
rect 1938 3693 1941 3716
rect 1898 3583 1909 3586
rect 1898 3513 1901 3576
rect 1906 3563 1909 3583
rect 1914 3556 1917 3576
rect 1914 3553 1921 3556
rect 1906 3513 1909 3536
rect 1890 3503 1905 3506
rect 1862 3423 1869 3426
rect 1842 3333 1845 3356
rect 1842 3223 1845 3316
rect 1850 3293 1853 3416
rect 1858 3303 1861 3406
rect 1866 3313 1869 3423
rect 1874 3296 1877 3466
rect 1882 3403 1885 3416
rect 1890 3333 1893 3496
rect 1902 3446 1905 3503
rect 1918 3496 1921 3553
rect 1914 3493 1921 3496
rect 1902 3443 1909 3446
rect 1898 3413 1901 3426
rect 1898 3343 1901 3366
rect 1898 3326 1901 3336
rect 1906 3333 1909 3443
rect 1914 3333 1917 3493
rect 1930 3476 1933 3516
rect 1938 3493 1941 3626
rect 1946 3573 1949 3743
rect 1954 3566 1957 3853
rect 1974 3836 1977 3903
rect 1974 3833 1981 3836
rect 1978 3813 1981 3833
rect 1986 3813 1989 3973
rect 1994 3813 1997 3936
rect 2002 3806 2005 4313
rect 2018 4256 2021 4323
rect 2010 4253 2021 4256
rect 2010 4003 2013 4253
rect 2018 4223 2021 4236
rect 2018 4163 2021 4206
rect 2034 4203 2037 4316
rect 2058 4196 2061 4337
rect 2090 4256 2093 4326
rect 2090 4253 2101 4256
rect 2050 4193 2061 4196
rect 2018 4133 2021 4146
rect 2018 4103 2021 4126
rect 2026 4063 2029 4186
rect 2034 4113 2037 4136
rect 2042 4093 2045 4126
rect 2010 3933 2013 3956
rect 2018 3936 2021 4016
rect 2050 4006 2053 4193
rect 2066 4173 2069 4236
rect 2082 4203 2085 4216
rect 2066 4033 2069 4136
rect 2042 3996 2045 4006
rect 2050 4003 2069 4006
rect 2074 4003 2077 4016
rect 2090 4006 2093 4126
rect 2098 4113 2101 4253
rect 2106 4043 2109 4246
rect 2114 4143 2117 4337
rect 2138 4313 2189 4316
rect 2122 4203 2125 4286
rect 2138 4236 2141 4313
rect 2138 4233 2149 4236
rect 2130 4183 2133 4216
rect 2138 4193 2141 4206
rect 2146 4176 2149 4233
rect 2130 4173 2149 4176
rect 2130 4093 2133 4173
rect 2154 4166 2157 4296
rect 2162 4203 2165 4306
rect 2186 4276 2189 4313
rect 2162 4176 2165 4196
rect 2170 4183 2173 4216
rect 2178 4203 2181 4276
rect 2186 4273 2197 4276
rect 2186 4213 2189 4273
rect 2194 4193 2197 4206
rect 2210 4203 2213 4316
rect 2226 4283 2229 4340
rect 2242 4293 2245 4340
rect 2322 4303 2325 4340
rect 2250 4226 2253 4286
rect 2274 4256 2277 4296
rect 2282 4293 2317 4296
rect 2282 4273 2285 4293
rect 2274 4253 2281 4256
rect 2242 4223 2253 4226
rect 2162 4173 2173 4176
rect 2138 4163 2157 4166
rect 2114 4036 2117 4066
rect 2106 4033 2117 4036
rect 2082 4003 2093 4006
rect 2042 3993 2053 3996
rect 2018 3933 2029 3936
rect 2010 3913 2013 3926
rect 2018 3903 2021 3926
rect 1986 3803 2005 3806
rect 1986 3773 1989 3803
rect 2010 3796 2013 3816
rect 2018 3813 2021 3886
rect 1962 3743 1989 3746
rect 1962 3656 1965 3743
rect 1970 3733 1981 3736
rect 1970 3703 1973 3733
rect 1978 3716 1981 3726
rect 1986 3723 1989 3743
rect 1994 3734 1997 3796
rect 2002 3793 2013 3796
rect 2018 3793 2021 3806
rect 2002 3723 2005 3793
rect 2010 3716 2013 3736
rect 1978 3713 2013 3716
rect 1962 3653 1981 3656
rect 1962 3573 1965 3616
rect 1954 3563 1965 3566
rect 1946 3513 1949 3536
rect 1922 3473 1933 3476
rect 1922 3383 1925 3473
rect 1930 3413 1949 3416
rect 1930 3403 1933 3413
rect 1954 3403 1957 3546
rect 1962 3403 1965 3563
rect 1978 3533 1981 3653
rect 1970 3513 1973 3526
rect 1970 3413 1973 3506
rect 1978 3396 1981 3496
rect 1930 3373 1933 3396
rect 1962 3393 1981 3396
rect 1870 3293 1877 3296
rect 1858 3206 1861 3266
rect 1870 3226 1873 3293
rect 1882 3253 1885 3316
rect 1890 3306 1893 3326
rect 1898 3323 1917 3326
rect 1890 3303 1901 3306
rect 1930 3303 1933 3346
rect 1946 3333 1949 3356
rect 1954 3343 1957 3366
rect 1870 3223 1877 3226
rect 1834 3203 1845 3206
rect 1854 3203 1861 3206
rect 1874 3203 1877 3223
rect 1834 3123 1837 3203
rect 1854 3156 1857 3203
rect 1866 3183 1869 3196
rect 1882 3193 1885 3206
rect 1898 3186 1901 3303
rect 1914 3223 1933 3226
rect 1938 3223 1941 3256
rect 1914 3213 1917 3223
rect 1930 3216 1933 3223
rect 1922 3196 1925 3216
rect 1930 3213 1941 3216
rect 1938 3203 1941 3213
rect 1946 3196 1949 3226
rect 1954 3203 1957 3246
rect 1922 3193 1949 3196
rect 1962 3193 1965 3393
rect 1970 3363 1981 3366
rect 1970 3323 1973 3363
rect 1978 3306 1981 3326
rect 1974 3303 1981 3306
rect 1974 3236 1977 3303
rect 1970 3233 1977 3236
rect 1970 3213 1973 3233
rect 1890 3183 1901 3186
rect 1854 3153 1861 3156
rect 1842 3123 1845 3136
rect 1858 3133 1861 3153
rect 1866 3143 1869 3166
rect 1818 3083 1829 3086
rect 1810 3013 1813 3076
rect 1818 3003 1821 3036
rect 1826 2986 1829 3006
rect 1874 3003 1877 3086
rect 1890 3016 1893 3183
rect 1906 3143 1909 3166
rect 1938 3143 1941 3193
rect 1906 3083 1909 3136
rect 1914 3133 1933 3136
rect 1946 3133 1949 3166
rect 1954 3146 1957 3176
rect 1954 3143 1973 3146
rect 1978 3133 1981 3226
rect 1826 2983 1865 2986
rect 1818 2896 1821 2936
rect 1810 2893 1821 2896
rect 1810 2843 1813 2893
rect 1842 2886 1845 2926
rect 1818 2883 1845 2886
rect 1810 2716 1813 2816
rect 1818 2803 1821 2883
rect 1826 2813 1829 2846
rect 1834 2813 1845 2816
rect 1818 2723 1821 2746
rect 1826 2733 1829 2776
rect 1834 2756 1837 2813
rect 1850 2806 1853 2926
rect 1862 2886 1865 2983
rect 1882 2966 1885 3016
rect 1890 3013 1901 3016
rect 1874 2963 1885 2966
rect 1890 2963 1893 3006
rect 1898 2946 1901 3013
rect 1914 3003 1917 3036
rect 1938 3013 1941 3096
rect 1946 2976 1949 3126
rect 1962 3123 1973 3126
rect 1962 3083 1965 3123
rect 1986 3106 1989 3696
rect 2018 3686 2021 3776
rect 1994 3683 2021 3686
rect 1994 3613 1997 3683
rect 2026 3676 2029 3926
rect 2034 3906 2037 3926
rect 2042 3913 2045 3936
rect 2050 3933 2053 3993
rect 2058 3923 2061 3956
rect 2066 3933 2069 3966
rect 2066 3906 2069 3926
rect 2034 3903 2069 3906
rect 2074 3903 2077 3956
rect 2082 3933 2085 4003
rect 2098 3966 2101 4016
rect 2106 4003 2109 4033
rect 2122 4023 2125 4046
rect 2090 3963 2101 3966
rect 2090 3923 2093 3963
rect 2098 3926 2101 3936
rect 2106 3933 2109 3956
rect 2098 3923 2109 3926
rect 2034 3813 2037 3836
rect 2042 3803 2045 3866
rect 2050 3823 2061 3826
rect 2050 3786 2053 3816
rect 2034 3783 2053 3786
rect 2034 3736 2037 3783
rect 2042 3743 2045 3756
rect 2034 3733 2045 3736
rect 2010 3673 2029 3676
rect 2002 3536 2005 3616
rect 2010 3603 2013 3673
rect 2034 3613 2037 3726
rect 2042 3683 2045 3733
rect 2050 3723 2053 3776
rect 2058 3753 2061 3816
rect 2066 3793 2069 3903
rect 2074 3773 2077 3886
rect 2082 3823 2085 3836
rect 2090 3766 2093 3916
rect 2114 3876 2117 4016
rect 2122 3983 2125 4006
rect 2138 4003 2141 4163
rect 2162 4156 2165 4166
rect 2146 4153 2165 4156
rect 2146 4123 2149 4153
rect 2154 4133 2157 4146
rect 2170 4143 2173 4173
rect 2242 4166 2245 4223
rect 2178 4163 2213 4166
rect 2242 4163 2253 4166
rect 2162 4133 2173 4136
rect 2154 4103 2157 4126
rect 2162 4123 2165 4133
rect 2146 3966 2149 4096
rect 2098 3873 2117 3876
rect 2122 3963 2149 3966
rect 2098 3803 2101 3873
rect 2122 3836 2125 3963
rect 2130 3916 2133 3926
rect 2146 3923 2149 3936
rect 2154 3933 2157 4016
rect 2154 3916 2157 3926
rect 2130 3913 2157 3916
rect 2110 3833 2125 3836
rect 2066 3763 2093 3766
rect 2066 3736 2069 3763
rect 2058 3733 2069 3736
rect 2058 3696 2061 3733
rect 2066 3703 2069 3726
rect 2050 3693 2061 3696
rect 2074 3693 2077 3736
rect 2082 3723 2085 3756
rect 2098 3723 2101 3796
rect 2110 3766 2113 3833
rect 2106 3763 2113 3766
rect 2106 3716 2109 3763
rect 2114 3723 2117 3746
rect 2082 3713 2093 3716
rect 2098 3713 2109 3716
rect 2050 3623 2053 3693
rect 2042 3613 2053 3616
rect 2018 3603 2029 3606
rect 2018 3573 2021 3603
rect 2034 3596 2037 3606
rect 2042 3603 2045 3613
rect 2026 3593 2037 3596
rect 1994 3413 1997 3536
rect 2002 3533 2013 3536
rect 2002 3483 2005 3526
rect 2002 3406 2005 3426
rect 2010 3413 2013 3533
rect 2018 3433 2021 3516
rect 1994 3403 2005 3406
rect 2018 3403 2021 3426
rect 1994 3223 1997 3403
rect 2002 3333 2005 3366
rect 2010 3323 2013 3346
rect 2018 3333 2021 3396
rect 2026 3316 2029 3593
rect 2034 3453 2037 3576
rect 2050 3563 2053 3606
rect 2042 3493 2045 3546
rect 2058 3533 2061 3686
rect 2082 3663 2085 3713
rect 2066 3553 2069 3606
rect 2050 3523 2069 3526
rect 2074 3486 2077 3546
rect 2082 3543 2085 3576
rect 2090 3536 2093 3656
rect 2098 3613 2101 3713
rect 2114 3703 2117 3716
rect 2098 3563 2101 3596
rect 2050 3483 2077 3486
rect 2034 3353 2037 3416
rect 2042 3413 2045 3426
rect 2050 3403 2053 3483
rect 2042 3323 2045 3366
rect 2002 3263 2005 3316
rect 2026 3313 2045 3316
rect 2058 3313 2061 3456
rect 2066 3403 2069 3476
rect 2066 3316 2069 3396
rect 2074 3323 2077 3483
rect 2082 3533 2093 3536
rect 2082 3466 2085 3533
rect 2090 3523 2101 3526
rect 2082 3463 2093 3466
rect 2106 3463 2109 3666
rect 2114 3613 2117 3686
rect 2122 3573 2125 3826
rect 2130 3803 2133 3846
rect 2138 3813 2141 3913
rect 2146 3796 2149 3906
rect 2162 3876 2165 4116
rect 2170 4103 2173 4126
rect 2170 4013 2173 4046
rect 2170 3903 2173 3976
rect 2178 3936 2181 4163
rect 2186 4133 2189 4146
rect 2194 4143 2205 4146
rect 2194 4103 2197 4143
rect 2202 4126 2205 4136
rect 2210 4133 2213 4163
rect 2226 4133 2229 4146
rect 2250 4143 2253 4163
rect 2258 4156 2261 4216
rect 2278 4186 2281 4253
rect 2290 4213 2293 4286
rect 2298 4203 2301 4276
rect 2314 4236 2317 4293
rect 2314 4233 2325 4236
rect 2274 4183 2281 4186
rect 2306 4183 2309 4216
rect 2274 4163 2277 4183
rect 2258 4153 2301 4156
rect 2202 4123 2213 4126
rect 2218 4106 2221 4126
rect 2210 4103 2221 4106
rect 2210 4026 2213 4103
rect 2210 4023 2221 4026
rect 2186 3953 2189 4016
rect 2202 4003 2213 4006
rect 2218 3996 2221 4023
rect 2210 3993 2221 3996
rect 2178 3933 2197 3936
rect 2210 3933 2213 3993
rect 2226 3986 2229 4126
rect 2242 4066 2245 4126
rect 2250 4086 2253 4136
rect 2266 4133 2269 4146
rect 2258 4123 2269 4126
rect 2258 4093 2261 4123
rect 2274 4086 2277 4126
rect 2250 4083 2277 4086
rect 2234 4063 2245 4066
rect 2218 3983 2229 3986
rect 2154 3873 2165 3876
rect 2154 3803 2157 3873
rect 2130 3793 2149 3796
rect 2162 3793 2165 3866
rect 2170 3803 2173 3836
rect 2178 3813 2181 3926
rect 2130 3706 2133 3793
rect 2186 3756 2189 3826
rect 2194 3776 2197 3933
rect 2210 3893 2213 3926
rect 2202 3786 2205 3816
rect 2210 3793 2213 3836
rect 2202 3783 2213 3786
rect 2194 3773 2205 3776
rect 2170 3753 2189 3756
rect 2138 3733 2141 3746
rect 2138 3723 2149 3726
rect 2130 3703 2141 3706
rect 2138 3646 2141 3703
rect 2130 3643 2141 3646
rect 2130 3603 2133 3643
rect 2138 3623 2157 3626
rect 2138 3613 2141 3623
rect 2154 3616 2157 3623
rect 2138 3583 2141 3606
rect 2114 3526 2117 3546
rect 2114 3523 2133 3526
rect 2122 3483 2125 3516
rect 2146 3473 2149 3616
rect 2154 3613 2165 3616
rect 2162 3603 2165 3613
rect 2154 3483 2157 3576
rect 2162 3533 2165 3546
rect 2170 3526 2173 3753
rect 2178 3723 2181 3736
rect 2186 3693 2189 3746
rect 2178 3613 2181 3626
rect 2186 3613 2189 3626
rect 2194 3533 2197 3766
rect 2202 3733 2205 3773
rect 2210 3763 2213 3783
rect 2218 3746 2221 3983
rect 2226 3933 2229 3976
rect 2234 3923 2237 4006
rect 2250 4003 2253 4066
rect 2274 4026 2277 4046
rect 2282 4036 2285 4136
rect 2290 4043 2293 4146
rect 2298 4133 2301 4153
rect 2314 4146 2317 4206
rect 2322 4163 2325 4233
rect 2306 4143 2317 4146
rect 2306 4133 2309 4143
rect 2314 4126 2317 4136
rect 2322 4133 2325 4146
rect 2306 4093 2309 4126
rect 2314 4123 2325 4126
rect 2330 4066 2333 4296
rect 2346 4203 2349 4316
rect 2362 4246 2365 4340
rect 2362 4243 2373 4246
rect 2370 4203 2373 4243
rect 2346 4133 2349 4196
rect 2362 4133 2365 4146
rect 2338 4113 2341 4126
rect 2330 4063 2341 4066
rect 2298 4053 2333 4056
rect 2282 4033 2293 4036
rect 2274 4023 2285 4026
rect 2274 3973 2277 4016
rect 2242 3933 2261 3936
rect 2250 3893 2253 3926
rect 2258 3923 2261 3933
rect 2242 3883 2253 3886
rect 2250 3866 2253 3883
rect 2246 3863 2253 3866
rect 2226 3823 2229 3836
rect 2234 3813 2237 3826
rect 2210 3743 2221 3746
rect 2210 3723 2213 3743
rect 2226 3736 2229 3766
rect 2246 3756 2249 3863
rect 2258 3803 2261 3836
rect 2266 3823 2269 3926
rect 2274 3813 2277 3866
rect 2282 3823 2285 4023
rect 2290 3933 2293 4033
rect 2298 3933 2301 4053
rect 2330 4043 2333 4053
rect 2330 4003 2333 4016
rect 2338 4003 2341 4063
rect 2354 4043 2357 4126
rect 2370 4123 2373 4136
rect 2378 4133 2381 4306
rect 2410 4293 2413 4340
rect 2426 4286 2429 4340
rect 2562 4337 2597 4340
rect 2394 4283 2429 4286
rect 2394 4273 2397 4283
rect 2434 4276 2437 4306
rect 2426 4273 2437 4276
rect 2378 4106 2381 4126
rect 2386 4123 2389 4196
rect 2394 4176 2397 4216
rect 2426 4213 2429 4273
rect 2394 4173 2421 4176
rect 2402 4123 2405 4136
rect 2418 4133 2421 4173
rect 2410 4116 2413 4126
rect 2426 4123 2429 4196
rect 2442 4193 2445 4316
rect 2434 4126 2437 4136
rect 2442 4133 2453 4136
rect 2434 4123 2445 4126
rect 2450 4116 2453 4133
rect 2458 4123 2461 4146
rect 2466 4133 2469 4276
rect 2474 4216 2477 4296
rect 2474 4213 2481 4216
rect 2478 4156 2481 4213
rect 2490 4176 2493 4216
rect 2522 4213 2525 4276
rect 2530 4223 2557 4226
rect 2530 4213 2533 4223
rect 2538 4213 2549 4216
rect 2554 4213 2557 4223
rect 2490 4173 2501 4176
rect 2474 4153 2481 4156
rect 2410 4113 2453 4116
rect 2370 4103 2381 4106
rect 2370 4086 2373 4103
rect 2450 4096 2453 4113
rect 2366 4083 2373 4086
rect 2446 4093 2453 4096
rect 2474 4093 2477 4153
rect 2482 4103 2485 4136
rect 2498 4133 2501 4173
rect 2522 4146 2525 4206
rect 2530 4203 2541 4206
rect 2490 4116 2493 4126
rect 2506 4123 2509 4146
rect 2522 4143 2541 4146
rect 2514 4126 2517 4136
rect 2522 4133 2533 4136
rect 2514 4123 2525 4126
rect 2530 4116 2533 4133
rect 2490 4113 2533 4116
rect 2366 4026 2369 4083
rect 2378 4053 2413 4056
rect 2366 4023 2373 4026
rect 2314 3926 2317 3986
rect 2322 3943 2341 3946
rect 2322 3933 2325 3943
rect 2298 3826 2301 3926
rect 2314 3923 2325 3926
rect 2330 3893 2333 3936
rect 2338 3923 2341 3943
rect 2346 3933 2349 4016
rect 2354 3926 2357 3956
rect 2362 3933 2365 3976
rect 2370 3943 2373 4023
rect 2378 4013 2381 4053
rect 2386 4003 2389 4046
rect 2410 4026 2413 4053
rect 2446 4036 2449 4093
rect 2442 4033 2449 4036
rect 2410 4023 2433 4026
rect 2394 4003 2397 4016
rect 2410 4013 2413 4023
rect 2418 4006 2421 4016
rect 2402 4003 2421 4006
rect 2354 3923 2365 3926
rect 2290 3823 2301 3826
rect 2306 3823 2309 3846
rect 2330 3833 2341 3836
rect 2290 3806 2293 3823
rect 2298 3813 2309 3816
rect 2266 3803 2293 3806
rect 2246 3753 2253 3756
rect 2218 3733 2229 3736
rect 2242 3726 2245 3736
rect 2218 3676 2221 3726
rect 2226 3683 2229 3726
rect 2234 3723 2245 3726
rect 2234 3676 2237 3723
rect 2218 3673 2237 3676
rect 2202 3603 2205 3616
rect 2210 3526 2213 3626
rect 2234 3603 2237 3656
rect 2242 3603 2245 3716
rect 2162 3523 2173 3526
rect 2194 3523 2213 3526
rect 2082 3413 2085 3456
rect 2082 3323 2085 3406
rect 2090 3376 2093 3463
rect 2130 3453 2141 3456
rect 2114 3433 2125 3436
rect 2098 3406 2101 3416
rect 2114 3406 2117 3433
rect 2098 3403 2117 3406
rect 2098 3386 2101 3396
rect 2114 3393 2117 3403
rect 2098 3383 2109 3386
rect 2090 3373 2101 3376
rect 2098 3343 2101 3373
rect 2106 3366 2109 3383
rect 2106 3363 2125 3366
rect 2106 3343 2109 3356
rect 2122 3353 2125 3363
rect 2130 3336 2133 3436
rect 2138 3423 2141 3453
rect 2162 3446 2165 3523
rect 2170 3513 2181 3516
rect 2210 3506 2213 3523
rect 2206 3503 2213 3506
rect 2178 3473 2189 3476
rect 2154 3443 2165 3446
rect 2138 3363 2141 3406
rect 2138 3346 2141 3356
rect 2154 3353 2157 3443
rect 2138 3343 2149 3346
rect 2126 3333 2133 3336
rect 2066 3313 2077 3316
rect 2018 3213 2037 3216
rect 2018 3203 2021 3213
rect 2042 3203 2045 3313
rect 2018 3173 2021 3196
rect 2050 3166 2053 3216
rect 2066 3203 2069 3246
rect 2074 3176 2077 3313
rect 2098 3306 2101 3326
rect 2098 3303 2105 3306
rect 2114 3303 2117 3316
rect 2082 3276 2085 3296
rect 2082 3273 2093 3276
rect 2082 3186 2085 3266
rect 2090 3243 2093 3273
rect 2102 3226 2105 3303
rect 2126 3236 2129 3333
rect 2138 3263 2141 3326
rect 2146 3323 2149 3343
rect 2154 3323 2157 3336
rect 2162 3333 2165 3436
rect 2170 3253 2173 3466
rect 2178 3423 2181 3436
rect 2178 3353 2181 3396
rect 2126 3233 2133 3236
rect 2098 3223 2105 3226
rect 2090 3193 2093 3206
rect 2098 3203 2101 3223
rect 2106 3193 2109 3206
rect 2122 3193 2125 3216
rect 2082 3183 2093 3186
rect 2074 3173 2081 3176
rect 1994 3113 1997 3126
rect 2002 3123 2005 3166
rect 2050 3163 2069 3166
rect 1986 3103 1997 3106
rect 1954 3016 1957 3036
rect 1954 3013 1961 3016
rect 1922 2973 1949 2976
rect 1898 2943 1917 2946
rect 1882 2886 1885 2936
rect 1890 2923 1901 2926
rect 1862 2883 1869 2886
rect 1842 2803 1853 2806
rect 1858 2803 1861 2866
rect 1834 2753 1845 2756
rect 1842 2733 1845 2753
rect 1810 2713 1829 2716
rect 1810 2703 1821 2706
rect 1810 2606 1813 2616
rect 1818 2613 1821 2636
rect 1810 2603 1821 2606
rect 1810 2583 1813 2596
rect 1818 2546 1821 2603
rect 1826 2576 1829 2713
rect 1834 2686 1837 2726
rect 1842 2703 1845 2726
rect 1850 2723 1853 2766
rect 1866 2756 1869 2883
rect 1874 2883 1885 2886
rect 1874 2773 1877 2883
rect 1898 2856 1901 2923
rect 1906 2873 1909 2936
rect 1914 2906 1917 2943
rect 1922 2923 1925 2973
rect 1958 2946 1961 3013
rect 1954 2943 1961 2946
rect 1914 2903 1921 2906
rect 1898 2853 1909 2856
rect 1882 2766 1885 2816
rect 1890 2803 1893 2826
rect 1898 2813 1901 2846
rect 1882 2763 1901 2766
rect 1858 2753 1869 2756
rect 1834 2683 1853 2686
rect 1834 2603 1837 2676
rect 1842 2613 1845 2626
rect 1826 2573 1845 2576
rect 1810 2543 1821 2546
rect 1818 2526 1821 2536
rect 1810 2503 1813 2526
rect 1818 2523 1829 2526
rect 1818 2496 1821 2516
rect 1810 2493 1821 2496
rect 1810 2396 1813 2493
rect 1818 2413 1821 2476
rect 1810 2393 1821 2396
rect 1810 2333 1813 2376
rect 1762 2283 1781 2286
rect 1762 2213 1773 2216
rect 1778 2206 1781 2283
rect 1794 2233 1797 2316
rect 1802 2313 1809 2316
rect 1786 2216 1789 2226
rect 1806 2216 1809 2313
rect 1818 2233 1821 2393
rect 1826 2383 1829 2523
rect 1834 2503 1837 2566
rect 1826 2343 1829 2356
rect 1834 2333 1837 2436
rect 1842 2406 1845 2573
rect 1850 2563 1853 2683
rect 1858 2546 1861 2753
rect 1850 2543 1861 2546
rect 1850 2523 1853 2543
rect 1866 2536 1869 2706
rect 1874 2686 1877 2756
rect 1898 2736 1901 2763
rect 1906 2753 1909 2853
rect 1918 2826 1921 2903
rect 1938 2866 1941 2926
rect 1946 2913 1949 2936
rect 1930 2863 1941 2866
rect 1930 2833 1933 2863
rect 1954 2856 1957 2943
rect 1938 2853 1957 2856
rect 1914 2823 1921 2826
rect 1914 2756 1917 2823
rect 1922 2773 1925 2806
rect 1914 2753 1921 2756
rect 1898 2733 1909 2736
rect 1874 2683 1893 2686
rect 1874 2666 1877 2676
rect 1890 2673 1893 2683
rect 1898 2666 1901 2726
rect 1874 2663 1901 2666
rect 1906 2656 1909 2733
rect 1918 2686 1921 2753
rect 1938 2723 1941 2853
rect 1962 2833 1965 2926
rect 1970 2923 1973 2966
rect 1994 2963 1997 3103
rect 2010 3093 2013 3136
rect 2018 3113 2021 3146
rect 2034 3133 2037 3146
rect 2042 3123 2045 3136
rect 2002 3003 2005 3046
rect 1978 2873 1981 2936
rect 1994 2856 1997 2926
rect 1986 2853 1997 2856
rect 1962 2813 1965 2826
rect 1978 2806 1981 2826
rect 1962 2803 1981 2806
rect 1946 2716 1949 2756
rect 1938 2713 1949 2716
rect 1918 2683 1933 2686
rect 1890 2653 1909 2656
rect 1858 2533 1869 2536
rect 1874 2516 1877 2616
rect 1882 2583 1885 2606
rect 1850 2493 1853 2506
rect 1850 2413 1853 2426
rect 1858 2413 1861 2516
rect 1870 2513 1877 2516
rect 1882 2513 1885 2566
rect 1842 2403 1853 2406
rect 1850 2386 1853 2403
rect 1870 2386 1873 2513
rect 1882 2433 1885 2506
rect 1850 2383 1857 2386
rect 1870 2383 1877 2386
rect 1842 2333 1845 2366
rect 1854 2326 1857 2383
rect 1874 2366 1877 2383
rect 1882 2373 1885 2426
rect 1874 2363 1885 2366
rect 1874 2333 1877 2356
rect 1842 2303 1845 2326
rect 1850 2323 1857 2326
rect 1850 2256 1853 2323
rect 1858 2263 1861 2306
rect 1850 2253 1861 2256
rect 1826 2216 1829 2246
rect 1842 2223 1845 2246
rect 1786 2213 1797 2216
rect 1806 2213 1813 2216
rect 1762 2183 1765 2206
rect 1770 2203 1781 2206
rect 1770 2143 1773 2203
rect 1786 2183 1789 2206
rect 1794 2166 1797 2213
rect 1786 2163 1797 2166
rect 1786 2156 1789 2163
rect 1810 2156 1813 2213
rect 1778 2153 1789 2156
rect 1794 2153 1813 2156
rect 1822 2213 1829 2216
rect 1762 2123 1765 2136
rect 1762 2013 1765 2036
rect 1770 2023 1773 2136
rect 1754 1933 1765 1936
rect 1754 1916 1757 1933
rect 1770 1926 1773 2016
rect 1738 1913 1757 1916
rect 1762 1923 1773 1926
rect 1738 1906 1741 1913
rect 1714 1903 1741 1906
rect 1706 1893 1717 1896
rect 1706 1763 1709 1816
rect 1714 1786 1717 1893
rect 1714 1783 1725 1786
rect 1722 1733 1725 1783
rect 1690 1713 1697 1716
rect 1682 1633 1685 1656
rect 1634 1563 1645 1566
rect 1642 1543 1645 1563
rect 1618 1483 1629 1486
rect 1586 1413 1605 1416
rect 1610 1413 1613 1426
rect 1586 1393 1589 1413
rect 1594 1373 1597 1406
rect 1602 1403 1621 1406
rect 1530 1183 1533 1206
rect 1546 1163 1549 1216
rect 1562 1213 1569 1216
rect 1554 1143 1557 1206
rect 1566 1166 1569 1213
rect 1578 1203 1581 1226
rect 1566 1163 1573 1166
rect 1570 1153 1573 1163
rect 1578 1136 1581 1186
rect 1586 1143 1589 1366
rect 1602 1333 1605 1403
rect 1610 1373 1613 1403
rect 1602 1213 1605 1286
rect 1610 1253 1613 1336
rect 1618 1223 1621 1336
rect 1522 1013 1525 1106
rect 1538 1076 1541 1126
rect 1534 1073 1541 1076
rect 1554 1076 1557 1136
rect 1578 1133 1589 1136
rect 1554 1073 1561 1076
rect 1534 1026 1537 1073
rect 1534 1023 1541 1026
rect 1522 996 1525 1006
rect 1538 1003 1541 1023
rect 1546 1013 1549 1066
rect 1522 993 1549 996
rect 1522 933 1525 946
rect 1522 923 1541 926
rect 1522 803 1525 906
rect 1530 853 1533 896
rect 1506 783 1525 786
rect 1466 763 1485 766
rect 1466 733 1469 746
rect 1454 723 1461 726
rect 1402 683 1413 686
rect 1434 713 1445 716
rect 1434 646 1437 713
rect 1426 643 1437 646
rect 1386 633 1393 636
rect 1346 503 1349 536
rect 1362 533 1365 586
rect 1354 523 1365 526
rect 1354 403 1357 466
rect 1370 446 1373 606
rect 1386 556 1389 633
rect 1394 563 1397 616
rect 1410 586 1413 606
rect 1418 603 1421 636
rect 1426 613 1429 643
rect 1434 593 1437 606
rect 1442 586 1445 616
rect 1450 603 1453 626
rect 1458 603 1461 723
rect 1410 583 1445 586
rect 1458 583 1461 596
rect 1418 556 1421 576
rect 1378 533 1381 556
rect 1386 553 1397 556
rect 1370 443 1381 446
rect 1330 386 1333 403
rect 1330 383 1349 386
rect 1314 373 1341 376
rect 1290 323 1301 326
rect 1314 316 1317 336
rect 1330 333 1333 346
rect 1338 326 1341 373
rect 1346 333 1349 383
rect 1354 333 1357 376
rect 1338 323 1357 326
rect 1314 313 1333 316
rect 1314 256 1317 296
rect 1314 253 1321 256
rect 1298 193 1301 216
rect 1318 176 1321 253
rect 1330 236 1333 313
rect 1330 233 1341 236
rect 1330 183 1333 216
rect 1338 203 1341 233
rect 1346 213 1349 296
rect 1354 286 1357 323
rect 1378 303 1381 443
rect 1386 403 1389 536
rect 1394 386 1397 553
rect 1410 553 1421 556
rect 1410 466 1413 553
rect 1410 463 1421 466
rect 1390 383 1397 386
rect 1354 283 1381 286
rect 1370 193 1373 206
rect 1378 203 1381 283
rect 1390 266 1393 383
rect 1402 353 1405 416
rect 1418 413 1421 463
rect 1426 456 1429 583
rect 1434 513 1437 536
rect 1442 516 1445 526
rect 1450 523 1453 536
rect 1466 533 1477 536
rect 1442 513 1453 516
rect 1426 453 1437 456
rect 1434 396 1437 453
rect 1450 403 1453 513
rect 1482 493 1485 763
rect 1498 716 1501 756
rect 1522 733 1525 783
rect 1506 723 1517 726
rect 1498 713 1509 716
rect 1490 593 1493 616
rect 1498 613 1501 636
rect 1506 606 1509 713
rect 1530 673 1533 716
rect 1530 623 1533 646
rect 1538 616 1541 726
rect 1530 613 1541 616
rect 1530 606 1533 613
rect 1498 603 1509 606
rect 1514 603 1533 606
rect 1490 426 1493 446
rect 1458 423 1477 426
rect 1458 413 1461 423
rect 1466 403 1469 416
rect 1474 403 1477 423
rect 1486 423 1493 426
rect 1434 393 1445 396
rect 1418 336 1421 386
rect 1390 263 1397 266
rect 1394 243 1397 263
rect 1386 203 1389 226
rect 1402 216 1405 336
rect 1418 333 1429 336
rect 1410 306 1413 326
rect 1418 323 1429 326
rect 1410 303 1421 306
rect 1434 286 1437 326
rect 1398 213 1405 216
rect 1426 283 1437 286
rect 1314 173 1321 176
rect 1298 113 1301 136
rect 1306 116 1309 126
rect 1314 123 1317 173
rect 1398 156 1401 213
rect 1398 153 1405 156
rect 1322 133 1325 146
rect 1330 123 1333 136
rect 1338 116 1341 136
rect 1378 123 1381 136
rect 1306 113 1341 116
rect 1402 113 1405 153
rect 1410 143 1413 206
rect 1418 123 1421 196
rect 1426 133 1429 283
rect 1434 203 1437 216
rect 1442 213 1445 393
rect 1450 303 1453 336
rect 1458 333 1461 396
rect 1486 356 1489 423
rect 1498 373 1501 603
rect 1546 576 1549 993
rect 1558 946 1561 1073
rect 1570 956 1573 1026
rect 1578 1003 1581 1133
rect 1594 1123 1597 1206
rect 1610 1163 1613 1206
rect 1586 1036 1589 1076
rect 1602 1073 1605 1146
rect 1618 1086 1621 1216
rect 1626 1093 1629 1483
rect 1634 1363 1637 1416
rect 1642 1333 1645 1536
rect 1650 1506 1653 1566
rect 1658 1546 1661 1623
rect 1658 1543 1669 1546
rect 1658 1523 1661 1536
rect 1666 1523 1669 1543
rect 1674 1523 1677 1616
rect 1650 1503 1661 1506
rect 1658 1436 1661 1503
rect 1650 1433 1661 1436
rect 1650 1376 1653 1433
rect 1658 1413 1669 1416
rect 1674 1413 1677 1426
rect 1666 1396 1669 1406
rect 1658 1393 1669 1396
rect 1674 1376 1677 1396
rect 1650 1373 1661 1376
rect 1658 1326 1661 1373
rect 1634 1283 1637 1326
rect 1650 1323 1661 1326
rect 1670 1373 1677 1376
rect 1634 1223 1637 1256
rect 1634 1153 1637 1216
rect 1642 1203 1645 1236
rect 1634 1123 1637 1136
rect 1610 1083 1621 1086
rect 1586 1033 1597 1036
rect 1570 953 1581 956
rect 1558 943 1565 946
rect 1554 833 1557 936
rect 1562 903 1565 943
rect 1570 923 1573 946
rect 1578 896 1581 953
rect 1586 933 1589 986
rect 1594 923 1597 1033
rect 1610 1023 1613 1083
rect 1602 993 1605 1016
rect 1610 986 1613 1006
rect 1618 993 1621 1046
rect 1626 1003 1629 1076
rect 1634 1013 1637 1036
rect 1610 983 1637 986
rect 1562 893 1581 896
rect 1562 826 1565 893
rect 1602 876 1605 936
rect 1610 923 1613 966
rect 1618 933 1621 946
rect 1634 936 1637 983
rect 1626 933 1637 936
rect 1558 823 1565 826
rect 1570 873 1605 876
rect 1558 756 1561 823
rect 1570 813 1573 873
rect 1602 813 1605 836
rect 1610 813 1613 826
rect 1618 796 1621 836
rect 1554 753 1561 756
rect 1614 793 1621 796
rect 1554 733 1557 753
rect 1578 733 1597 736
rect 1554 673 1557 696
rect 1538 573 1549 576
rect 1538 533 1541 573
rect 1554 563 1557 646
rect 1562 623 1565 716
rect 1562 553 1565 616
rect 1570 603 1573 726
rect 1578 693 1581 733
rect 1578 593 1581 626
rect 1530 513 1533 526
rect 1578 523 1581 536
rect 1586 503 1589 726
rect 1594 683 1597 716
rect 1602 703 1605 726
rect 1594 623 1597 676
rect 1614 636 1617 793
rect 1602 633 1617 636
rect 1506 386 1509 486
rect 1522 403 1525 466
rect 1546 446 1549 496
rect 1594 486 1597 616
rect 1590 483 1597 486
rect 1546 443 1557 446
rect 1554 396 1557 443
rect 1590 426 1593 483
rect 1602 463 1605 633
rect 1626 626 1629 926
rect 1634 913 1637 933
rect 1642 856 1645 1146
rect 1650 1123 1653 1323
rect 1670 1286 1673 1373
rect 1670 1283 1677 1286
rect 1650 976 1653 1036
rect 1658 1023 1661 1216
rect 1666 1203 1669 1266
rect 1674 1133 1677 1283
rect 1682 1126 1685 1626
rect 1694 1586 1697 1713
rect 1706 1613 1709 1726
rect 1730 1716 1733 1856
rect 1722 1713 1733 1716
rect 1690 1583 1697 1586
rect 1690 1546 1693 1583
rect 1698 1556 1701 1566
rect 1722 1563 1725 1713
rect 1698 1553 1717 1556
rect 1690 1543 1709 1546
rect 1690 1483 1693 1536
rect 1690 1413 1693 1436
rect 1690 1323 1693 1406
rect 1698 1316 1701 1406
rect 1706 1393 1709 1543
rect 1714 1533 1717 1553
rect 1722 1446 1725 1546
rect 1730 1523 1733 1636
rect 1738 1623 1741 1736
rect 1746 1716 1749 1766
rect 1754 1733 1757 1906
rect 1746 1713 1753 1716
rect 1750 1646 1753 1713
rect 1746 1643 1753 1646
rect 1746 1533 1749 1643
rect 1762 1636 1765 1923
rect 1770 1813 1773 1916
rect 1770 1723 1773 1756
rect 1770 1653 1773 1716
rect 1762 1633 1769 1636
rect 1754 1613 1757 1626
rect 1722 1443 1733 1446
rect 1730 1406 1733 1443
rect 1738 1423 1741 1496
rect 1714 1396 1717 1406
rect 1730 1403 1741 1406
rect 1746 1403 1749 1526
rect 1754 1486 1757 1606
rect 1766 1546 1769 1633
rect 1778 1603 1781 2153
rect 1786 1943 1789 2146
rect 1794 2033 1797 2153
rect 1822 2146 1825 2213
rect 1834 2146 1837 2216
rect 1802 2133 1805 2146
rect 1822 2143 1829 2146
rect 1834 2143 1845 2146
rect 1810 2046 1813 2126
rect 1826 2106 1829 2143
rect 1822 2103 1829 2106
rect 1822 2046 1825 2103
rect 1834 2083 1837 2136
rect 1842 2123 1845 2143
rect 1850 2063 1853 2216
rect 1802 2043 1813 2046
rect 1818 2043 1825 2046
rect 1794 2013 1797 2026
rect 1802 2006 1805 2043
rect 1794 2003 1805 2006
rect 1786 1896 1789 1926
rect 1794 1916 1797 1956
rect 1810 1936 1813 1956
rect 1802 1933 1813 1936
rect 1810 1916 1813 1926
rect 1794 1913 1813 1916
rect 1786 1893 1797 1896
rect 1794 1836 1797 1893
rect 1794 1833 1801 1836
rect 1798 1766 1801 1833
rect 1794 1763 1801 1766
rect 1794 1746 1797 1763
rect 1794 1743 1805 1746
rect 1802 1733 1805 1743
rect 1810 1726 1813 1896
rect 1762 1543 1769 1546
rect 1762 1523 1765 1543
rect 1770 1493 1773 1526
rect 1754 1483 1773 1486
rect 1714 1393 1725 1396
rect 1690 1313 1701 1316
rect 1690 1213 1693 1313
rect 1698 1296 1701 1313
rect 1698 1293 1709 1296
rect 1714 1276 1717 1336
rect 1738 1316 1741 1403
rect 1754 1396 1757 1406
rect 1746 1393 1757 1396
rect 1762 1393 1765 1416
rect 1770 1386 1773 1483
rect 1778 1396 1781 1536
rect 1786 1413 1789 1726
rect 1794 1723 1813 1726
rect 1794 1603 1797 1723
rect 1802 1613 1805 1666
rect 1818 1653 1821 2043
rect 1826 1986 1829 2036
rect 1834 1996 1837 2016
rect 1842 2003 1845 2026
rect 1850 2013 1853 2056
rect 1834 1993 1845 1996
rect 1826 1983 1837 1986
rect 1826 1933 1829 1976
rect 1834 1926 1837 1983
rect 1826 1923 1837 1926
rect 1826 1746 1829 1923
rect 1834 1756 1837 1916
rect 1842 1853 1845 1993
rect 1850 1933 1853 1946
rect 1850 1813 1853 1926
rect 1842 1763 1845 1806
rect 1858 1786 1861 2253
rect 1866 2196 1869 2326
rect 1882 2323 1885 2363
rect 1890 2276 1893 2653
rect 1914 2636 1917 2676
rect 1898 2633 1917 2636
rect 1898 2503 1901 2633
rect 1914 2613 1917 2626
rect 1922 2616 1925 2636
rect 1930 2623 1933 2683
rect 1938 2633 1941 2713
rect 1954 2706 1957 2726
rect 1946 2703 1957 2706
rect 1962 2633 1965 2803
rect 1986 2786 1989 2853
rect 1970 2783 1989 2786
rect 1922 2613 1933 2616
rect 1946 2613 1957 2616
rect 1962 2613 1965 2626
rect 1906 2563 1909 2606
rect 1922 2583 1925 2606
rect 1930 2576 1933 2613
rect 1970 2606 1973 2783
rect 1978 2696 1981 2776
rect 1994 2733 1997 2776
rect 2002 2766 2005 2936
rect 2010 2773 2013 3086
rect 2058 3073 2061 3136
rect 2066 3123 2069 3163
rect 2078 3066 2081 3173
rect 2090 3153 2093 3183
rect 2130 3136 2133 3233
rect 2138 3216 2141 3246
rect 2138 3213 2157 3216
rect 2090 3116 2093 3136
rect 2106 3123 2109 3136
rect 2122 3126 2125 3136
rect 2130 3133 2141 3136
rect 2122 3123 2133 3126
rect 2122 3116 2125 3123
rect 2090 3113 2125 3116
rect 2018 2943 2021 3066
rect 2078 3063 2085 3066
rect 2018 2913 2021 2926
rect 2018 2813 2021 2826
rect 2026 2813 2029 3016
rect 2034 3013 2045 3016
rect 2034 2933 2037 3013
rect 2066 3003 2069 3036
rect 2074 3013 2077 3046
rect 2002 2763 2013 2766
rect 2010 2753 2013 2763
rect 1978 2693 1985 2696
rect 1982 2646 1985 2693
rect 1994 2676 1997 2726
rect 2026 2723 2029 2776
rect 1994 2673 2013 2676
rect 1982 2643 1989 2646
rect 1914 2573 1933 2576
rect 1954 2603 1973 2606
rect 1914 2556 1917 2573
rect 1906 2553 1917 2556
rect 1906 2436 1909 2553
rect 1914 2516 1917 2536
rect 1922 2523 1925 2536
rect 1930 2523 1941 2526
rect 1914 2513 1921 2516
rect 1918 2456 1921 2513
rect 1918 2453 1925 2456
rect 1930 2453 1933 2523
rect 1946 2513 1949 2536
rect 1898 2433 1909 2436
rect 1922 2436 1925 2453
rect 1922 2433 1933 2436
rect 1898 2413 1901 2433
rect 1906 2413 1917 2416
rect 1882 2273 1893 2276
rect 1874 2213 1877 2246
rect 1882 2203 1885 2273
rect 1890 2203 1893 2216
rect 1866 2193 1885 2196
rect 1866 2143 1869 2186
rect 1882 2143 1885 2193
rect 1898 2156 1901 2406
rect 1906 2386 1909 2406
rect 1914 2403 1925 2406
rect 1906 2383 1925 2386
rect 1906 2226 1909 2376
rect 1922 2373 1925 2383
rect 1930 2366 1933 2433
rect 1938 2393 1941 2506
rect 1914 2363 1933 2366
rect 1914 2263 1917 2363
rect 1922 2343 1925 2356
rect 1922 2303 1925 2336
rect 1930 2316 1933 2336
rect 1938 2323 1941 2346
rect 1930 2313 1941 2316
rect 1946 2313 1949 2416
rect 1954 2323 1957 2603
rect 1962 2533 1973 2536
rect 1970 2503 1973 2526
rect 1978 2496 1981 2636
rect 1986 2603 1989 2643
rect 1994 2586 1997 2666
rect 1986 2523 1989 2586
rect 1994 2583 2005 2586
rect 1994 2533 1997 2546
rect 2002 2526 2005 2536
rect 2010 2533 2013 2673
rect 2018 2526 2021 2546
rect 2034 2536 2037 2926
rect 2042 2816 2045 2936
rect 2050 2826 2053 2926
rect 2058 2883 2061 2936
rect 2082 2933 2085 3063
rect 2090 3013 2093 3066
rect 2138 3046 2141 3133
rect 2146 3116 2149 3213
rect 2154 3193 2157 3206
rect 2162 3133 2165 3246
rect 2178 3193 2181 3336
rect 2186 3203 2189 3473
rect 2194 3306 2197 3476
rect 2206 3436 2209 3503
rect 2206 3433 2213 3436
rect 2202 3393 2205 3416
rect 2202 3323 2205 3356
rect 2210 3336 2213 3433
rect 2218 3346 2221 3556
rect 2226 3533 2229 3576
rect 2234 3533 2237 3556
rect 2250 3546 2253 3753
rect 2258 3653 2261 3766
rect 2290 3746 2293 3766
rect 2286 3743 2293 3746
rect 2274 3713 2277 3726
rect 2258 3613 2261 3636
rect 2250 3543 2257 3546
rect 2226 3473 2229 3526
rect 2226 3423 2237 3426
rect 2242 3423 2245 3536
rect 2254 3456 2257 3543
rect 2266 3533 2269 3696
rect 2274 3573 2277 3656
rect 2286 3646 2289 3743
rect 2298 3703 2301 3716
rect 2306 3696 2309 3813
rect 2298 3693 2309 3696
rect 2286 3643 2293 3646
rect 2282 3603 2285 3626
rect 2274 3536 2277 3556
rect 2282 3543 2285 3596
rect 2274 3533 2285 3536
rect 2274 3513 2277 3526
rect 2282 3473 2285 3533
rect 2290 3513 2293 3643
rect 2298 3506 2301 3693
rect 2306 3613 2309 3626
rect 2314 3603 2317 3826
rect 2346 3753 2349 3886
rect 2354 3803 2357 3826
rect 2322 3743 2349 3746
rect 2362 3743 2365 3923
rect 2370 3893 2373 3926
rect 2370 3763 2373 3886
rect 2378 3843 2381 3966
rect 2430 3956 2433 4023
rect 2430 3953 2437 3956
rect 2378 3793 2381 3806
rect 2322 3726 2325 3736
rect 2322 3723 2341 3726
rect 2338 3613 2341 3626
rect 2346 3616 2349 3743
rect 2354 3623 2357 3736
rect 2362 3683 2365 3726
rect 2378 3703 2381 3716
rect 2346 3613 2357 3616
rect 2362 3613 2365 3626
rect 2306 3583 2309 3596
rect 2314 3533 2317 3546
rect 2314 3516 2317 3526
rect 2290 3503 2301 3506
rect 2306 3513 2317 3516
rect 2322 3513 2325 3556
rect 2250 3453 2257 3456
rect 2226 3353 2229 3416
rect 2250 3406 2253 3453
rect 2246 3403 2253 3406
rect 2218 3343 2229 3346
rect 2210 3333 2221 3336
rect 2194 3303 2201 3306
rect 2210 3303 2213 3326
rect 2198 3196 2201 3303
rect 2194 3193 2201 3196
rect 2146 3113 2157 3116
rect 2114 3043 2141 3046
rect 2154 3046 2157 3113
rect 2154 3043 2165 3046
rect 2114 3026 2117 3043
rect 2110 3023 2117 3026
rect 2122 3033 2157 3036
rect 2066 2893 2069 2926
rect 2090 2916 2093 3006
rect 2082 2913 2093 2916
rect 2082 2846 2085 2913
rect 2082 2843 2089 2846
rect 2098 2843 2101 3016
rect 2110 2966 2113 3023
rect 2122 2983 2125 3033
rect 2130 3013 2157 3016
rect 2138 2976 2141 3006
rect 2122 2973 2141 2976
rect 2110 2963 2117 2966
rect 2114 2943 2117 2963
rect 2106 2913 2109 2936
rect 2122 2933 2125 2973
rect 2050 2823 2077 2826
rect 2042 2813 2053 2816
rect 2058 2813 2077 2816
rect 2002 2523 2021 2526
rect 2026 2533 2037 2536
rect 2026 2516 2029 2533
rect 2010 2513 2029 2516
rect 1962 2493 1981 2496
rect 1962 2413 1965 2493
rect 1938 2306 1941 2313
rect 1938 2303 1949 2306
rect 1962 2266 1965 2406
rect 1970 2373 1973 2446
rect 1978 2413 1989 2416
rect 1978 2403 1989 2406
rect 1978 2333 1981 2366
rect 1994 2333 1997 2506
rect 1970 2283 1973 2316
rect 1954 2263 1965 2266
rect 1906 2223 1941 2226
rect 1906 2166 1909 2206
rect 1914 2203 1917 2216
rect 1922 2213 1933 2216
rect 1922 2203 1925 2213
rect 1930 2176 1933 2206
rect 1938 2183 1941 2223
rect 1946 2213 1949 2226
rect 1954 2206 1957 2263
rect 1946 2203 1957 2206
rect 1946 2176 1949 2203
rect 1930 2173 1949 2176
rect 1906 2163 1941 2166
rect 1898 2153 1917 2156
rect 1866 2123 1869 2136
rect 1874 2116 1877 2136
rect 1870 2113 1877 2116
rect 1870 1966 1873 2113
rect 1882 2093 1885 2126
rect 1890 2053 1893 2146
rect 1898 2046 1901 2146
rect 1914 2076 1917 2153
rect 1938 2123 1941 2163
rect 1946 2106 1949 2173
rect 1890 2043 1901 2046
rect 1906 2073 1917 2076
rect 1942 2103 1949 2106
rect 1890 2013 1893 2043
rect 1898 2006 1901 2036
rect 1882 2003 1901 2006
rect 1866 1963 1873 1966
rect 1866 1906 1869 1963
rect 1882 1933 1885 1976
rect 1906 1973 1909 2073
rect 1906 1923 1909 1956
rect 1866 1903 1885 1906
rect 1866 1866 1869 1896
rect 1882 1886 1885 1903
rect 1882 1883 1901 1886
rect 1866 1863 1877 1866
rect 1874 1816 1877 1863
rect 1890 1833 1893 1856
rect 1866 1813 1877 1816
rect 1866 1793 1869 1813
rect 1858 1783 1877 1786
rect 1834 1753 1861 1756
rect 1826 1743 1837 1746
rect 1834 1723 1837 1743
rect 1858 1733 1861 1753
rect 1874 1733 1877 1783
rect 1794 1506 1797 1526
rect 1794 1503 1801 1506
rect 1798 1426 1801 1503
rect 1794 1423 1801 1426
rect 1794 1396 1797 1423
rect 1810 1413 1813 1606
rect 1818 1516 1821 1546
rect 1826 1533 1829 1566
rect 1834 1533 1837 1616
rect 1842 1613 1845 1726
rect 1850 1653 1853 1716
rect 1858 1603 1861 1726
rect 1866 1713 1885 1716
rect 1866 1696 1869 1713
rect 1866 1693 1873 1696
rect 1870 1606 1873 1693
rect 1866 1603 1873 1606
rect 1866 1586 1869 1603
rect 1858 1583 1869 1586
rect 1818 1513 1829 1516
rect 1826 1436 1829 1513
rect 1858 1446 1861 1583
rect 1882 1546 1885 1706
rect 1890 1613 1893 1806
rect 1898 1796 1901 1883
rect 1906 1803 1909 1916
rect 1898 1793 1909 1796
rect 1906 1723 1909 1793
rect 1914 1716 1917 2066
rect 1922 2013 1925 2046
rect 1942 2036 1945 2103
rect 1942 2033 1949 2036
rect 1930 2013 1941 2016
rect 1922 2003 1933 2006
rect 1922 1893 1925 2003
rect 1938 1966 1941 2013
rect 1946 2003 1949 2033
rect 1930 1963 1941 1966
rect 1930 1923 1933 1963
rect 1954 1923 1957 2186
rect 1922 1813 1925 1836
rect 1938 1823 1949 1826
rect 1930 1813 1941 1816
rect 1938 1783 1941 1813
rect 1946 1736 1949 1816
rect 1954 1803 1957 1836
rect 1922 1733 1933 1736
rect 1906 1713 1917 1716
rect 1922 1713 1925 1726
rect 1906 1646 1909 1713
rect 1898 1643 1909 1646
rect 1898 1603 1901 1643
rect 1906 1613 1909 1626
rect 1874 1543 1885 1546
rect 1914 1546 1917 1606
rect 1922 1583 1925 1616
rect 1914 1543 1925 1546
rect 1874 1523 1877 1543
rect 1858 1443 1869 1446
rect 1818 1433 1829 1436
rect 1802 1403 1813 1406
rect 1778 1393 1785 1396
rect 1794 1393 1805 1396
rect 1754 1383 1773 1386
rect 1738 1313 1749 1316
rect 1706 1273 1717 1276
rect 1706 1156 1709 1273
rect 1730 1196 1733 1246
rect 1698 1153 1709 1156
rect 1722 1193 1733 1196
rect 1674 1123 1685 1126
rect 1674 1056 1677 1123
rect 1690 1106 1693 1136
rect 1666 1053 1677 1056
rect 1686 1103 1693 1106
rect 1658 996 1661 1016
rect 1666 1006 1669 1053
rect 1686 1036 1689 1103
rect 1698 1043 1701 1153
rect 1706 1123 1709 1146
rect 1674 1023 1677 1036
rect 1686 1033 1693 1036
rect 1674 1013 1685 1016
rect 1666 1003 1685 1006
rect 1658 993 1669 996
rect 1650 973 1657 976
rect 1654 866 1657 973
rect 1666 923 1669 993
rect 1674 933 1677 956
rect 1682 933 1685 1003
rect 1654 863 1669 866
rect 1642 853 1661 856
rect 1666 846 1669 863
rect 1658 843 1669 846
rect 1690 846 1693 1033
rect 1698 913 1701 1006
rect 1706 996 1709 1036
rect 1714 1003 1717 1126
rect 1722 1123 1725 1193
rect 1730 1133 1733 1146
rect 1738 1123 1741 1216
rect 1746 1166 1749 1313
rect 1754 1286 1757 1383
rect 1762 1323 1765 1336
rect 1782 1316 1785 1393
rect 1778 1313 1785 1316
rect 1754 1283 1773 1286
rect 1754 1183 1757 1216
rect 1770 1176 1773 1283
rect 1762 1173 1773 1176
rect 1746 1163 1757 1166
rect 1746 1133 1749 1156
rect 1754 1123 1757 1163
rect 1722 1013 1725 1096
rect 1762 1073 1765 1173
rect 1746 1013 1749 1036
rect 1706 993 1717 996
rect 1706 873 1709 946
rect 1714 853 1717 993
rect 1730 936 1733 1006
rect 1754 996 1757 1046
rect 1762 1013 1765 1036
rect 1722 933 1733 936
rect 1746 993 1757 996
rect 1722 896 1725 933
rect 1730 903 1733 926
rect 1722 893 1741 896
rect 1690 843 1725 846
rect 1650 816 1653 826
rect 1642 813 1653 816
rect 1642 796 1645 813
rect 1610 623 1629 626
rect 1634 793 1645 796
rect 1610 533 1613 623
rect 1618 613 1629 616
rect 1634 613 1637 793
rect 1618 533 1621 556
rect 1610 513 1613 526
rect 1626 483 1629 606
rect 1642 553 1645 746
rect 1658 733 1661 843
rect 1674 803 1677 836
rect 1674 733 1677 786
rect 1682 743 1701 746
rect 1714 743 1717 816
rect 1650 623 1653 676
rect 1650 583 1653 616
rect 1658 596 1661 606
rect 1666 603 1669 636
rect 1682 613 1685 743
rect 1690 716 1693 726
rect 1698 723 1701 743
rect 1690 713 1701 716
rect 1698 603 1701 713
rect 1706 703 1709 736
rect 1722 726 1725 843
rect 1738 826 1741 893
rect 1746 833 1749 993
rect 1762 943 1765 1006
rect 1770 986 1773 1146
rect 1778 1013 1781 1313
rect 1794 1296 1797 1326
rect 1786 1293 1797 1296
rect 1802 1293 1805 1393
rect 1786 1096 1789 1236
rect 1794 1153 1797 1206
rect 1802 1116 1805 1216
rect 1810 1153 1813 1396
rect 1818 1226 1821 1433
rect 1866 1426 1869 1443
rect 1826 1373 1829 1406
rect 1826 1273 1829 1366
rect 1818 1223 1829 1226
rect 1818 1193 1821 1216
rect 1818 1153 1821 1186
rect 1826 1176 1829 1223
rect 1834 1213 1837 1416
rect 1850 1413 1853 1426
rect 1866 1423 1873 1426
rect 1842 1333 1845 1406
rect 1850 1363 1853 1406
rect 1858 1393 1861 1406
rect 1870 1366 1873 1423
rect 1882 1376 1885 1536
rect 1890 1533 1917 1536
rect 1890 1523 1893 1533
rect 1898 1523 1917 1526
rect 1898 1433 1901 1523
rect 1914 1483 1917 1516
rect 1922 1463 1925 1543
rect 1930 1506 1933 1733
rect 1938 1523 1941 1736
rect 1946 1733 1957 1736
rect 1946 1706 1949 1726
rect 1954 1723 1957 1733
rect 1946 1703 1953 1706
rect 1950 1636 1953 1703
rect 1946 1633 1953 1636
rect 1946 1523 1949 1633
rect 1954 1563 1957 1616
rect 1962 1556 1965 2256
rect 1970 2203 1973 2216
rect 1978 2083 1981 2326
rect 1986 2203 1989 2216
rect 1994 2203 1997 2216
rect 2002 2183 2005 2436
rect 2010 2403 2013 2513
rect 2010 2333 2013 2356
rect 2018 2323 2021 2506
rect 2034 2503 2037 2526
rect 2042 2476 2045 2806
rect 2050 2766 2053 2813
rect 2074 2773 2077 2806
rect 2050 2763 2061 2766
rect 2058 2663 2061 2763
rect 2086 2756 2089 2843
rect 2106 2816 2109 2866
rect 2114 2826 2117 2926
rect 2130 2836 2133 2936
rect 2138 2923 2141 2946
rect 2146 2843 2149 3006
rect 2130 2833 2141 2836
rect 2114 2823 2125 2826
rect 2106 2813 2125 2816
rect 2098 2786 2101 2806
rect 2098 2783 2117 2786
rect 2066 2656 2069 2756
rect 2082 2753 2089 2756
rect 2074 2696 2077 2726
rect 2082 2703 2085 2753
rect 2098 2733 2101 2776
rect 2114 2753 2117 2783
rect 2098 2696 2101 2726
rect 2122 2723 2125 2806
rect 2130 2773 2133 2816
rect 2138 2756 2141 2833
rect 2154 2826 2157 3013
rect 2162 2943 2165 3043
rect 2170 3023 2173 3146
rect 2186 3036 2189 3126
rect 2194 3053 2197 3193
rect 2202 3123 2205 3136
rect 2210 3126 2213 3246
rect 2218 3133 2221 3333
rect 2226 3193 2229 3343
rect 2234 3263 2237 3326
rect 2246 3296 2249 3403
rect 2258 3303 2261 3436
rect 2266 3393 2269 3426
rect 2274 3353 2277 3416
rect 2246 3293 2253 3296
rect 2250 3236 2253 3293
rect 2266 3246 2269 3316
rect 2274 3253 2277 3316
rect 2282 3263 2285 3326
rect 2290 3246 2293 3503
rect 2298 3413 2301 3436
rect 2306 3423 2309 3513
rect 2330 3506 2333 3536
rect 2314 3503 2333 3506
rect 2346 3526 2349 3606
rect 2354 3533 2357 3613
rect 2346 3523 2357 3526
rect 2314 3403 2317 3503
rect 2266 3243 2277 3246
rect 2250 3233 2269 3236
rect 2234 3213 2253 3216
rect 2258 3213 2261 3226
rect 2234 3203 2237 3213
rect 2266 3206 2269 3233
rect 2258 3203 2269 3206
rect 2226 3126 2229 3136
rect 2234 3133 2237 3196
rect 2274 3193 2277 3243
rect 2282 3243 2293 3246
rect 2282 3203 2285 3243
rect 2290 3186 2293 3236
rect 2266 3183 2293 3186
rect 2210 3123 2229 3126
rect 2186 3033 2205 3036
rect 2170 2983 2173 3006
rect 2178 2936 2181 3016
rect 2186 3013 2197 3016
rect 2202 3006 2205 3033
rect 2170 2933 2181 2936
rect 2186 3003 2205 3006
rect 2186 2933 2189 3003
rect 2162 2836 2165 2916
rect 2170 2883 2173 2933
rect 2178 2843 2181 2926
rect 2194 2923 2197 2956
rect 2202 2863 2205 2996
rect 2210 2976 2213 3036
rect 2234 3016 2237 3126
rect 2266 3123 2269 3183
rect 2298 3166 2301 3316
rect 2306 3303 2309 3326
rect 2314 3313 2317 3396
rect 2322 3353 2325 3416
rect 2314 3223 2317 3276
rect 2330 3243 2333 3436
rect 2338 3403 2341 3496
rect 2346 3366 2349 3523
rect 2362 3473 2365 3596
rect 2370 3586 2373 3606
rect 2386 3603 2389 3936
rect 2394 3933 2397 3946
rect 2410 3926 2413 3936
rect 2418 3933 2429 3936
rect 2402 3893 2405 3926
rect 2410 3923 2421 3926
rect 2426 3863 2429 3896
rect 2394 3673 2397 3826
rect 2402 3823 2429 3826
rect 2402 3793 2405 3823
rect 2410 3793 2413 3806
rect 2418 3746 2421 3816
rect 2402 3743 2421 3746
rect 2402 3733 2405 3743
rect 2402 3713 2405 3726
rect 2410 3663 2413 3736
rect 2418 3633 2421 3726
rect 2426 3716 2429 3823
rect 2434 3803 2437 3953
rect 2442 3896 2445 4033
rect 2458 4003 2461 4066
rect 2482 4013 2485 4046
rect 2490 3976 2493 4036
rect 2458 3973 2493 3976
rect 2458 3933 2461 3973
rect 2498 3953 2501 4086
rect 2482 3923 2485 3946
rect 2442 3893 2449 3896
rect 2446 3836 2449 3893
rect 2498 3886 2501 3936
rect 2466 3883 2501 3886
rect 2442 3833 2449 3836
rect 2434 3726 2437 3796
rect 2442 3793 2445 3833
rect 2450 3733 2453 3816
rect 2458 3793 2461 3866
rect 2466 3803 2469 3883
rect 2506 3863 2509 4113
rect 2538 4106 2541 4143
rect 2554 4133 2557 4196
rect 2562 4166 2565 4337
rect 2578 4213 2581 4236
rect 2586 4213 2589 4276
rect 2610 4266 2613 4340
rect 2722 4296 2725 4340
rect 2674 4293 2725 4296
rect 2610 4263 2621 4266
rect 2610 4216 2613 4226
rect 2594 4213 2613 4216
rect 2594 4173 2597 4213
rect 2602 4203 2613 4206
rect 2602 4166 2605 4196
rect 2562 4163 2581 4166
rect 2522 4103 2541 4106
rect 2522 3973 2525 4103
rect 2522 3886 2525 3946
rect 2530 3933 2533 4086
rect 2514 3883 2525 3886
rect 2474 3753 2477 3816
rect 2482 3806 2485 3856
rect 2490 3823 2509 3826
rect 2490 3813 2493 3823
rect 2482 3803 2493 3806
rect 2498 3773 2501 3816
rect 2514 3806 2517 3883
rect 2522 3813 2525 3866
rect 2530 3823 2533 3846
rect 2514 3803 2525 3806
rect 2434 3723 2445 3726
rect 2426 3713 2437 3716
rect 2394 3586 2397 3616
rect 2370 3583 2397 3586
rect 2402 3576 2405 3616
rect 2370 3573 2405 3576
rect 2370 3533 2373 3573
rect 2378 3546 2381 3566
rect 2378 3543 2385 3546
rect 2370 3493 2373 3516
rect 2382 3476 2385 3543
rect 2394 3533 2405 3536
rect 2394 3523 2405 3526
rect 2410 3496 2413 3616
rect 2434 3603 2437 3713
rect 2442 3693 2445 3723
rect 2450 3703 2453 3716
rect 2458 3663 2461 3736
rect 2466 3726 2469 3746
rect 2466 3723 2477 3726
rect 2498 3723 2501 3746
rect 2506 3726 2509 3736
rect 2514 3733 2517 3796
rect 2530 3773 2533 3816
rect 2538 3733 2541 4036
rect 2546 4013 2549 4096
rect 2554 4033 2557 4116
rect 2546 3923 2549 3976
rect 2554 3943 2557 4016
rect 2562 4003 2565 4046
rect 2562 3936 2565 3996
rect 2570 3976 2573 4016
rect 2578 3993 2581 4163
rect 2594 4163 2605 4166
rect 2586 4003 2589 4106
rect 2594 4083 2597 4163
rect 2618 4146 2621 4263
rect 2634 4213 2637 4236
rect 2650 4203 2653 4216
rect 2658 4196 2661 4276
rect 2666 4223 2669 4266
rect 2666 4203 2669 4216
rect 2642 4193 2661 4196
rect 2642 4183 2645 4193
rect 2674 4186 2677 4293
rect 2682 4213 2685 4276
rect 2690 4203 2693 4286
rect 2618 4143 2637 4146
rect 2570 3973 2581 3976
rect 2554 3933 2565 3936
rect 2578 3933 2581 3973
rect 2594 3946 2597 4016
rect 2602 4003 2605 4126
rect 2618 4043 2621 4143
rect 2634 4123 2637 4143
rect 2642 4123 2645 4136
rect 2658 4133 2661 4186
rect 2666 4183 2677 4186
rect 2666 4143 2669 4183
rect 2698 4163 2701 4216
rect 2674 4153 2701 4156
rect 2674 4133 2677 4153
rect 2682 4133 2685 4146
rect 2594 3943 2605 3946
rect 2610 3943 2613 4016
rect 2634 3993 2637 4006
rect 2546 3806 2549 3896
rect 2554 3813 2557 3846
rect 2546 3803 2557 3806
rect 2562 3803 2565 3926
rect 2602 3836 2605 3943
rect 2626 3923 2629 3946
rect 2598 3833 2605 3836
rect 2506 3723 2525 3726
rect 2466 3646 2469 3716
rect 2482 3713 2493 3716
rect 2482 3666 2485 3713
rect 2474 3663 2485 3666
rect 2474 3653 2477 3663
rect 2482 3653 2493 3656
rect 2482 3646 2485 3653
rect 2498 3646 2501 3666
rect 2466 3643 2485 3646
rect 2490 3643 2501 3646
rect 2450 3616 2453 3626
rect 2442 3603 2445 3616
rect 2450 3613 2477 3616
rect 2402 3493 2413 3496
rect 2382 3473 2389 3476
rect 2354 3413 2357 3426
rect 2354 3393 2357 3406
rect 2338 3323 2341 3366
rect 2346 3363 2357 3366
rect 2362 3336 2365 3456
rect 2378 3423 2381 3456
rect 2386 3403 2389 3473
rect 2394 3396 2397 3406
rect 2346 3333 2365 3336
rect 2378 3393 2397 3396
rect 2346 3306 2349 3333
rect 2342 3303 2349 3306
rect 2354 3323 2365 3326
rect 2322 3213 2325 3236
rect 2282 3163 2301 3166
rect 2250 3053 2253 3116
rect 2258 3083 2269 3086
rect 2274 3083 2277 3136
rect 2282 3123 2285 3163
rect 2290 3133 2301 3136
rect 2306 3123 2309 3196
rect 2314 3153 2325 3156
rect 2330 3153 2333 3236
rect 2342 3226 2345 3303
rect 2342 3223 2349 3226
rect 2314 3083 2317 3136
rect 2322 3126 2325 3153
rect 2346 3136 2349 3223
rect 2354 3146 2357 3323
rect 2362 3303 2365 3323
rect 2378 3313 2381 3393
rect 2394 3346 2397 3366
rect 2390 3343 2397 3346
rect 2378 3286 2381 3306
rect 2370 3283 2381 3286
rect 2362 3203 2365 3266
rect 2370 3213 2373 3283
rect 2390 3226 2393 3343
rect 2402 3263 2405 3493
rect 2418 3486 2421 3536
rect 2426 3523 2429 3546
rect 2434 3523 2437 3536
rect 2442 3523 2445 3536
rect 2450 3493 2453 3526
rect 2410 3483 2421 3486
rect 2458 3483 2461 3536
rect 2466 3486 2469 3606
rect 2482 3563 2485 3606
rect 2490 3543 2493 3643
rect 2498 3603 2501 3636
rect 2506 3556 2509 3616
rect 2498 3553 2509 3556
rect 2466 3483 2477 3486
rect 2482 3483 2485 3526
rect 2410 3386 2413 3483
rect 2418 3403 2421 3476
rect 2450 3423 2453 3476
rect 2474 3466 2477 3483
rect 2458 3463 2477 3466
rect 2458 3416 2461 3463
rect 2474 3423 2485 3426
rect 2410 3383 2421 3386
rect 2410 3333 2413 3376
rect 2418 3256 2421 3383
rect 2426 3373 2429 3416
rect 2426 3353 2429 3366
rect 2426 3313 2429 3336
rect 2434 3263 2437 3406
rect 2442 3353 2445 3416
rect 2458 3413 2477 3416
rect 2450 3403 2461 3406
rect 2458 3333 2469 3336
rect 2450 3323 2461 3326
rect 2418 3253 2429 3256
rect 2390 3223 2397 3226
rect 2378 3203 2389 3206
rect 2354 3143 2381 3146
rect 2338 3133 2349 3136
rect 2362 3126 2365 3136
rect 2322 3123 2365 3126
rect 2242 3023 2245 3046
rect 2250 3043 2261 3046
rect 2226 3013 2237 3016
rect 2250 3003 2253 3043
rect 2266 3003 2269 3083
rect 2330 3063 2333 3116
rect 2362 3083 2365 3116
rect 2370 3093 2373 3126
rect 2282 3043 2293 3046
rect 2290 3013 2293 3043
rect 2210 2973 2237 2976
rect 2226 2893 2229 2936
rect 2162 2833 2181 2836
rect 2154 2823 2173 2826
rect 2134 2753 2141 2756
rect 2074 2693 2101 2696
rect 2066 2653 2077 2656
rect 2074 2636 2077 2653
rect 2074 2633 2081 2636
rect 2050 2563 2053 2616
rect 2050 2486 2053 2536
rect 2058 2513 2061 2626
rect 2078 2576 2081 2633
rect 2074 2573 2081 2576
rect 2066 2496 2069 2536
rect 2074 2533 2077 2573
rect 2082 2503 2085 2546
rect 2090 2543 2093 2616
rect 2098 2563 2101 2693
rect 2134 2686 2137 2753
rect 2134 2683 2141 2686
rect 2130 2636 2133 2666
rect 2114 2633 2133 2636
rect 2138 2633 2141 2683
rect 2146 2663 2149 2806
rect 2170 2803 2173 2816
rect 2178 2796 2181 2833
rect 2170 2793 2181 2796
rect 2066 2493 2077 2496
rect 2050 2483 2069 2486
rect 2034 2466 2037 2476
rect 2042 2473 2053 2476
rect 2034 2463 2061 2466
rect 2026 2346 2029 2416
rect 2034 2413 2045 2416
rect 2042 2373 2045 2406
rect 2050 2356 2053 2416
rect 2058 2403 2061 2463
rect 2042 2353 2053 2356
rect 2026 2343 2037 2346
rect 2026 2303 2029 2336
rect 2034 2276 2037 2343
rect 2018 2273 2037 2276
rect 2002 2133 2005 2146
rect 1986 2123 1997 2126
rect 2002 2083 2005 2126
rect 2010 2063 2013 2266
rect 2018 2203 2021 2273
rect 2010 2013 2013 2026
rect 1978 1973 1981 2006
rect 1970 1913 1973 1956
rect 1978 1896 1981 1946
rect 1994 1933 1997 1956
rect 2010 1933 2013 1946
rect 1986 1913 1989 1926
rect 1994 1906 1997 1926
rect 2002 1923 2013 1926
rect 1994 1903 2001 1906
rect 1974 1893 1981 1896
rect 1974 1816 1977 1893
rect 1970 1813 1977 1816
rect 1970 1796 1973 1813
rect 1986 1803 1989 1866
rect 1998 1826 2001 1903
rect 1994 1823 2001 1826
rect 1970 1793 1981 1796
rect 1970 1733 1973 1746
rect 1978 1713 1981 1793
rect 1986 1613 1989 1746
rect 1994 1716 1997 1823
rect 2002 1763 2005 1806
rect 2002 1723 2005 1736
rect 2010 1733 2013 1896
rect 1994 1713 2001 1716
rect 1978 1593 1981 1606
rect 1954 1553 1965 1556
rect 1954 1526 1957 1553
rect 1970 1536 1973 1576
rect 1962 1533 1973 1536
rect 1978 1526 1981 1586
rect 1998 1556 2001 1713
rect 2010 1613 2013 1726
rect 2010 1583 2013 1606
rect 2018 1593 2021 2196
rect 2034 2193 2037 2273
rect 2042 2243 2045 2353
rect 2050 2273 2053 2346
rect 2058 2333 2061 2356
rect 2066 2266 2069 2483
rect 2074 2393 2077 2493
rect 2074 2323 2077 2386
rect 2050 2263 2069 2266
rect 2026 2123 2029 2186
rect 2050 2146 2053 2263
rect 2074 2213 2077 2226
rect 2034 2133 2037 2146
rect 2042 2143 2053 2146
rect 2026 1983 2029 2066
rect 2042 2023 2045 2143
rect 2050 2016 2053 2136
rect 2066 2133 2069 2196
rect 2074 2126 2077 2206
rect 2058 2123 2077 2126
rect 2058 2113 2061 2123
rect 2082 2036 2085 2406
rect 2090 2343 2093 2476
rect 2098 2353 2101 2526
rect 2106 2473 2109 2616
rect 2090 2316 2093 2336
rect 2106 2323 2109 2366
rect 2090 2313 2097 2316
rect 2094 2246 2097 2313
rect 2106 2293 2109 2316
rect 2090 2243 2097 2246
rect 2090 2223 2093 2243
rect 2090 2113 2093 2176
rect 2098 2113 2101 2126
rect 2106 2093 2109 2106
rect 2042 2013 2053 2016
rect 2058 2013 2061 2036
rect 2066 2033 2085 2036
rect 2042 1943 2045 2013
rect 2066 1953 2069 2033
rect 2082 1983 2085 2026
rect 2106 2013 2109 2056
rect 2026 1913 2029 1936
rect 2106 1933 2109 1976
rect 2114 1933 2117 2633
rect 2130 2626 2133 2633
rect 2130 2623 2149 2626
rect 2146 2613 2149 2623
rect 2122 2373 2125 2416
rect 2130 2366 2133 2416
rect 2138 2403 2141 2456
rect 2138 2373 2141 2396
rect 2146 2386 2149 2526
rect 2162 2516 2165 2756
rect 2170 2523 2173 2793
rect 2194 2773 2197 2806
rect 2218 2756 2221 2876
rect 2234 2836 2237 2973
rect 2250 2946 2253 2996
rect 2250 2943 2261 2946
rect 2250 2926 2253 2936
rect 2242 2923 2253 2926
rect 2242 2913 2245 2923
rect 2250 2883 2253 2916
rect 2234 2833 2241 2836
rect 2226 2813 2229 2826
rect 2238 2776 2241 2833
rect 2258 2823 2261 2943
rect 2266 2896 2269 2996
rect 2298 2993 2301 3056
rect 2378 3053 2381 3143
rect 2306 2986 2309 3016
rect 2282 2983 2309 2986
rect 2266 2893 2273 2896
rect 2270 2836 2273 2893
rect 2282 2876 2285 2983
rect 2346 2966 2349 3016
rect 2346 2963 2353 2966
rect 2306 2913 2309 2926
rect 2322 2876 2325 2896
rect 2350 2886 2353 2963
rect 2362 2936 2365 3026
rect 2370 3013 2373 3026
rect 2378 2996 2381 3036
rect 2386 3006 2389 3026
rect 2394 3013 2397 3223
rect 2402 3216 2405 3246
rect 2410 3223 2421 3226
rect 2402 3213 2413 3216
rect 2410 3123 2413 3213
rect 2418 3133 2421 3206
rect 2426 3203 2429 3253
rect 2434 3213 2437 3226
rect 2442 3203 2445 3256
rect 2450 3146 2453 3226
rect 2458 3203 2461 3266
rect 2466 3213 2469 3316
rect 2474 3223 2477 3413
rect 2482 3403 2485 3416
rect 2490 3356 2493 3536
rect 2498 3513 2501 3553
rect 2506 3523 2509 3546
rect 2498 3413 2501 3426
rect 2482 3353 2493 3356
rect 2482 3296 2485 3353
rect 2498 3323 2501 3336
rect 2506 3323 2509 3506
rect 2514 3416 2517 3566
rect 2530 3543 2533 3626
rect 2538 3613 2541 3696
rect 2546 3616 2549 3726
rect 2554 3656 2557 3803
rect 2570 3783 2573 3806
rect 2570 3726 2573 3766
rect 2578 3733 2581 3796
rect 2586 3753 2589 3816
rect 2598 3736 2601 3833
rect 2610 3823 2637 3826
rect 2610 3793 2613 3816
rect 2618 3783 2621 3816
rect 2634 3813 2637 3823
rect 2594 3733 2601 3736
rect 2610 3733 2613 3776
rect 2562 3663 2565 3726
rect 2570 3723 2577 3726
rect 2554 3653 2565 3656
rect 2546 3613 2557 3616
rect 2562 3606 2565 3653
rect 2574 3646 2577 3723
rect 2586 3673 2589 3726
rect 2594 3703 2597 3733
rect 2574 3643 2581 3646
rect 2578 3623 2581 3643
rect 2546 3603 2565 3606
rect 2570 3613 2581 3616
rect 2570 3576 2573 3613
rect 2586 3603 2589 3636
rect 2538 3573 2573 3576
rect 2530 3516 2533 3536
rect 2538 3523 2541 3573
rect 2594 3563 2597 3616
rect 2602 3556 2605 3726
rect 2610 3613 2613 3726
rect 2618 3606 2621 3766
rect 2626 3753 2629 3806
rect 2626 3673 2629 3726
rect 2546 3523 2549 3546
rect 2562 3523 2565 3556
rect 2594 3553 2605 3556
rect 2610 3603 2621 3606
rect 2570 3516 2573 3536
rect 2530 3513 2541 3516
rect 2522 3423 2525 3506
rect 2530 3483 2533 3506
rect 2514 3413 2525 3416
rect 2514 3316 2517 3326
rect 2490 3313 2517 3316
rect 2482 3293 2493 3296
rect 2490 3236 2493 3293
rect 2522 3253 2525 3413
rect 2530 3403 2533 3426
rect 2538 3336 2541 3513
rect 2554 3513 2573 3516
rect 2546 3413 2549 3476
rect 2554 3406 2557 3513
rect 2562 3486 2565 3506
rect 2578 3503 2581 3526
rect 2586 3493 2589 3536
rect 2594 3486 2597 3553
rect 2602 3523 2605 3546
rect 2562 3483 2597 3486
rect 2562 3413 2565 3483
rect 2570 3406 2573 3476
rect 2610 3473 2613 3603
rect 2618 3523 2621 3596
rect 2626 3576 2629 3666
rect 2634 3653 2637 3726
rect 2642 3646 2645 4086
rect 2650 3896 2653 4126
rect 2666 4123 2685 4126
rect 2658 4003 2661 4106
rect 2682 4056 2685 4123
rect 2690 4116 2693 4136
rect 2698 4123 2701 4153
rect 2706 4146 2709 4286
rect 2722 4213 2725 4293
rect 2746 4283 2749 4340
rect 2722 4176 2725 4206
rect 2754 4183 2757 4216
rect 2762 4176 2765 4316
rect 2786 4196 2789 4326
rect 2826 4306 2829 4340
rect 2802 4303 2829 4306
rect 2802 4236 2805 4303
rect 2802 4233 2813 4236
rect 2794 4213 2805 4216
rect 2786 4193 2793 4196
rect 2770 4176 2773 4186
rect 2722 4173 2773 4176
rect 2706 4143 2717 4146
rect 2690 4113 2701 4116
rect 2706 4113 2709 4136
rect 2682 4053 2693 4056
rect 2666 4013 2669 4036
rect 2682 3993 2685 4016
rect 2690 4003 2693 4053
rect 2698 4013 2701 4113
rect 2658 3923 2661 3936
rect 2666 3906 2669 3956
rect 2682 3953 2701 3956
rect 2706 3953 2709 4016
rect 2714 4003 2717 4143
rect 2722 4143 2749 4146
rect 2722 4106 2725 4143
rect 2730 4133 2741 4136
rect 2730 4123 2733 4133
rect 2722 4103 2729 4106
rect 2726 4006 2729 4103
rect 2738 4096 2741 4126
rect 2746 4123 2749 4143
rect 2754 4113 2757 4136
rect 2762 4103 2765 4126
rect 2770 4096 2773 4136
rect 2778 4133 2781 4146
rect 2778 4103 2781 4126
rect 2790 4096 2793 4193
rect 2810 4143 2813 4233
rect 2818 4213 2821 4296
rect 2834 4253 2837 4276
rect 2818 4203 2829 4206
rect 2834 4163 2837 4216
rect 2738 4093 2773 4096
rect 2786 4093 2793 4096
rect 2726 4003 2733 4006
rect 2746 4003 2749 4066
rect 2674 3923 2677 3936
rect 2682 3923 2685 3953
rect 2698 3946 2701 3953
rect 2690 3933 2693 3946
rect 2698 3943 2717 3946
rect 2706 3926 2709 3936
rect 2714 3933 2717 3943
rect 2722 3936 2725 3996
rect 2730 3943 2733 4003
rect 2722 3933 2733 3936
rect 2698 3916 2701 3926
rect 2706 3923 2717 3926
rect 2698 3913 2709 3916
rect 2666 3903 2701 3906
rect 2650 3893 2677 3896
rect 2650 3773 2653 3816
rect 2658 3813 2661 3866
rect 2666 3856 2669 3886
rect 2674 3866 2677 3893
rect 2674 3863 2685 3866
rect 2666 3853 2677 3856
rect 2658 3783 2661 3806
rect 2666 3803 2669 3846
rect 2674 3786 2677 3853
rect 2682 3806 2685 3863
rect 2690 3813 2693 3866
rect 2682 3803 2693 3806
rect 2674 3783 2681 3786
rect 2634 3643 2645 3646
rect 2634 3603 2637 3643
rect 2650 3636 2653 3736
rect 2658 3713 2661 3766
rect 2666 3723 2669 3776
rect 2678 3726 2681 3783
rect 2690 3733 2693 3803
rect 2698 3756 2701 3903
rect 2706 3863 2709 3913
rect 2730 3843 2733 3926
rect 2746 3906 2749 3946
rect 2754 3913 2757 3936
rect 2762 3923 2765 3996
rect 2770 3973 2773 4016
rect 2786 3983 2789 4093
rect 2810 4063 2813 4136
rect 2834 4113 2837 4126
rect 2826 4013 2829 4046
rect 2842 3996 2845 4340
rect 2922 4326 2925 4340
rect 2918 4323 2925 4326
rect 2850 4203 2853 4256
rect 2858 4196 2861 4216
rect 2866 4203 2869 4306
rect 2874 4213 2877 4276
rect 2890 4213 2893 4276
rect 2906 4223 2909 4316
rect 2918 4236 2921 4323
rect 2918 4233 2925 4236
rect 2922 4216 2925 4233
rect 2898 4213 2909 4216
rect 2914 4213 2925 4216
rect 2930 4213 2933 4326
rect 2898 4206 2901 4213
rect 2882 4203 2901 4206
rect 2906 4196 2909 4206
rect 2850 4063 2853 4196
rect 2858 4193 2909 4196
rect 2914 4193 2917 4213
rect 2858 4086 2861 4186
rect 2890 4123 2893 4146
rect 2906 4133 2909 4186
rect 2922 4146 2925 4213
rect 2938 4176 2941 4340
rect 2954 4306 2957 4326
rect 2954 4303 2965 4306
rect 2946 4193 2949 4266
rect 2962 4246 2965 4303
rect 2994 4263 2997 4340
rect 3002 4286 3005 4306
rect 3002 4283 3013 4286
rect 2954 4243 2965 4246
rect 2954 4213 2957 4243
rect 2962 4223 2989 4226
rect 2938 4173 2945 4176
rect 2962 4173 2965 4223
rect 2970 4213 2981 4216
rect 2994 4213 2997 4256
rect 3010 4236 3013 4283
rect 3002 4233 3013 4236
rect 3002 4213 3005 4233
rect 2922 4143 2933 4146
rect 2858 4083 2869 4086
rect 2866 4003 2869 4083
rect 2810 3993 2845 3996
rect 2746 3903 2757 3906
rect 2706 3766 2709 3836
rect 2714 3813 2717 3826
rect 2722 3823 2733 3826
rect 2738 3803 2741 3866
rect 2746 3793 2749 3816
rect 2706 3763 2733 3766
rect 2698 3753 2709 3756
rect 2674 3723 2681 3726
rect 2642 3633 2653 3636
rect 2642 3613 2645 3633
rect 2650 3613 2661 3616
rect 2626 3573 2645 3576
rect 2530 3333 2541 3336
rect 2546 3403 2557 3406
rect 2562 3403 2573 3406
rect 2578 3403 2581 3466
rect 2586 3463 2621 3466
rect 2626 3463 2629 3556
rect 2634 3533 2637 3566
rect 2642 3553 2645 3573
rect 2650 3546 2653 3613
rect 2666 3606 2669 3666
rect 2642 3543 2653 3546
rect 2658 3603 2669 3606
rect 2642 3526 2645 3543
rect 2634 3523 2645 3526
rect 2634 3506 2637 3523
rect 2634 3503 2645 3506
rect 2650 3503 2653 3536
rect 2530 3246 2533 3333
rect 2486 3233 2493 3236
rect 2514 3243 2533 3246
rect 2450 3143 2461 3146
rect 2426 3123 2429 3136
rect 2434 3093 2437 3136
rect 2442 3063 2445 3126
rect 2458 3043 2461 3143
rect 2466 3063 2469 3206
rect 2474 3193 2477 3216
rect 2486 3186 2489 3233
rect 2482 3183 2489 3186
rect 2498 3213 2509 3216
rect 2474 3106 2477 3136
rect 2482 3123 2485 3183
rect 2498 3123 2501 3213
rect 2506 3183 2509 3206
rect 2474 3103 2485 3106
rect 2482 3046 2485 3103
rect 2514 3093 2517 3243
rect 2522 3133 2525 3226
rect 2530 3203 2533 3226
rect 2538 3223 2541 3326
rect 2546 3296 2549 3403
rect 2562 3396 2565 3403
rect 2554 3393 2565 3396
rect 2554 3316 2557 3393
rect 2562 3323 2565 3336
rect 2570 3333 2573 3396
rect 2578 3323 2581 3366
rect 2586 3333 2589 3463
rect 2602 3413 2605 3456
rect 2618 3413 2621 3463
rect 2594 3363 2597 3406
rect 2602 3333 2605 3406
rect 2610 3343 2613 3406
rect 2618 3363 2621 3406
rect 2626 3383 2629 3456
rect 2634 3413 2637 3496
rect 2642 3473 2645 3503
rect 2642 3406 2645 3426
rect 2634 3403 2645 3406
rect 2634 3336 2637 3403
rect 2650 3396 2653 3416
rect 2642 3393 2653 3396
rect 2642 3373 2645 3393
rect 2658 3386 2661 3603
rect 2666 3563 2669 3596
rect 2666 3413 2669 3466
rect 2610 3333 2637 3336
rect 2586 3316 2589 3326
rect 2594 3316 2597 3326
rect 2554 3313 2597 3316
rect 2610 3306 2613 3333
rect 2546 3293 2553 3296
rect 2550 3236 2553 3293
rect 2546 3233 2553 3236
rect 2538 3183 2541 3216
rect 2546 3176 2549 3233
rect 2554 3203 2557 3216
rect 2562 3203 2565 3256
rect 2578 3223 2581 3306
rect 2586 3303 2613 3306
rect 2586 3216 2589 3303
rect 2530 3173 2549 3176
rect 2522 3083 2525 3126
rect 2530 3063 2533 3173
rect 2570 3146 2573 3216
rect 2582 3213 2589 3216
rect 2582 3156 2585 3213
rect 2562 3143 2573 3146
rect 2578 3153 2585 3156
rect 2562 3133 2565 3143
rect 2570 3076 2573 3136
rect 2578 3123 2581 3153
rect 2586 3083 2589 3136
rect 2594 3123 2597 3256
rect 2618 3223 2621 3326
rect 2602 3196 2605 3206
rect 2626 3203 2629 3286
rect 2634 3196 2637 3246
rect 2602 3193 2637 3196
rect 2602 3133 2637 3136
rect 2602 3113 2605 3133
rect 2570 3073 2597 3076
rect 2482 3043 2501 3046
rect 2386 3003 2397 3006
rect 2402 3003 2413 3006
rect 2402 2996 2405 3003
rect 2378 2993 2405 2996
rect 2410 2963 2413 2996
rect 2418 2976 2421 3026
rect 2426 2993 2429 3016
rect 2418 2973 2425 2976
rect 2378 2953 2397 2956
rect 2362 2933 2373 2936
rect 2378 2933 2381 2953
rect 2394 2933 2397 2953
rect 2282 2873 2293 2876
rect 2266 2833 2273 2836
rect 2266 2776 2269 2833
rect 2210 2753 2221 2756
rect 2178 2743 2189 2746
rect 2178 2613 2181 2743
rect 2186 2723 2189 2736
rect 2210 2696 2213 2753
rect 2226 2743 2229 2776
rect 2234 2773 2241 2776
rect 2250 2773 2269 2776
rect 2234 2753 2237 2773
rect 2226 2733 2245 2736
rect 2226 2723 2229 2733
rect 2242 2723 2245 2733
rect 2210 2693 2221 2696
rect 2186 2673 2213 2676
rect 2186 2613 2189 2673
rect 2194 2623 2197 2666
rect 2210 2663 2213 2673
rect 2194 2606 2197 2616
rect 2178 2603 2197 2606
rect 2210 2576 2213 2616
rect 2194 2573 2213 2576
rect 2178 2526 2181 2566
rect 2178 2523 2185 2526
rect 2162 2513 2173 2516
rect 2154 2393 2157 2406
rect 2146 2383 2157 2386
rect 2130 2363 2149 2366
rect 2122 2303 2125 2326
rect 2130 2286 2133 2336
rect 2146 2293 2149 2363
rect 2130 2283 2141 2286
rect 2122 2186 2125 2246
rect 2130 2193 2133 2216
rect 2122 2183 2129 2186
rect 2126 2116 2129 2183
rect 2138 2173 2141 2236
rect 2126 2113 2133 2116
rect 2138 2113 2141 2126
rect 2146 2113 2149 2126
rect 2026 1796 2029 1846
rect 2034 1823 2037 1836
rect 2026 1793 2037 1796
rect 2026 1653 2029 1746
rect 2034 1723 2037 1793
rect 2034 1626 2037 1676
rect 2042 1663 2045 1846
rect 2050 1666 2053 1926
rect 2058 1923 2077 1926
rect 2058 1906 2061 1923
rect 2058 1903 2065 1906
rect 2062 1846 2065 1903
rect 2082 1853 2085 1926
rect 2122 1866 2125 2096
rect 2130 1936 2133 2113
rect 2138 2093 2141 2106
rect 2154 1936 2157 2383
rect 2162 2353 2165 2456
rect 2162 2223 2165 2346
rect 2170 2216 2173 2513
rect 2182 2426 2185 2523
rect 2194 2516 2197 2573
rect 2202 2523 2205 2566
rect 2210 2533 2213 2546
rect 2218 2533 2221 2693
rect 2226 2563 2229 2666
rect 2234 2633 2237 2706
rect 2242 2626 2245 2666
rect 2234 2623 2245 2626
rect 2210 2523 2229 2526
rect 2194 2513 2205 2516
rect 2178 2423 2185 2426
rect 2178 2363 2181 2423
rect 2186 2393 2189 2406
rect 2186 2313 2189 2356
rect 2178 2303 2189 2306
rect 2178 2223 2181 2236
rect 2162 2213 2189 2216
rect 2162 2113 2165 2206
rect 2170 2013 2173 2146
rect 2194 2136 2197 2476
rect 2186 2133 2197 2136
rect 2178 2113 2181 2126
rect 2178 2063 2181 2106
rect 2186 2103 2189 2133
rect 2194 2113 2197 2126
rect 2202 2123 2205 2513
rect 2210 2413 2213 2523
rect 2218 2413 2221 2436
rect 2226 2406 2229 2506
rect 2234 2453 2237 2623
rect 2242 2553 2245 2616
rect 2250 2563 2253 2773
rect 2274 2766 2277 2816
rect 2282 2813 2285 2866
rect 2290 2833 2293 2873
rect 2318 2873 2325 2876
rect 2346 2883 2353 2886
rect 2290 2806 2293 2826
rect 2258 2763 2277 2766
rect 2282 2803 2293 2806
rect 2258 2556 2261 2763
rect 2266 2723 2269 2756
rect 2266 2706 2269 2716
rect 2282 2713 2285 2803
rect 2290 2706 2293 2736
rect 2298 2723 2301 2866
rect 2318 2816 2321 2873
rect 2330 2823 2333 2846
rect 2318 2813 2325 2816
rect 2306 2736 2309 2806
rect 2322 2796 2325 2813
rect 2338 2803 2341 2816
rect 2322 2793 2341 2796
rect 2338 2776 2341 2793
rect 2346 2786 2349 2883
rect 2362 2863 2365 2926
rect 2370 2886 2373 2933
rect 2370 2883 2389 2886
rect 2362 2803 2365 2836
rect 2386 2796 2389 2883
rect 2422 2876 2425 2973
rect 2378 2793 2389 2796
rect 2346 2783 2365 2786
rect 2306 2733 2325 2736
rect 2330 2733 2333 2776
rect 2338 2773 2357 2776
rect 2266 2703 2293 2706
rect 2266 2603 2269 2636
rect 2274 2633 2301 2636
rect 2274 2613 2277 2633
rect 2306 2623 2309 2733
rect 2250 2553 2261 2556
rect 2210 2403 2229 2406
rect 2210 2236 2213 2336
rect 2226 2333 2229 2346
rect 2234 2333 2237 2386
rect 2226 2283 2229 2326
rect 2210 2233 2229 2236
rect 2210 2203 2213 2216
rect 2218 2213 2221 2226
rect 2226 2206 2229 2233
rect 2234 2213 2237 2296
rect 2242 2263 2245 2546
rect 2250 2423 2253 2546
rect 2258 2433 2261 2506
rect 2266 2376 2269 2566
rect 2282 2563 2285 2616
rect 2298 2613 2309 2616
rect 2290 2546 2293 2606
rect 2282 2543 2293 2546
rect 2274 2496 2277 2506
rect 2282 2503 2285 2516
rect 2290 2513 2293 2543
rect 2290 2496 2293 2506
rect 2274 2493 2293 2496
rect 2298 2486 2301 2613
rect 2314 2546 2317 2726
rect 2322 2723 2325 2733
rect 2330 2716 2333 2726
rect 2322 2713 2333 2716
rect 2322 2616 2325 2713
rect 2330 2623 2333 2666
rect 2322 2613 2333 2616
rect 2330 2603 2333 2613
rect 2290 2483 2301 2486
rect 2306 2543 2317 2546
rect 2274 2433 2277 2456
rect 2282 2423 2285 2466
rect 2266 2373 2273 2376
rect 2250 2323 2253 2336
rect 2258 2316 2261 2366
rect 2270 2326 2273 2373
rect 2250 2313 2261 2316
rect 2266 2323 2273 2326
rect 2250 2206 2253 2313
rect 2266 2296 2269 2323
rect 2282 2313 2285 2366
rect 2262 2293 2269 2296
rect 2262 2236 2265 2293
rect 2262 2233 2269 2236
rect 2218 2203 2229 2206
rect 2234 2203 2253 2206
rect 2130 1933 2141 1936
rect 2146 1933 2157 1936
rect 2098 1863 2125 1866
rect 2058 1843 2065 1846
rect 2058 1803 2061 1843
rect 2066 1813 2069 1826
rect 2082 1803 2085 1836
rect 2058 1733 2061 1776
rect 2066 1763 2069 1786
rect 2090 1783 2093 1816
rect 2066 1723 2077 1726
rect 2050 1663 2073 1666
rect 2034 1623 2045 1626
rect 2034 1583 2037 1616
rect 1998 1553 2005 1556
rect 1954 1523 1965 1526
rect 1970 1523 1981 1526
rect 1930 1503 1937 1506
rect 1914 1426 1917 1436
rect 1934 1426 1937 1503
rect 1898 1423 1917 1426
rect 1930 1423 1937 1426
rect 1898 1403 1901 1423
rect 1882 1373 1893 1376
rect 1870 1363 1901 1366
rect 1906 1363 1909 1406
rect 1914 1396 1917 1416
rect 1922 1403 1925 1416
rect 1914 1393 1925 1396
rect 1850 1313 1853 1336
rect 1866 1286 1869 1336
rect 1890 1286 1893 1316
rect 1850 1213 1853 1286
rect 1866 1283 1893 1286
rect 1842 1183 1845 1206
rect 1858 1193 1861 1206
rect 1826 1173 1861 1176
rect 1810 1123 1813 1146
rect 1818 1123 1821 1136
rect 1826 1123 1829 1136
rect 1834 1133 1837 1146
rect 1842 1123 1845 1166
rect 1802 1113 1813 1116
rect 1786 1093 1797 1096
rect 1794 1036 1797 1093
rect 1810 1056 1813 1113
rect 1850 1106 1853 1126
rect 1846 1103 1853 1106
rect 1810 1053 1821 1056
rect 1786 1033 1797 1036
rect 1786 1013 1789 1033
rect 1778 1003 1789 1006
rect 1770 983 1777 986
rect 1786 983 1789 1003
rect 1774 856 1777 983
rect 1738 823 1757 826
rect 1754 783 1757 823
rect 1762 776 1765 856
rect 1770 853 1777 856
rect 1770 833 1773 853
rect 1786 816 1789 946
rect 1794 923 1797 1006
rect 1802 966 1805 1016
rect 1810 1003 1813 1036
rect 1802 963 1813 966
rect 1810 873 1813 963
rect 1818 906 1821 1053
rect 1826 1013 1829 1026
rect 1834 1003 1837 1076
rect 1846 986 1849 1103
rect 1858 1003 1861 1173
rect 1866 1126 1869 1276
rect 1874 1203 1877 1246
rect 1882 1176 1885 1216
rect 1874 1173 1885 1176
rect 1874 1133 1877 1173
rect 1866 1123 1877 1126
rect 1874 1096 1877 1123
rect 1866 1013 1869 1096
rect 1874 1093 1881 1096
rect 1878 1026 1881 1093
rect 1890 1086 1893 1283
rect 1898 1273 1901 1363
rect 1914 1323 1917 1336
rect 1898 1213 1909 1216
rect 1898 1183 1901 1206
rect 1914 1203 1917 1266
rect 1914 1123 1917 1156
rect 1922 1143 1925 1206
rect 1930 1086 1933 1423
rect 1946 1413 1949 1426
rect 1938 1333 1941 1406
rect 1954 1393 1957 1406
rect 1946 1306 1949 1376
rect 1954 1333 1957 1366
rect 1942 1303 1949 1306
rect 1942 1236 1945 1303
rect 1942 1233 1949 1236
rect 1938 1123 1941 1216
rect 1946 1213 1949 1233
rect 1890 1083 1901 1086
rect 1930 1083 1937 1086
rect 1954 1083 1957 1286
rect 1874 1023 1881 1026
rect 1874 1006 1877 1023
rect 1870 1003 1877 1006
rect 1846 983 1853 986
rect 1850 966 1853 983
rect 1850 963 1861 966
rect 1858 936 1861 963
rect 1870 936 1873 1003
rect 1842 933 1861 936
rect 1866 933 1873 936
rect 1826 913 1829 926
rect 1818 903 1837 906
rect 1778 813 1789 816
rect 1718 723 1725 726
rect 1730 773 1765 776
rect 1718 626 1721 723
rect 1718 623 1725 626
rect 1706 596 1709 616
rect 1658 593 1709 596
rect 1714 593 1717 606
rect 1634 503 1637 546
rect 1658 526 1661 593
rect 1642 466 1645 526
rect 1634 463 1645 466
rect 1650 523 1661 526
rect 1602 436 1605 456
rect 1602 433 1613 436
rect 1590 423 1597 426
rect 1570 403 1573 416
rect 1546 393 1557 396
rect 1506 383 1517 386
rect 1486 353 1493 356
rect 1482 256 1485 336
rect 1490 323 1493 353
rect 1498 333 1501 356
rect 1514 333 1517 383
rect 1546 376 1549 393
rect 1542 373 1549 376
rect 1482 253 1493 256
rect 1450 186 1453 246
rect 1458 193 1461 206
rect 1466 203 1469 216
rect 1474 203 1477 226
rect 1482 213 1485 236
rect 1490 203 1493 253
rect 1506 213 1509 326
rect 1522 216 1525 346
rect 1530 293 1533 326
rect 1542 246 1545 373
rect 1542 243 1549 246
rect 1514 213 1525 216
rect 1538 213 1541 226
rect 1514 206 1517 213
rect 1506 203 1517 206
rect 1522 203 1533 206
rect 1450 183 1477 186
rect 1458 123 1461 146
rect 1466 113 1469 136
rect 1474 123 1477 183
rect 1498 133 1501 146
rect 1506 123 1509 203
rect 1546 196 1549 243
rect 1538 193 1549 196
rect 1538 133 1541 193
rect 1554 186 1557 376
rect 1570 323 1573 336
rect 1586 333 1589 396
rect 1594 313 1597 423
rect 1610 366 1613 433
rect 1602 363 1613 366
rect 1634 366 1637 463
rect 1650 413 1653 523
rect 1666 516 1669 536
rect 1682 533 1685 546
rect 1658 413 1661 516
rect 1666 513 1673 516
rect 1670 436 1673 513
rect 1666 433 1673 436
rect 1666 413 1669 433
rect 1634 363 1645 366
rect 1570 203 1573 286
rect 1554 183 1573 186
rect 1570 123 1573 183
rect 1594 123 1597 146
rect 1602 63 1605 363
rect 1642 346 1645 363
rect 1650 356 1653 406
rect 1658 403 1669 406
rect 1650 353 1661 356
rect 1610 343 1653 346
rect 1610 323 1613 343
rect 1618 323 1621 336
rect 1634 316 1637 336
rect 1650 333 1653 343
rect 1630 313 1637 316
rect 1630 256 1633 313
rect 1642 303 1645 326
rect 1618 253 1633 256
rect 1618 213 1621 253
rect 1650 213 1653 326
rect 1658 213 1661 353
rect 1666 203 1669 396
rect 1674 316 1677 416
rect 1682 386 1685 446
rect 1690 433 1693 526
rect 1698 513 1701 536
rect 1706 506 1709 593
rect 1722 513 1725 623
rect 1702 503 1709 506
rect 1702 446 1705 503
rect 1698 443 1705 446
rect 1698 403 1701 443
rect 1714 403 1717 466
rect 1730 443 1733 773
rect 1738 733 1741 746
rect 1746 733 1757 736
rect 1762 726 1765 736
rect 1746 723 1765 726
rect 1746 693 1749 723
rect 1746 616 1749 676
rect 1738 613 1749 616
rect 1754 613 1757 646
rect 1770 626 1773 806
rect 1794 803 1797 836
rect 1786 733 1789 786
rect 1770 623 1781 626
rect 1746 553 1749 606
rect 1770 583 1773 616
rect 1778 566 1781 623
rect 1786 603 1789 636
rect 1794 613 1797 726
rect 1802 643 1805 826
rect 1818 803 1821 866
rect 1842 753 1845 933
rect 1850 913 1853 926
rect 1858 826 1861 906
rect 1866 853 1869 933
rect 1882 926 1885 1006
rect 1898 943 1901 1083
rect 1890 933 1901 936
rect 1882 923 1901 926
rect 1874 903 1877 916
rect 1882 856 1885 916
rect 1882 853 1889 856
rect 1858 823 1865 826
rect 1810 693 1813 736
rect 1834 733 1837 746
rect 1850 743 1853 816
rect 1862 756 1865 823
rect 1886 796 1889 853
rect 1882 793 1889 796
rect 1882 773 1885 793
rect 1898 783 1901 923
rect 1906 913 1909 926
rect 1906 803 1909 856
rect 1914 823 1917 966
rect 1922 933 1925 1076
rect 1934 1006 1937 1083
rect 1930 1003 1937 1006
rect 1930 833 1933 1003
rect 1938 933 1941 986
rect 1946 963 1949 1016
rect 1962 993 1965 1523
rect 1986 1506 1989 1536
rect 1982 1503 1989 1506
rect 1970 1403 1973 1446
rect 1982 1426 1985 1503
rect 1982 1423 1989 1426
rect 1970 1253 1973 1396
rect 1978 1243 1981 1406
rect 1986 1313 1989 1423
rect 1994 1393 1997 1536
rect 2002 1496 2005 1553
rect 2018 1533 2021 1576
rect 2042 1533 2045 1623
rect 2058 1613 2061 1656
rect 2042 1496 2045 1526
rect 2002 1493 2013 1496
rect 2010 1436 2013 1493
rect 2002 1433 2013 1436
rect 2034 1493 2045 1496
rect 1994 1256 1997 1376
rect 2002 1346 2005 1433
rect 2010 1393 2013 1416
rect 2018 1363 2021 1406
rect 2026 1366 2029 1416
rect 2034 1403 2037 1493
rect 2050 1463 2053 1606
rect 2026 1363 2037 1366
rect 2002 1343 2025 1346
rect 1986 1253 1997 1256
rect 2002 1253 2005 1336
rect 2010 1323 2013 1336
rect 1970 1186 1973 1226
rect 1978 1193 1981 1216
rect 1970 1183 1981 1186
rect 1970 1123 1973 1146
rect 1978 1123 1981 1183
rect 1970 1013 1981 1016
rect 1986 1006 1989 1253
rect 1994 1093 1997 1246
rect 2002 1203 2005 1216
rect 2010 1213 2013 1276
rect 2022 1226 2025 1343
rect 2034 1283 2037 1363
rect 2042 1333 2045 1426
rect 2050 1393 2053 1406
rect 2050 1333 2053 1366
rect 2022 1223 2029 1226
rect 2018 1193 2021 1206
rect 2026 1186 2029 1223
rect 2034 1203 2037 1246
rect 2042 1196 2045 1276
rect 2058 1266 2061 1596
rect 2070 1566 2073 1663
rect 2066 1563 2073 1566
rect 2066 1453 2069 1563
rect 2082 1476 2085 1736
rect 2078 1473 2085 1476
rect 2078 1396 2081 1473
rect 2090 1403 2093 1726
rect 2098 1673 2101 1863
rect 2106 1706 2109 1806
rect 2114 1803 2117 1826
rect 2122 1786 2125 1856
rect 2130 1793 2133 1926
rect 2122 1783 2133 1786
rect 2130 1733 2133 1783
rect 2138 1733 2141 1933
rect 2146 1793 2149 1926
rect 2154 1916 2157 1933
rect 2154 1913 2161 1916
rect 2158 1856 2161 1913
rect 2154 1853 2161 1856
rect 2154 1836 2157 1853
rect 2154 1833 2165 1836
rect 2154 1813 2157 1833
rect 2162 1783 2165 1806
rect 2146 1733 2157 1736
rect 2114 1723 2125 1726
rect 2106 1703 2113 1706
rect 2110 1626 2113 1703
rect 2122 1676 2125 1723
rect 2138 1703 2141 1726
rect 2122 1673 2141 1676
rect 2110 1623 2117 1626
rect 2098 1593 2101 1606
rect 2106 1583 2109 1616
rect 2098 1443 2101 1526
rect 2114 1443 2117 1623
rect 2122 1603 2125 1673
rect 2078 1393 2085 1396
rect 2066 1273 2069 1366
rect 2082 1336 2085 1393
rect 2078 1333 2085 1336
rect 2002 1183 2029 1186
rect 2034 1193 2045 1196
rect 2050 1263 2061 1266
rect 1978 1003 1989 1006
rect 1946 863 1949 946
rect 1938 813 1941 856
rect 1906 793 1917 796
rect 1946 783 1949 816
rect 1954 803 1957 936
rect 1962 933 1965 946
rect 1962 873 1965 926
rect 1970 903 1973 926
rect 1978 923 1981 1003
rect 1986 953 1989 986
rect 1986 916 1989 946
rect 1978 913 1989 916
rect 1962 786 1965 816
rect 1970 803 1973 826
rect 1978 793 1981 913
rect 1986 786 1989 836
rect 1994 823 1997 1016
rect 1962 783 1989 786
rect 1858 753 1865 756
rect 1826 706 1829 726
rect 1842 723 1845 736
rect 1826 703 1833 706
rect 1850 703 1853 736
rect 1818 643 1821 676
rect 1830 646 1833 703
rect 1830 643 1845 646
rect 1802 613 1821 616
rect 1802 596 1805 613
rect 1786 593 1805 596
rect 1778 563 1789 566
rect 1746 463 1749 536
rect 1770 523 1773 546
rect 1738 396 1741 416
rect 1730 393 1741 396
rect 1682 383 1693 386
rect 1690 376 1693 383
rect 1682 333 1685 376
rect 1690 373 1725 376
rect 1698 316 1701 336
rect 1674 313 1681 316
rect 1678 236 1681 313
rect 1690 313 1701 316
rect 1714 316 1717 326
rect 1722 323 1725 373
rect 1730 333 1733 393
rect 1778 356 1781 556
rect 1786 403 1789 563
rect 1794 543 1797 586
rect 1802 566 1805 593
rect 1810 586 1813 606
rect 1826 593 1829 606
rect 1810 583 1837 586
rect 1802 563 1821 566
rect 1794 373 1797 536
rect 1802 403 1805 416
rect 1770 353 1781 356
rect 1738 323 1741 346
rect 1746 316 1749 336
rect 1714 313 1749 316
rect 1690 293 1693 313
rect 1674 233 1681 236
rect 1674 203 1677 233
rect 1682 173 1685 216
rect 1706 213 1709 306
rect 1770 296 1773 353
rect 1762 293 1773 296
rect 1762 236 1765 293
rect 1762 233 1773 236
rect 1650 123 1653 156
rect 1674 133 1677 166
rect 1698 123 1701 206
rect 1746 176 1749 206
rect 1762 203 1765 216
rect 1770 213 1773 233
rect 1746 173 1757 176
rect 1778 173 1781 216
rect 1754 123 1757 173
rect 1786 133 1789 336
rect 1810 293 1813 546
rect 1818 496 1821 563
rect 1826 513 1829 526
rect 1818 493 1825 496
rect 1834 493 1837 536
rect 1822 436 1825 493
rect 1842 486 1845 643
rect 1858 603 1861 753
rect 1866 693 1869 736
rect 1882 673 1885 726
rect 1850 556 1853 596
rect 1874 583 1877 616
rect 1882 613 1885 666
rect 1882 593 1885 606
rect 1850 553 1869 556
rect 1866 533 1869 553
rect 1834 483 1845 486
rect 1822 433 1829 436
rect 1802 146 1805 206
rect 1810 203 1813 216
rect 1818 173 1821 416
rect 1826 406 1829 433
rect 1834 413 1837 483
rect 1850 413 1853 436
rect 1826 403 1837 406
rect 1826 323 1829 386
rect 1834 213 1837 403
rect 1842 383 1845 406
rect 1858 403 1861 526
rect 1874 523 1877 556
rect 1890 516 1893 756
rect 1898 733 1901 746
rect 1906 706 1909 736
rect 1938 733 1941 756
rect 1970 733 1973 776
rect 1906 703 1917 706
rect 1898 596 1901 676
rect 1914 603 1917 703
rect 1922 603 1925 636
rect 1898 593 1917 596
rect 1914 546 1917 593
rect 1914 543 1921 546
rect 1874 513 1893 516
rect 1874 346 1877 513
rect 1898 503 1901 536
rect 1906 496 1909 536
rect 1898 493 1909 496
rect 1918 486 1921 543
rect 1930 533 1933 626
rect 1946 613 1949 726
rect 1954 583 1957 606
rect 1938 533 1941 556
rect 1930 516 1933 526
rect 1938 523 1949 526
rect 1930 513 1949 516
rect 1914 483 1921 486
rect 1882 413 1893 416
rect 1890 403 1893 413
rect 1914 406 1917 483
rect 1938 413 1941 436
rect 1898 403 1917 406
rect 1866 343 1877 346
rect 1866 323 1869 343
rect 1874 286 1877 336
rect 1866 283 1877 286
rect 1866 226 1869 283
rect 1882 246 1885 326
rect 1898 323 1901 403
rect 1930 393 1933 406
rect 1906 333 1909 346
rect 1882 243 1893 246
rect 1866 223 1885 226
rect 1842 203 1869 206
rect 1874 203 1877 216
rect 1802 143 1813 146
rect 1810 123 1813 143
rect 1866 123 1869 203
rect 1874 123 1877 176
rect 1882 133 1885 223
rect 1890 213 1893 243
rect 1898 193 1901 206
rect 1906 203 1909 216
rect 1906 133 1909 146
rect 1914 123 1917 336
rect 1938 196 1941 406
rect 1946 403 1949 513
rect 1954 503 1957 536
rect 1962 486 1965 616
rect 1970 593 1973 606
rect 1978 533 1981 636
rect 1986 613 1989 656
rect 1994 626 1997 786
rect 2002 683 2005 1183
rect 2034 1156 2037 1193
rect 2050 1156 2053 1263
rect 2078 1256 2081 1333
rect 2090 1283 2093 1326
rect 2018 1153 2037 1156
rect 2042 1153 2053 1156
rect 2058 1253 2081 1256
rect 2010 1133 2013 1146
rect 2018 1123 2021 1153
rect 2026 1123 2037 1126
rect 2010 993 2013 1016
rect 2018 1013 2021 1096
rect 2042 1026 2045 1153
rect 2050 1133 2053 1146
rect 2058 1033 2061 1253
rect 2066 1133 2069 1186
rect 2074 1166 2077 1206
rect 2074 1163 2093 1166
rect 2042 1023 2061 1026
rect 2026 1013 2045 1016
rect 2018 983 2021 1006
rect 2026 976 2029 1013
rect 2018 973 2029 976
rect 2010 913 2013 936
rect 2018 893 2021 973
rect 2034 963 2037 1006
rect 2026 903 2029 936
rect 2026 843 2029 856
rect 2010 706 2013 836
rect 2026 783 2029 806
rect 2034 763 2037 816
rect 2018 723 2021 746
rect 2010 703 2017 706
rect 2014 646 2017 703
rect 2042 663 2045 1006
rect 2050 993 2053 1006
rect 2058 1003 2061 1023
rect 2074 1013 2077 1126
rect 2082 1093 2085 1136
rect 2090 1006 2093 1163
rect 2098 1116 2101 1396
rect 2106 1343 2109 1436
rect 2114 1333 2117 1416
rect 2122 1406 2125 1596
rect 2130 1413 2133 1616
rect 2138 1556 2141 1673
rect 2146 1563 2149 1733
rect 2162 1723 2165 1756
rect 2154 1656 2157 1676
rect 2154 1653 2161 1656
rect 2158 1556 2161 1653
rect 2138 1553 2149 1556
rect 2138 1453 2141 1546
rect 2146 1523 2149 1553
rect 2154 1553 2161 1556
rect 2138 1426 2141 1446
rect 2154 1443 2157 1553
rect 2138 1423 2149 1426
rect 2122 1403 2133 1406
rect 2122 1293 2125 1396
rect 2130 1323 2133 1403
rect 2146 1356 2149 1423
rect 2162 1413 2165 1536
rect 2162 1393 2165 1406
rect 2138 1353 2149 1356
rect 2138 1316 2141 1353
rect 2146 1333 2157 1336
rect 2130 1313 2141 1316
rect 2106 1153 2109 1276
rect 2114 1213 2117 1256
rect 2106 1123 2109 1146
rect 2114 1123 2117 1136
rect 2098 1113 2109 1116
rect 2074 1003 2093 1006
rect 2074 996 2077 1003
rect 2058 993 2077 996
rect 2058 773 2061 993
rect 2082 936 2085 996
rect 2106 966 2109 1113
rect 2122 1093 2125 1266
rect 2138 1236 2141 1256
rect 2138 1233 2145 1236
rect 2142 1176 2145 1233
rect 2138 1173 2145 1176
rect 2138 1106 2141 1173
rect 2154 1133 2157 1326
rect 2162 1323 2165 1356
rect 2162 1213 2165 1276
rect 2170 1173 2173 1966
rect 2178 1893 2181 2036
rect 2210 2026 2213 2116
rect 2218 2113 2221 2203
rect 2226 2103 2229 2146
rect 2234 2083 2237 2203
rect 2258 2186 2261 2216
rect 2242 2183 2261 2186
rect 2242 2113 2245 2183
rect 2266 2176 2269 2233
rect 2250 2173 2269 2176
rect 2250 2096 2253 2173
rect 2274 2143 2277 2306
rect 2282 2233 2285 2306
rect 2290 2233 2293 2483
rect 2306 2456 2309 2543
rect 2314 2473 2317 2526
rect 2330 2513 2333 2546
rect 2298 2423 2301 2456
rect 2306 2453 2317 2456
rect 2306 2416 2309 2436
rect 2322 2433 2325 2506
rect 2338 2433 2341 2773
rect 2346 2723 2349 2736
rect 2354 2723 2357 2773
rect 2362 2676 2365 2783
rect 2346 2673 2365 2676
rect 2314 2423 2325 2426
rect 2306 2413 2317 2416
rect 2306 2323 2309 2413
rect 2322 2396 2325 2423
rect 2330 2403 2333 2426
rect 2346 2406 2349 2673
rect 2370 2666 2373 2756
rect 2362 2663 2373 2666
rect 2378 2656 2381 2793
rect 2394 2786 2397 2876
rect 2418 2873 2425 2876
rect 2418 2856 2421 2873
rect 2434 2856 2437 3036
rect 2458 3033 2477 3036
rect 2450 2996 2453 3016
rect 2458 3003 2461 3033
rect 2466 2996 2469 3016
rect 2450 2993 2469 2996
rect 2458 2966 2461 2986
rect 2458 2963 2465 2966
rect 2474 2963 2477 3026
rect 2482 3013 2485 3026
rect 2498 3023 2501 3043
rect 2506 2993 2509 3026
rect 2538 3023 2549 3026
rect 2530 3013 2541 3016
rect 2530 2983 2533 3013
rect 2538 2996 2541 3006
rect 2546 3003 2549 3023
rect 2554 3013 2557 3026
rect 2562 2996 2565 3036
rect 2570 3013 2573 3026
rect 2586 3016 2589 3036
rect 2594 3023 2597 3073
rect 2602 3016 2605 3106
rect 2610 3033 2613 3126
rect 2626 3083 2629 3116
rect 2634 3096 2637 3133
rect 2642 3123 2645 3366
rect 2650 3313 2653 3386
rect 2658 3383 2669 3386
rect 2658 3343 2661 3383
rect 2666 3343 2669 3376
rect 2666 3326 2669 3336
rect 2674 3333 2677 3723
rect 2682 3603 2685 3706
rect 2690 3663 2693 3726
rect 2690 3623 2693 3656
rect 2698 3606 2701 3746
rect 2706 3663 2709 3753
rect 2706 3613 2709 3626
rect 2714 3613 2717 3646
rect 2722 3606 2725 3736
rect 2730 3673 2733 3763
rect 2738 3723 2741 3766
rect 2746 3723 2749 3746
rect 2690 3603 2701 3606
rect 2706 3603 2725 3606
rect 2690 3586 2693 3603
rect 2682 3583 2693 3586
rect 2682 3533 2685 3583
rect 2690 3523 2693 3546
rect 2682 3513 2693 3516
rect 2682 3333 2685 3506
rect 2690 3493 2693 3513
rect 2690 3353 2693 3416
rect 2698 3396 2701 3536
rect 2706 3493 2709 3526
rect 2714 3476 2717 3566
rect 2730 3553 2733 3666
rect 2738 3623 2741 3706
rect 2746 3603 2749 3626
rect 2754 3603 2757 3903
rect 2762 3823 2765 3846
rect 2762 3803 2765 3816
rect 2762 3733 2765 3766
rect 2770 3726 2773 3946
rect 2786 3936 2789 3956
rect 2778 3923 2781 3936
rect 2786 3933 2797 3936
rect 2794 3893 2797 3926
rect 2802 3923 2805 3946
rect 2810 3823 2813 3993
rect 2818 3916 2821 3986
rect 2834 3933 2837 3966
rect 2842 3923 2845 3956
rect 2850 3933 2853 3976
rect 2874 3936 2877 3956
rect 2890 3953 2893 4016
rect 2818 3913 2829 3916
rect 2826 3836 2829 3913
rect 2850 3896 2853 3926
rect 2858 3923 2861 3936
rect 2866 3926 2869 3936
rect 2874 3933 2893 3936
rect 2898 3933 2901 3986
rect 2906 3966 2909 4096
rect 2914 3976 2917 4016
rect 2930 3983 2933 4143
rect 2942 4036 2945 4173
rect 2954 4103 2957 4126
rect 2994 4123 2997 4206
rect 3010 4203 3013 4216
rect 3018 4163 3021 4216
rect 3026 4203 3029 4296
rect 3034 4203 3037 4216
rect 3042 4213 3045 4306
rect 3050 4203 3053 4276
rect 3058 4236 3061 4340
rect 3082 4293 3085 4340
rect 3098 4286 3101 4340
rect 3258 4326 3261 4340
rect 3298 4326 3301 4340
rect 3250 4323 3261 4326
rect 3274 4323 3301 4326
rect 3074 4283 3101 4286
rect 3058 4233 3069 4236
rect 3034 4193 3045 4196
rect 3010 4133 3013 4146
rect 2938 4033 2945 4036
rect 2914 3973 2933 3976
rect 2906 3963 2917 3966
rect 2866 3923 2877 3926
rect 2890 3916 2893 3933
rect 2886 3913 2893 3916
rect 2850 3893 2861 3896
rect 2818 3833 2829 3836
rect 2786 3805 2789 3816
rect 2810 3766 2813 3816
rect 2778 3733 2781 3766
rect 2794 3763 2813 3766
rect 2818 3763 2821 3833
rect 2794 3733 2797 3763
rect 2810 3743 2829 3746
rect 2810 3733 2813 3743
rect 2770 3723 2781 3726
rect 2786 3716 2789 3726
rect 2794 3723 2805 3726
rect 2818 3716 2821 3736
rect 2826 3723 2829 3743
rect 2834 3723 2837 3796
rect 2850 3776 2853 3886
rect 2842 3773 2853 3776
rect 2762 3706 2765 3716
rect 2786 3713 2821 3716
rect 2762 3703 2797 3706
rect 2762 3693 2765 3703
rect 2746 3563 2749 3596
rect 2706 3473 2717 3476
rect 2722 3473 2725 3526
rect 2706 3403 2709 3473
rect 2714 3423 2717 3466
rect 2722 3413 2725 3426
rect 2714 3396 2717 3406
rect 2698 3393 2717 3396
rect 2666 3323 2685 3326
rect 2690 3316 2693 3346
rect 2658 3313 2693 3316
rect 2650 3283 2653 3306
rect 2650 3203 2653 3226
rect 2658 3193 2661 3313
rect 2674 3293 2701 3296
rect 2650 3116 2653 3136
rect 2650 3113 2657 3116
rect 2634 3093 2645 3096
rect 2618 3043 2621 3066
rect 2538 2993 2565 2996
rect 2410 2853 2421 2856
rect 2430 2853 2437 2856
rect 2402 2813 2405 2826
rect 2386 2783 2397 2786
rect 2386 2723 2389 2783
rect 2410 2746 2413 2853
rect 2430 2766 2433 2853
rect 2442 2843 2445 2926
rect 2462 2886 2465 2963
rect 2578 2936 2581 3016
rect 2586 3013 2605 3016
rect 2610 3016 2613 3026
rect 2610 3013 2621 3016
rect 2626 3013 2629 3036
rect 2602 2936 2605 3006
rect 2474 2906 2477 2926
rect 2474 2903 2485 2906
rect 2506 2903 2509 2936
rect 2578 2933 2605 2936
rect 2618 2933 2621 3013
rect 2634 2926 2637 3093
rect 2642 3083 2645 3093
rect 2654 3046 2657 3113
rect 2650 3043 2657 3046
rect 2642 3016 2645 3036
rect 2650 3023 2653 3043
rect 2642 3013 2653 3016
rect 2650 2996 2653 3013
rect 2666 3003 2669 3226
rect 2674 3166 2677 3293
rect 2682 3213 2685 3256
rect 2706 3243 2709 3336
rect 2714 3236 2717 3393
rect 2690 3233 2717 3236
rect 2682 3173 2685 3206
rect 2690 3203 2693 3233
rect 2722 3226 2725 3336
rect 2698 3223 2709 3226
rect 2714 3223 2725 3226
rect 2714 3173 2717 3223
rect 2722 3203 2725 3216
rect 2674 3163 2701 3166
rect 2698 3146 2701 3163
rect 2698 3143 2705 3146
rect 2682 3116 2685 3126
rect 2674 3043 2677 3116
rect 2682 3113 2693 3116
rect 2674 3013 2677 3026
rect 2682 3003 2685 3106
rect 2690 3036 2693 3113
rect 2702 3076 2705 3143
rect 2730 3123 2733 3546
rect 2738 3503 2741 3536
rect 2738 3413 2741 3466
rect 2746 3403 2749 3526
rect 2754 3523 2757 3586
rect 2738 3333 2741 3376
rect 2754 3373 2757 3486
rect 2762 3403 2765 3636
rect 2770 3613 2773 3626
rect 2778 3613 2781 3686
rect 2786 3606 2789 3626
rect 2794 3623 2797 3703
rect 2810 3626 2813 3713
rect 2826 3706 2829 3716
rect 2818 3703 2829 3706
rect 2818 3633 2821 3703
rect 2778 3586 2781 3606
rect 2786 3603 2797 3606
rect 2802 3586 2805 3626
rect 2810 3623 2821 3626
rect 2778 3583 2805 3586
rect 2770 3533 2773 3566
rect 2778 3526 2781 3576
rect 2770 3523 2781 3526
rect 2786 3523 2789 3583
rect 2818 3536 2821 3623
rect 2834 3613 2837 3636
rect 2826 3543 2829 3566
rect 2842 3553 2845 3773
rect 2858 3766 2861 3893
rect 2886 3846 2889 3913
rect 2886 3843 2893 3846
rect 2866 3813 2869 3826
rect 2850 3763 2861 3766
rect 2850 3733 2853 3763
rect 2866 3733 2869 3806
rect 2858 3723 2869 3726
rect 2874 3723 2877 3816
rect 2882 3803 2885 3826
rect 2890 3746 2893 3843
rect 2898 3753 2901 3926
rect 2906 3866 2909 3956
rect 2914 3933 2917 3963
rect 2930 3933 2933 3973
rect 2938 3933 2941 4033
rect 2946 3983 2949 4016
rect 2954 3953 2957 3996
rect 2962 3966 2965 4006
rect 2970 3973 2973 4016
rect 2978 4003 2981 4096
rect 2986 3966 2989 4016
rect 2994 4003 2997 4106
rect 3002 4013 3005 4126
rect 3010 3973 3013 4006
rect 3018 3983 3021 4136
rect 3026 4133 3029 4186
rect 3034 4056 3037 4193
rect 3058 4163 3061 4216
rect 3066 4203 3069 4233
rect 3074 4203 3077 4283
rect 3146 4236 3149 4256
rect 3138 4233 3149 4236
rect 3082 4193 3085 4216
rect 3098 4186 3101 4206
rect 3122 4186 3125 4216
rect 3082 4183 3101 4186
rect 3114 4183 3125 4186
rect 3042 4126 3045 4136
rect 3050 4133 3061 4136
rect 3042 4123 3053 4126
rect 3082 4123 3085 4183
rect 3138 4176 3141 4233
rect 3138 4173 3149 4176
rect 3146 4156 3149 4173
rect 3146 4153 3153 4156
rect 3026 4053 3037 4056
rect 3026 4003 3029 4053
rect 3034 4033 3045 4036
rect 3050 4013 3061 4016
rect 3026 3973 3045 3976
rect 2962 3963 2989 3966
rect 2946 3943 2965 3946
rect 2946 3933 2949 3943
rect 2922 3876 2925 3926
rect 2938 3883 2941 3926
rect 2954 3876 2957 3936
rect 2962 3923 2965 3943
rect 2922 3873 2957 3876
rect 2906 3863 2917 3866
rect 2914 3803 2917 3863
rect 2946 3826 2949 3873
rect 2946 3823 2957 3826
rect 2978 3823 2981 3936
rect 2986 3916 2989 3963
rect 2994 3933 2997 3956
rect 2986 3913 2993 3916
rect 2990 3846 2993 3913
rect 3002 3863 3005 3926
rect 3010 3913 3013 3936
rect 2986 3843 2993 3846
rect 2938 3803 2941 3816
rect 2914 3763 2917 3786
rect 2954 3776 2957 3823
rect 2986 3776 2989 3843
rect 2994 3813 2997 3826
rect 2922 3773 2957 3776
rect 2970 3773 2989 3776
rect 2890 3743 2909 3746
rect 2882 3726 2885 3736
rect 2890 3733 2901 3736
rect 2882 3723 2893 3726
rect 2898 3723 2901 3733
rect 2850 3623 2853 3656
rect 2858 3633 2861 3723
rect 2906 3716 2909 3743
rect 2866 3616 2869 3716
rect 2890 3713 2909 3716
rect 2850 3613 2869 3616
rect 2794 3523 2797 3536
rect 2770 3506 2773 3523
rect 2802 3516 2805 3526
rect 2778 3513 2805 3516
rect 2770 3503 2781 3506
rect 2770 3396 2773 3406
rect 2778 3403 2781 3503
rect 2802 3423 2805 3506
rect 2810 3416 2813 3536
rect 2818 3533 2825 3536
rect 2834 3533 2845 3536
rect 2822 3456 2825 3533
rect 2834 3456 2837 3526
rect 2842 3513 2845 3533
rect 2822 3453 2829 3456
rect 2834 3453 2845 3456
rect 2794 3413 2813 3416
rect 2770 3393 2781 3396
rect 2746 3343 2773 3346
rect 2738 3303 2741 3326
rect 2746 3313 2749 3343
rect 2754 3303 2757 3336
rect 2762 3306 2765 3336
rect 2770 3323 2773 3343
rect 2778 3333 2781 3393
rect 2778 3323 2789 3326
rect 2794 3316 2797 3413
rect 2786 3313 2797 3316
rect 2762 3303 2773 3306
rect 2738 3243 2741 3286
rect 2738 3203 2741 3216
rect 2746 3186 2749 3216
rect 2762 3186 2765 3206
rect 2770 3193 2773 3303
rect 2778 3213 2781 3226
rect 2786 3186 2789 3313
rect 2802 3306 2805 3406
rect 2818 3403 2821 3436
rect 2826 3403 2829 3453
rect 2834 3413 2837 3436
rect 2818 3343 2821 3396
rect 2834 3393 2837 3406
rect 2842 3346 2845 3453
rect 2850 3403 2853 3613
rect 2874 3606 2877 3616
rect 2882 3613 2885 3646
rect 2858 3603 2877 3606
rect 2858 3533 2861 3596
rect 2882 3576 2885 3606
rect 2890 3603 2893 3713
rect 2898 3663 2901 3706
rect 2914 3666 2917 3736
rect 2922 3706 2925 3773
rect 2930 3726 2933 3746
rect 2930 3723 2941 3726
rect 2946 3716 2949 3766
rect 2954 3743 2957 3756
rect 2954 3733 2965 3736
rect 2970 3733 2973 3773
rect 2962 3726 2965 3733
rect 2962 3723 2973 3726
rect 2978 3716 2981 3746
rect 2938 3713 2949 3716
rect 2922 3703 2941 3706
rect 2906 3663 2917 3666
rect 2906 3646 2909 3663
rect 2898 3643 2909 3646
rect 2898 3603 2901 3643
rect 2906 3583 2909 3626
rect 2882 3573 2909 3576
rect 2858 3523 2869 3526
rect 2882 3523 2885 3536
rect 2834 3343 2845 3346
rect 2798 3303 2805 3306
rect 2798 3246 2801 3303
rect 2746 3183 2757 3186
rect 2762 3183 2789 3186
rect 2794 3243 2801 3246
rect 2698 3073 2705 3076
rect 2714 3083 2725 3086
rect 2698 3053 2701 3073
rect 2690 3033 2709 3036
rect 2698 3013 2701 3033
rect 2706 3013 2709 3026
rect 2714 3003 2717 3083
rect 2738 3056 2741 3136
rect 2746 3123 2749 3176
rect 2754 3123 2757 3183
rect 2794 3176 2797 3243
rect 2802 3213 2805 3226
rect 2762 3173 2797 3176
rect 2762 3126 2765 3173
rect 2770 3133 2781 3136
rect 2762 3123 2769 3126
rect 2738 3053 2749 3056
rect 2458 2883 2465 2886
rect 2458 2866 2461 2883
rect 2450 2863 2461 2866
rect 2442 2773 2445 2816
rect 2450 2766 2453 2863
rect 2430 2763 2437 2766
rect 2394 2743 2413 2746
rect 2394 2706 2397 2743
rect 2362 2653 2381 2656
rect 2390 2703 2397 2706
rect 2354 2613 2357 2636
rect 2362 2606 2365 2653
rect 2390 2646 2393 2703
rect 2378 2643 2393 2646
rect 2354 2603 2365 2606
rect 2354 2536 2357 2603
rect 2362 2563 2365 2596
rect 2370 2556 2373 2606
rect 2378 2563 2381 2643
rect 2402 2636 2405 2736
rect 2418 2723 2421 2756
rect 2434 2746 2437 2763
rect 2426 2743 2437 2746
rect 2434 2733 2437 2743
rect 2442 2763 2453 2766
rect 2402 2633 2413 2636
rect 2394 2613 2397 2626
rect 2402 2586 2405 2616
rect 2386 2583 2405 2586
rect 2362 2553 2381 2556
rect 2362 2543 2365 2553
rect 2354 2533 2361 2536
rect 2358 2476 2361 2533
rect 2358 2473 2365 2476
rect 2342 2403 2349 2406
rect 2322 2393 2333 2396
rect 2314 2316 2317 2356
rect 2298 2283 2301 2316
rect 2306 2313 2317 2316
rect 2282 2213 2285 2226
rect 2282 2136 2285 2176
rect 2298 2156 2301 2226
rect 2306 2173 2309 2313
rect 2314 2273 2317 2306
rect 2322 2253 2325 2346
rect 2330 2223 2333 2393
rect 2342 2336 2345 2403
rect 2342 2333 2349 2336
rect 2338 2303 2341 2316
rect 2346 2306 2349 2333
rect 2354 2313 2357 2456
rect 2346 2303 2357 2306
rect 2354 2283 2357 2303
rect 2298 2153 2317 2156
rect 2274 2133 2285 2136
rect 2274 2116 2277 2133
rect 2282 2123 2293 2126
rect 2246 2093 2253 2096
rect 2246 2026 2249 2093
rect 2258 2053 2261 2116
rect 2274 2113 2285 2116
rect 2266 2033 2269 2096
rect 2274 2083 2277 2106
rect 2186 2023 2197 2026
rect 2210 2023 2237 2026
rect 2246 2023 2253 2026
rect 2186 1936 2189 2023
rect 2194 2013 2213 2016
rect 2194 2003 2197 2013
rect 2202 1983 2205 2006
rect 2210 2003 2229 2006
rect 2186 1933 2197 1936
rect 2178 1813 2181 1836
rect 2186 1743 2189 1926
rect 2178 1673 2181 1736
rect 2186 1653 2189 1736
rect 2194 1706 2197 1933
rect 2202 1913 2205 1926
rect 2202 1726 2205 1826
rect 2210 1813 2213 2003
rect 2234 1976 2237 2023
rect 2226 1973 2237 1976
rect 2226 1926 2229 1973
rect 2242 1933 2245 1966
rect 2250 1943 2253 2023
rect 2226 1923 2237 1926
rect 2218 1753 2221 1896
rect 2210 1733 2221 1736
rect 2202 1723 2213 1726
rect 2218 1723 2221 1733
rect 2194 1703 2205 1706
rect 2202 1646 2205 1703
rect 2226 1656 2229 1806
rect 2178 1643 2205 1646
rect 2218 1653 2229 1656
rect 2178 1613 2181 1643
rect 2194 1573 2197 1606
rect 2202 1593 2205 1616
rect 2186 1546 2189 1566
rect 2178 1403 2181 1546
rect 2186 1543 2193 1546
rect 2218 1543 2221 1653
rect 2226 1603 2229 1646
rect 2190 1456 2193 1543
rect 2202 1503 2205 1536
rect 2210 1523 2213 1536
rect 2218 1533 2229 1536
rect 2186 1453 2193 1456
rect 2178 1243 2181 1356
rect 2186 1323 2189 1453
rect 2194 1403 2197 1436
rect 2186 1203 2189 1316
rect 2202 1243 2205 1376
rect 2210 1163 2213 1446
rect 2218 1413 2221 1533
rect 2234 1516 2237 1923
rect 2250 1863 2253 1926
rect 2258 1916 2261 2016
rect 2266 2013 2269 2026
rect 2274 1933 2277 2066
rect 2282 1983 2285 2113
rect 2298 2103 2301 2146
rect 2290 2003 2293 2036
rect 2298 2033 2301 2086
rect 2306 2016 2309 2116
rect 2302 2013 2309 2016
rect 2282 1923 2285 1936
rect 2258 1913 2269 1916
rect 2290 1913 2293 1926
rect 2302 1916 2305 2013
rect 2314 1973 2317 2153
rect 2330 2136 2333 2186
rect 2338 2173 2341 2256
rect 2346 2203 2349 2226
rect 2354 2186 2357 2216
rect 2346 2183 2357 2186
rect 2330 2133 2341 2136
rect 2322 2016 2325 2126
rect 2346 2123 2349 2183
rect 2354 2116 2357 2176
rect 2338 2113 2357 2116
rect 2338 2096 2341 2113
rect 2362 2106 2365 2473
rect 2370 2416 2373 2536
rect 2378 2533 2381 2553
rect 2386 2533 2389 2583
rect 2410 2576 2413 2633
rect 2402 2573 2413 2576
rect 2378 2433 2381 2456
rect 2370 2413 2377 2416
rect 2374 2356 2377 2413
rect 2386 2373 2389 2436
rect 2370 2353 2377 2356
rect 2370 2336 2373 2353
rect 2370 2333 2389 2336
rect 2370 2273 2373 2306
rect 2378 2293 2381 2316
rect 2370 2203 2373 2226
rect 2386 2223 2389 2333
rect 2370 2133 2373 2146
rect 2334 2093 2341 2096
rect 2334 2036 2337 2093
rect 2346 2083 2349 2106
rect 2358 2103 2365 2106
rect 2334 2033 2341 2036
rect 2322 2013 2333 2016
rect 2322 1966 2325 2006
rect 2314 1963 2325 1966
rect 2314 1933 2317 1963
rect 2302 1913 2309 1916
rect 2266 1856 2269 1913
rect 2306 1893 2309 1913
rect 2322 1876 2325 1956
rect 2330 1903 2333 1976
rect 2314 1873 2325 1876
rect 2258 1853 2269 1856
rect 2242 1743 2245 1826
rect 2258 1756 2261 1853
rect 2274 1813 2277 1826
rect 2250 1753 2261 1756
rect 2230 1513 2237 1516
rect 2230 1396 2233 1513
rect 2242 1443 2245 1736
rect 2250 1546 2253 1753
rect 2258 1726 2261 1746
rect 2258 1723 2265 1726
rect 2262 1626 2265 1723
rect 2274 1673 2277 1806
rect 2282 1733 2285 1866
rect 2282 1706 2285 1726
rect 2290 1723 2293 1836
rect 2298 1733 2301 1846
rect 2306 1803 2309 1826
rect 2314 1733 2317 1873
rect 2322 1743 2325 1816
rect 2330 1793 2333 1806
rect 2306 1723 2317 1726
rect 2306 1706 2309 1723
rect 2282 1703 2309 1706
rect 2322 1663 2325 1736
rect 2262 1623 2285 1626
rect 2258 1566 2261 1616
rect 2282 1613 2285 1623
rect 2266 1603 2277 1606
rect 2290 1593 2293 1656
rect 2258 1563 2285 1566
rect 2250 1543 2257 1546
rect 2254 1416 2257 1543
rect 2250 1413 2257 1416
rect 2230 1393 2237 1396
rect 2242 1393 2245 1406
rect 2234 1373 2237 1393
rect 2242 1346 2245 1386
rect 2250 1363 2253 1413
rect 2266 1403 2269 1526
rect 2274 1506 2277 1536
rect 2282 1523 2285 1563
rect 2290 1533 2293 1546
rect 2298 1523 2301 1586
rect 2306 1576 2309 1596
rect 2322 1593 2325 1616
rect 2306 1573 2325 1576
rect 2330 1556 2333 1756
rect 2338 1743 2341 2033
rect 2346 2003 2349 2046
rect 2358 2036 2361 2103
rect 2378 2086 2381 2216
rect 2394 2206 2397 2566
rect 2402 2253 2405 2573
rect 2410 2543 2413 2566
rect 2410 2323 2413 2456
rect 2390 2203 2397 2206
rect 2402 2203 2405 2226
rect 2410 2223 2413 2306
rect 2390 2106 2393 2203
rect 2402 2133 2405 2196
rect 2390 2103 2397 2106
rect 2378 2083 2389 2086
rect 2354 2033 2361 2036
rect 2346 1803 2349 1986
rect 2354 1863 2357 2033
rect 2362 1973 2365 2016
rect 2354 1813 2357 1846
rect 2362 1786 2365 1946
rect 2370 1863 2373 2056
rect 2358 1783 2365 1786
rect 2338 1706 2341 1736
rect 2346 1723 2349 1756
rect 2358 1736 2361 1783
rect 2370 1743 2373 1776
rect 2358 1733 2365 1736
rect 2338 1703 2349 1706
rect 2346 1626 2349 1703
rect 2362 1653 2365 1733
rect 2338 1623 2349 1626
rect 2338 1573 2341 1623
rect 2346 1566 2349 1606
rect 2354 1593 2357 1606
rect 2346 1563 2357 1566
rect 2314 1553 2333 1556
rect 2274 1503 2285 1506
rect 2282 1396 2285 1503
rect 2242 1343 2253 1346
rect 2226 1273 2229 1336
rect 2250 1293 2253 1343
rect 2178 1123 2181 1156
rect 2138 1103 2157 1106
rect 2154 1076 2157 1103
rect 2154 1073 2165 1076
rect 2122 1053 2141 1056
rect 2122 1013 2125 1053
rect 2130 1013 2133 1026
rect 2102 963 2109 966
rect 2122 966 2125 1006
rect 2138 1003 2141 1053
rect 2122 963 2129 966
rect 2082 933 2093 936
rect 2082 913 2085 926
rect 2090 906 2093 933
rect 2082 903 2093 906
rect 2066 766 2069 826
rect 2050 763 2069 766
rect 2014 643 2045 646
rect 1994 623 2005 626
rect 1958 483 1965 486
rect 1958 356 1961 483
rect 1958 353 1965 356
rect 1946 333 1957 336
rect 1962 316 1965 353
rect 1954 313 1965 316
rect 1954 236 1957 313
rect 1970 263 1973 526
rect 1986 513 1989 606
rect 2002 546 2005 623
rect 2018 613 2021 636
rect 2026 613 2037 616
rect 1994 543 2005 546
rect 2018 543 2021 556
rect 1994 456 1997 543
rect 2026 526 2029 613
rect 2034 593 2037 606
rect 2002 513 2005 526
rect 2022 523 2029 526
rect 1994 453 2013 456
rect 1986 256 1989 406
rect 2010 386 2013 453
rect 2022 436 2025 523
rect 2022 433 2029 436
rect 2018 393 2021 416
rect 2010 383 2021 386
rect 2010 323 2013 346
rect 2018 333 2021 383
rect 2026 256 2029 433
rect 2034 353 2037 536
rect 2042 533 2045 643
rect 2050 633 2053 763
rect 2074 756 2077 866
rect 2082 803 2085 903
rect 2102 886 2105 963
rect 2126 886 2129 963
rect 2146 933 2149 1056
rect 2162 976 2165 1073
rect 2186 1003 2189 1126
rect 2202 1013 2205 1106
rect 2218 1103 2221 1226
rect 2234 1193 2237 1216
rect 2226 1123 2237 1126
rect 2154 973 2165 976
rect 2102 883 2109 886
rect 2090 816 2093 846
rect 2090 813 2101 816
rect 2090 793 2093 806
rect 2098 783 2101 813
rect 2106 803 2109 883
rect 2122 883 2129 886
rect 2114 813 2117 836
rect 2122 816 2125 883
rect 2122 813 2133 816
rect 2058 723 2061 756
rect 2066 753 2077 756
rect 2122 753 2125 806
rect 2050 416 2053 606
rect 2058 523 2061 586
rect 2066 486 2069 753
rect 2082 686 2085 736
rect 2122 723 2125 746
rect 2082 683 2105 686
rect 2102 606 2105 683
rect 2114 613 2117 636
rect 2102 603 2109 606
rect 2130 603 2133 813
rect 2138 793 2141 926
rect 2154 856 2157 973
rect 2194 946 2197 1006
rect 2210 993 2213 1006
rect 2218 983 2221 1066
rect 2234 1046 2237 1066
rect 2230 1043 2237 1046
rect 2230 976 2233 1043
rect 2242 1003 2245 1176
rect 2230 973 2237 976
rect 2194 943 2205 946
rect 2170 863 2173 936
rect 2202 896 2205 943
rect 2218 923 2221 946
rect 2194 893 2205 896
rect 2194 876 2197 893
rect 2234 886 2237 973
rect 2218 883 2237 886
rect 2190 873 2197 876
rect 2154 853 2181 856
rect 2154 773 2157 806
rect 2170 776 2173 796
rect 2162 773 2173 776
rect 2162 756 2165 773
rect 2178 766 2181 853
rect 2190 816 2193 873
rect 2190 813 2197 816
rect 2202 813 2205 876
rect 2194 793 2197 813
rect 2154 753 2165 756
rect 2170 763 2181 766
rect 2154 676 2157 753
rect 2170 686 2173 763
rect 2178 723 2181 756
rect 2170 683 2177 686
rect 2154 673 2165 676
rect 2154 613 2157 656
rect 2162 613 2165 673
rect 2174 636 2177 683
rect 2170 633 2177 636
rect 2074 493 2077 526
rect 2106 486 2109 603
rect 2170 563 2173 633
rect 2178 603 2181 616
rect 2186 603 2189 736
rect 2202 733 2205 746
rect 2194 703 2197 726
rect 2194 596 2197 616
rect 2202 603 2205 636
rect 2210 613 2213 726
rect 2218 703 2221 883
rect 2226 776 2229 846
rect 2234 796 2237 866
rect 2242 853 2245 996
rect 2250 913 2253 1246
rect 2258 986 2261 1396
rect 2274 1393 2285 1396
rect 2266 1323 2269 1366
rect 2266 1173 2269 1246
rect 2274 1166 2277 1393
rect 2290 1286 2293 1376
rect 2298 1306 2301 1486
rect 2314 1456 2317 1553
rect 2354 1546 2357 1563
rect 2362 1556 2365 1616
rect 2362 1553 2373 1556
rect 2354 1543 2365 1546
rect 2314 1453 2325 1456
rect 2322 1433 2325 1453
rect 2306 1393 2309 1416
rect 2306 1323 2309 1386
rect 2298 1303 2309 1306
rect 2266 1163 2277 1166
rect 2282 1283 2293 1286
rect 2266 1003 2269 1163
rect 2282 1156 2285 1283
rect 2290 1206 2293 1266
rect 2298 1213 2301 1296
rect 2306 1253 2309 1303
rect 2314 1213 2317 1426
rect 2330 1413 2333 1476
rect 2322 1253 2325 1406
rect 2330 1263 2333 1406
rect 2338 1256 2341 1536
rect 2346 1423 2349 1446
rect 2354 1413 2357 1426
rect 2346 1393 2349 1406
rect 2362 1386 2365 1543
rect 2370 1503 2373 1553
rect 2346 1383 2365 1386
rect 2346 1316 2349 1383
rect 2370 1376 2373 1406
rect 2378 1403 2381 2046
rect 2386 2013 2389 2083
rect 2386 1973 2389 2006
rect 2394 1933 2397 2103
rect 2402 2023 2405 2126
rect 2410 1983 2413 2206
rect 2418 2043 2421 2706
rect 2434 2703 2437 2726
rect 2442 2696 2445 2763
rect 2458 2736 2461 2856
rect 2482 2836 2485 2903
rect 2450 2733 2461 2736
rect 2466 2816 2469 2836
rect 2474 2833 2485 2836
rect 2474 2816 2477 2833
rect 2466 2813 2477 2816
rect 2458 2706 2461 2726
rect 2466 2716 2469 2813
rect 2474 2733 2477 2806
rect 2482 2753 2485 2806
rect 2490 2796 2493 2816
rect 2498 2813 2501 2876
rect 2506 2803 2509 2846
rect 2514 2813 2517 2836
rect 2522 2796 2525 2806
rect 2490 2793 2525 2796
rect 2498 2733 2501 2746
rect 2466 2713 2473 2716
rect 2450 2703 2461 2706
rect 2434 2693 2445 2696
rect 2434 2616 2437 2693
rect 2426 2613 2437 2616
rect 2426 2556 2429 2613
rect 2434 2596 2437 2606
rect 2442 2603 2445 2666
rect 2458 2636 2461 2666
rect 2470 2636 2473 2713
rect 2450 2633 2461 2636
rect 2466 2633 2473 2636
rect 2482 2636 2485 2726
rect 2482 2633 2493 2636
rect 2450 2613 2453 2633
rect 2458 2596 2461 2606
rect 2434 2593 2461 2596
rect 2426 2553 2453 2556
rect 2426 2473 2429 2536
rect 2434 2533 2437 2546
rect 2442 2466 2445 2536
rect 2450 2523 2453 2553
rect 2442 2463 2449 2466
rect 2434 2413 2437 2456
rect 2446 2406 2449 2463
rect 2426 2383 2429 2406
rect 2442 2403 2449 2406
rect 2458 2403 2461 2536
rect 2466 2513 2469 2633
rect 2474 2516 2477 2616
rect 2490 2613 2493 2633
rect 2498 2586 2501 2726
rect 2506 2623 2509 2786
rect 2538 2753 2541 2906
rect 2554 2903 2557 2926
rect 2570 2923 2589 2926
rect 2618 2923 2637 2926
rect 2642 2993 2653 2996
rect 2658 2993 2677 2996
rect 2642 2923 2645 2993
rect 2658 2983 2661 2993
rect 2658 2923 2661 2936
rect 2554 2793 2557 2806
rect 2562 2803 2565 2816
rect 2570 2776 2573 2923
rect 2602 2813 2605 2826
rect 2610 2813 2613 2846
rect 2546 2773 2573 2776
rect 2498 2583 2509 2586
rect 2482 2523 2485 2566
rect 2474 2513 2485 2516
rect 2466 2463 2469 2496
rect 2442 2376 2445 2403
rect 2426 2373 2445 2376
rect 2426 2306 2429 2373
rect 2450 2316 2453 2386
rect 2434 2313 2453 2316
rect 2426 2303 2437 2306
rect 2426 2216 2429 2276
rect 2434 2223 2437 2303
rect 2442 2283 2445 2313
rect 2458 2306 2461 2376
rect 2466 2343 2469 2416
rect 2450 2303 2461 2306
rect 2474 2303 2477 2476
rect 2490 2473 2493 2536
rect 2498 2446 2501 2576
rect 2506 2533 2509 2583
rect 2490 2443 2501 2446
rect 2490 2403 2493 2443
rect 2498 2386 2501 2416
rect 2482 2383 2501 2386
rect 2506 2383 2509 2526
rect 2482 2343 2485 2383
rect 2514 2376 2517 2656
rect 2522 2443 2525 2736
rect 2546 2693 2549 2773
rect 2594 2766 2597 2796
rect 2602 2776 2605 2806
rect 2618 2803 2621 2906
rect 2626 2813 2629 2836
rect 2634 2803 2637 2826
rect 2602 2773 2613 2776
rect 2530 2663 2541 2666
rect 2530 2603 2533 2636
rect 2530 2523 2533 2566
rect 2538 2526 2541 2663
rect 2554 2653 2557 2756
rect 2562 2706 2565 2766
rect 2594 2763 2605 2766
rect 2570 2723 2573 2756
rect 2594 2716 2597 2726
rect 2602 2723 2605 2763
rect 2610 2733 2613 2773
rect 2594 2713 2605 2716
rect 2562 2703 2569 2706
rect 2566 2636 2569 2703
rect 2562 2633 2569 2636
rect 2546 2596 2549 2616
rect 2562 2603 2565 2633
rect 2570 2596 2573 2616
rect 2586 2603 2589 2686
rect 2594 2596 2597 2696
rect 2546 2593 2597 2596
rect 2546 2563 2549 2593
rect 2546 2533 2557 2536
rect 2586 2533 2589 2556
rect 2602 2526 2605 2713
rect 2610 2703 2613 2726
rect 2610 2533 2613 2606
rect 2538 2523 2597 2526
rect 2602 2523 2613 2526
rect 2594 2506 2597 2523
rect 2586 2503 2597 2506
rect 2490 2373 2517 2376
rect 2490 2336 2493 2373
rect 2522 2366 2525 2396
rect 2530 2393 2533 2436
rect 2538 2423 2541 2466
rect 2538 2376 2541 2416
rect 2482 2333 2493 2336
rect 2506 2363 2525 2366
rect 2530 2373 2541 2376
rect 2506 2333 2509 2363
rect 2514 2326 2517 2346
rect 2490 2323 2517 2326
rect 2530 2323 2533 2373
rect 2546 2356 2549 2486
rect 2586 2436 2589 2503
rect 2586 2433 2597 2436
rect 2562 2416 2565 2426
rect 2562 2413 2581 2416
rect 2594 2413 2597 2433
rect 2554 2403 2565 2406
rect 2546 2353 2557 2356
rect 2450 2286 2453 2303
rect 2490 2296 2493 2323
rect 2458 2293 2493 2296
rect 2450 2283 2461 2286
rect 2426 2213 2433 2216
rect 2430 2156 2433 2213
rect 2442 2156 2445 2216
rect 2450 2163 2453 2216
rect 2430 2153 2437 2156
rect 2442 2153 2453 2156
rect 2418 2013 2421 2026
rect 2426 2013 2429 2136
rect 2434 2133 2437 2153
rect 2434 2016 2437 2126
rect 2442 2023 2445 2116
rect 2434 2013 2445 2016
rect 2450 2013 2453 2153
rect 2386 1813 2389 1926
rect 2394 1903 2397 1926
rect 2386 1773 2389 1796
rect 2394 1783 2397 1886
rect 2402 1873 2405 1936
rect 2410 1856 2413 1946
rect 2418 1943 2421 1956
rect 2426 1936 2429 1976
rect 2406 1853 2413 1856
rect 2422 1933 2429 1936
rect 2406 1806 2409 1853
rect 2422 1846 2425 1933
rect 2434 1883 2437 2006
rect 2418 1843 2425 1846
rect 2418 1813 2421 1843
rect 2442 1826 2445 2013
rect 2450 1926 2453 2006
rect 2458 1933 2461 2283
rect 2466 2083 2469 2206
rect 2474 2076 2477 2286
rect 2538 2263 2541 2336
rect 2546 2323 2549 2346
rect 2554 2256 2557 2353
rect 2562 2333 2565 2386
rect 2570 2323 2573 2346
rect 2578 2306 2581 2413
rect 2602 2343 2605 2486
rect 2610 2423 2613 2523
rect 2610 2403 2613 2416
rect 2586 2333 2605 2336
rect 2610 2333 2613 2366
rect 2618 2326 2621 2796
rect 2642 2766 2645 2866
rect 2626 2763 2645 2766
rect 2626 2716 2629 2763
rect 2634 2733 2637 2756
rect 2650 2733 2653 2806
rect 2658 2803 2661 2916
rect 2666 2726 2669 2836
rect 2682 2823 2693 2826
rect 2682 2813 2685 2823
rect 2674 2773 2677 2806
rect 2690 2783 2693 2816
rect 2698 2803 2701 2926
rect 2706 2813 2709 2836
rect 2682 2733 2685 2756
rect 2642 2723 2669 2726
rect 2706 2723 2709 2806
rect 2714 2803 2717 2826
rect 2722 2786 2725 2966
rect 2730 2896 2733 3036
rect 2738 2986 2741 3036
rect 2746 3023 2749 3053
rect 2754 3033 2757 3086
rect 2766 3066 2769 3123
rect 2766 3063 2773 3066
rect 2754 3013 2757 3026
rect 2762 3013 2765 3046
rect 2738 2983 2757 2986
rect 2738 2913 2741 2976
rect 2754 2973 2757 2983
rect 2770 2913 2773 3063
rect 2778 3023 2781 3133
rect 2786 3043 2789 3136
rect 2794 3123 2797 3136
rect 2802 3083 2805 3136
rect 2810 3133 2813 3336
rect 2818 3333 2829 3336
rect 2818 3203 2821 3333
rect 2826 3243 2829 3326
rect 2834 3283 2837 3343
rect 2842 3313 2845 3336
rect 2850 3333 2853 3366
rect 2858 3323 2861 3523
rect 2890 3496 2893 3526
rect 2866 3493 2893 3496
rect 2866 3403 2869 3416
rect 2874 3343 2877 3406
rect 2882 3323 2885 3426
rect 2890 3413 2893 3426
rect 2898 3406 2901 3536
rect 2906 3503 2909 3573
rect 2914 3483 2917 3636
rect 2922 3633 2933 3636
rect 2922 3623 2925 3633
rect 2938 3626 2941 3703
rect 2946 3633 2949 3713
rect 2962 3713 2981 3716
rect 2986 3743 2997 3746
rect 2938 3623 2957 3626
rect 2930 3613 2949 3616
rect 2930 3603 2933 3613
rect 2954 3603 2957 3623
rect 2922 3556 2925 3586
rect 2930 3566 2933 3596
rect 2930 3563 2949 3566
rect 2922 3553 2933 3556
rect 2922 3463 2925 3526
rect 2930 3506 2933 3553
rect 2938 3523 2941 3556
rect 2930 3503 2937 3506
rect 2934 3436 2937 3503
rect 2906 3413 2909 3436
rect 2930 3433 2937 3436
rect 2914 3413 2925 3416
rect 2890 3396 2893 3406
rect 2898 3403 2909 3406
rect 2890 3393 2901 3396
rect 2890 3333 2893 3386
rect 2842 3266 2845 3296
rect 2834 3263 2845 3266
rect 2834 3226 2837 3263
rect 2842 3236 2845 3256
rect 2858 3253 2861 3316
rect 2842 3233 2861 3236
rect 2826 3186 2829 3226
rect 2834 3223 2853 3226
rect 2850 3203 2853 3223
rect 2822 3183 2829 3186
rect 2810 3093 2813 3126
rect 2822 3086 2825 3183
rect 2822 3083 2829 3086
rect 2826 3063 2829 3083
rect 2818 3013 2821 3026
rect 2834 3006 2837 3196
rect 2842 3123 2845 3186
rect 2850 3133 2853 3176
rect 2858 3123 2861 3226
rect 2842 3023 2845 3096
rect 2850 3033 2853 3066
rect 2858 3023 2861 3046
rect 2866 3023 2869 3316
rect 2898 3266 2901 3393
rect 2906 3323 2909 3403
rect 2914 3373 2917 3413
rect 2922 3336 2925 3406
rect 2930 3343 2933 3433
rect 2946 3416 2949 3563
rect 2954 3523 2957 3556
rect 2962 3533 2965 3713
rect 2970 3613 2973 3666
rect 2978 3606 2981 3636
rect 2970 3603 2981 3606
rect 2970 3573 2973 3603
rect 2970 3523 2973 3536
rect 2954 3506 2957 3516
rect 2978 3506 2981 3526
rect 2954 3503 2981 3506
rect 2986 3486 2989 3743
rect 2994 3693 2997 3726
rect 2994 3623 2997 3656
rect 3002 3636 3005 3846
rect 3018 3843 3021 3936
rect 3026 3863 3029 3973
rect 3034 3906 3037 3966
rect 3042 3933 3045 3973
rect 3050 3953 3053 4013
rect 3066 4003 3069 4046
rect 3074 4003 3077 4086
rect 3106 4046 3109 4126
rect 3150 4086 3153 4153
rect 3082 4003 3085 4046
rect 3102 4043 3109 4046
rect 3146 4083 3153 4086
rect 3050 3923 3053 3936
rect 3058 3916 3061 3986
rect 3090 3956 3093 4016
rect 3102 3956 3105 4043
rect 3122 3983 3125 4016
rect 3074 3953 3093 3956
rect 3074 3933 3077 3953
rect 3082 3933 3085 3946
rect 3090 3933 3093 3953
rect 3098 3953 3105 3956
rect 3098 3933 3101 3953
rect 3050 3913 3061 3916
rect 3034 3903 3041 3906
rect 3038 3846 3041 3903
rect 3050 3856 3053 3913
rect 3066 3893 3069 3926
rect 3090 3916 3093 3926
rect 3106 3923 3109 3936
rect 3114 3926 3117 3936
rect 3122 3933 3133 3936
rect 3114 3923 3125 3926
rect 3130 3916 3133 3933
rect 3090 3913 3133 3916
rect 3050 3853 3057 3856
rect 3038 3843 3045 3846
rect 3018 3793 3021 3806
rect 3042 3783 3045 3843
rect 3054 3766 3057 3853
rect 3066 3813 3069 3826
rect 3090 3806 3093 3913
rect 3138 3876 3141 3946
rect 3098 3813 3101 3846
rect 3090 3803 3101 3806
rect 3050 3763 3057 3766
rect 3018 3743 3045 3746
rect 3018 3726 3021 3736
rect 3018 3723 3037 3726
rect 3010 3703 3013 3716
rect 3002 3633 3037 3636
rect 2994 3603 2997 3616
rect 3002 3613 3005 3626
rect 3026 3616 3029 3626
rect 3018 3613 3029 3616
rect 3002 3583 3005 3606
rect 3010 3576 3013 3606
rect 2994 3533 2997 3576
rect 3002 3573 3013 3576
rect 3002 3533 3005 3573
rect 3010 3526 3013 3536
rect 2954 3423 2957 3436
rect 2938 3353 2941 3416
rect 2946 3413 2957 3416
rect 2954 3403 2957 3413
rect 2962 3403 2965 3486
rect 2978 3483 2989 3486
rect 2978 3436 2981 3483
rect 2994 3473 2997 3526
rect 3002 3523 3013 3526
rect 3018 3523 3021 3613
rect 3034 3606 3037 3633
rect 3026 3603 3037 3606
rect 3042 3603 3045 3743
rect 3050 3733 3053 3763
rect 3058 3733 3061 3746
rect 3050 3683 3053 3726
rect 3066 3663 3069 3776
rect 3074 3743 3093 3746
rect 3074 3696 3077 3743
rect 3098 3733 3101 3803
rect 3106 3736 3109 3876
rect 3114 3873 3141 3876
rect 3114 3803 3117 3873
rect 3122 3796 3125 3816
rect 3130 3803 3133 3826
rect 3138 3813 3141 3866
rect 3146 3843 3149 4083
rect 3154 3943 3157 4066
rect 3162 4043 3165 4296
rect 3170 4213 3181 4216
rect 3194 4203 3197 4286
rect 3250 4256 3253 4323
rect 3234 4253 3253 4256
rect 3170 4133 3173 4146
rect 3186 4133 3189 4186
rect 3218 4183 3221 4216
rect 3202 4143 3221 4146
rect 3202 4133 3205 4143
rect 3178 4106 3181 4126
rect 3194 4123 3205 4126
rect 3202 4113 3205 4123
rect 3210 4106 3213 4136
rect 3218 4123 3221 4143
rect 3226 4133 3229 4146
rect 3178 4103 3213 4106
rect 3202 4086 3205 4103
rect 3218 4096 3221 4106
rect 3194 4083 3205 4086
rect 3210 4093 3221 4096
rect 3146 3813 3157 3816
rect 3146 3803 3149 3813
rect 3154 3796 3157 3806
rect 3122 3793 3157 3796
rect 3106 3733 3117 3736
rect 3090 3723 3109 3726
rect 3082 3706 3085 3716
rect 3082 3703 3093 3706
rect 3074 3693 3085 3696
rect 3026 3533 3029 3603
rect 3050 3583 3053 3606
rect 3034 3523 3037 3566
rect 3042 3476 3045 3536
rect 3034 3473 3045 3476
rect 2994 3443 3013 3446
rect 2978 3433 2989 3436
rect 2986 3403 2989 3433
rect 2994 3413 2997 3443
rect 2962 3376 2965 3396
rect 2962 3373 2997 3376
rect 2922 3333 2957 3336
rect 2970 3333 2973 3346
rect 2994 3333 2997 3373
rect 2914 3303 2917 3326
rect 2882 3263 2901 3266
rect 2874 3203 2877 3216
rect 2874 3123 2877 3196
rect 2882 3173 2885 3263
rect 2890 3213 2893 3256
rect 2906 3213 2909 3226
rect 2898 3133 2901 3206
rect 2914 3153 2917 3236
rect 2922 3203 2925 3333
rect 2946 3293 2949 3326
rect 2954 3323 2965 3326
rect 2930 3206 2933 3276
rect 2946 3233 2949 3276
rect 2954 3223 2957 3266
rect 2978 3246 2981 3326
rect 2986 3313 2997 3316
rect 3002 3313 3005 3436
rect 3010 3416 3013 3443
rect 3018 3423 3021 3456
rect 3034 3416 3037 3473
rect 3050 3463 3053 3526
rect 3058 3513 3061 3616
rect 3074 3606 3077 3626
rect 3082 3613 3085 3693
rect 3090 3653 3093 3703
rect 3114 3686 3117 3733
rect 3106 3683 3117 3686
rect 3122 3683 3125 3726
rect 3090 3613 3101 3616
rect 3106 3606 3109 3683
rect 3130 3676 3133 3746
rect 3122 3673 3133 3676
rect 3122 3636 3125 3673
rect 3114 3633 3125 3636
rect 3066 3603 3077 3606
rect 3094 3603 3109 3606
rect 3114 3603 3117 3616
rect 3122 3603 3125 3633
rect 3130 3606 3133 3636
rect 3138 3613 3141 3793
rect 3146 3733 3149 3786
rect 3154 3733 3157 3756
rect 3162 3736 3165 3956
rect 3170 3933 3173 4016
rect 3194 3976 3197 4083
rect 3194 3973 3205 3976
rect 3178 3923 3181 3936
rect 3186 3926 3189 3936
rect 3194 3933 3197 3956
rect 3202 3936 3205 3973
rect 3210 3953 3213 4093
rect 3226 4086 3229 4126
rect 3234 4103 3237 4253
rect 3242 4133 3245 4186
rect 3266 4166 3269 4216
rect 3274 4176 3277 4323
rect 3290 4193 3293 4206
rect 3314 4183 3317 4216
rect 3274 4173 3309 4176
rect 3266 4163 3285 4166
rect 3258 4133 3277 4136
rect 3282 4133 3285 4163
rect 3226 4083 3237 4086
rect 3202 3933 3209 3936
rect 3186 3923 3197 3926
rect 3170 3753 3173 3826
rect 3178 3813 3181 3886
rect 3186 3796 3189 3916
rect 3194 3803 3197 3876
rect 3206 3856 3209 3933
rect 3218 3863 3221 3986
rect 3226 3946 3229 4083
rect 3250 4076 3253 4126
rect 3266 4083 3269 4126
rect 3274 4123 3277 4133
rect 3282 4076 3285 4126
rect 3298 4083 3301 4166
rect 3306 4136 3309 4173
rect 3306 4133 3325 4136
rect 3306 4113 3309 4126
rect 3250 4073 3285 4076
rect 3266 4056 3269 4073
rect 3330 4063 3333 4306
rect 3370 4216 3373 4326
rect 3394 4276 3397 4296
rect 3362 4213 3373 4216
rect 3386 4273 3397 4276
rect 3386 4193 3389 4273
rect 3434 4266 3437 4340
rect 3458 4283 3461 4340
rect 3434 4263 3445 4266
rect 3338 4133 3349 4136
rect 3346 4083 3349 4126
rect 3354 4103 3357 4136
rect 3362 4056 3365 4146
rect 3378 4136 3381 4186
rect 3410 4176 3413 4216
rect 3394 4173 3413 4176
rect 3370 4133 3381 4136
rect 3370 4123 3373 4133
rect 3378 4116 3381 4126
rect 3386 4123 3389 4146
rect 3394 4133 3397 4173
rect 3394 4123 3405 4126
rect 3410 4116 3413 4136
rect 3378 4113 3413 4116
rect 3418 4113 3421 4136
rect 3426 4123 3429 4216
rect 3434 4116 3437 4263
rect 3466 4196 3469 4236
rect 3474 4206 3477 4340
rect 3490 4296 3493 4340
rect 3506 4323 3509 4340
rect 3490 4293 3541 4296
rect 3490 4263 3509 4266
rect 3490 4213 3493 4263
rect 3498 4213 3501 4256
rect 3506 4213 3509 4263
rect 3474 4203 3493 4206
rect 3506 4196 3509 4206
rect 3466 4193 3509 4196
rect 3514 4196 3517 4216
rect 3522 4203 3525 4266
rect 3538 4213 3541 4293
rect 3514 4193 3525 4196
rect 3426 4113 3437 4116
rect 3266 4053 3277 4056
rect 3242 3983 3245 4006
rect 3274 3996 3277 4053
rect 3338 4053 3365 4056
rect 3338 4036 3341 4053
rect 3334 4033 3341 4036
rect 3418 4033 3421 4106
rect 3266 3993 3277 3996
rect 3226 3943 3253 3946
rect 3226 3933 3245 3936
rect 3226 3923 3229 3933
rect 3234 3893 3237 3916
rect 3206 3853 3213 3856
rect 3162 3733 3169 3736
rect 3146 3703 3149 3716
rect 3154 3693 3157 3726
rect 3166 3686 3169 3733
rect 3178 3726 3181 3796
rect 3186 3793 3197 3796
rect 3186 3733 3189 3756
rect 3194 3733 3197 3793
rect 3202 3783 3205 3816
rect 3210 3803 3213 3853
rect 3242 3836 3245 3926
rect 3250 3873 3253 3943
rect 3266 3933 3269 3993
rect 3290 3976 3293 4016
rect 3314 4013 3325 4016
rect 3334 3986 3337 4033
rect 3334 3983 3341 3986
rect 3354 3983 3357 4006
rect 3274 3933 3277 3966
rect 3282 3946 3285 3976
rect 3290 3973 3309 3976
rect 3282 3943 3293 3946
rect 3258 3893 3261 3926
rect 3266 3923 3277 3926
rect 3266 3873 3269 3923
rect 3282 3916 3285 3936
rect 3278 3913 3285 3916
rect 3234 3833 3245 3836
rect 3226 3813 3229 3826
rect 3234 3813 3237 3833
rect 3250 3803 3253 3866
rect 3278 3796 3281 3913
rect 3210 3793 3237 3796
rect 3210 3783 3221 3786
rect 3178 3723 3197 3726
rect 3178 3703 3181 3716
rect 3186 3696 3189 3716
rect 3162 3683 3169 3686
rect 3178 3693 3189 3696
rect 3146 3623 3149 3656
rect 3162 3633 3165 3683
rect 3154 3613 3173 3616
rect 3178 3613 3181 3693
rect 3130 3603 3157 3606
rect 3162 3603 3173 3606
rect 3066 3523 3069 3603
rect 3074 3496 3077 3576
rect 3082 3533 3085 3596
rect 3094 3546 3097 3603
rect 3090 3543 3097 3546
rect 3082 3503 3085 3526
rect 3090 3496 3093 3543
rect 3066 3493 3077 3496
rect 3082 3493 3093 3496
rect 3066 3426 3069 3493
rect 3010 3413 3021 3416
rect 3018 3403 3021 3413
rect 3026 3413 3037 3416
rect 3042 3423 3069 3426
rect 3026 3403 3029 3413
rect 3034 3363 3037 3406
rect 3018 3316 3021 3346
rect 3042 3333 3045 3423
rect 3050 3413 3061 3416
rect 3066 3413 3069 3423
rect 3058 3383 3061 3406
rect 3066 3393 3069 3406
rect 3050 3343 3069 3346
rect 3074 3343 3077 3416
rect 3050 3333 3053 3343
rect 3026 3323 3053 3326
rect 2986 3293 2989 3313
rect 2994 3303 3005 3306
rect 2978 3243 2985 3246
rect 2938 3213 2965 3216
rect 2930 3203 2949 3206
rect 2930 3173 2941 3176
rect 2946 3173 2949 3203
rect 2970 3193 2973 3236
rect 2982 3186 2985 3243
rect 2994 3216 2997 3303
rect 3002 3233 3005 3256
rect 3010 3226 3013 3316
rect 3018 3313 3045 3316
rect 3050 3313 3053 3323
rect 3058 3306 3061 3336
rect 3034 3303 3061 3306
rect 3002 3223 3013 3226
rect 3018 3223 3021 3286
rect 3034 3226 3037 3303
rect 3066 3233 3069 3343
rect 3082 3333 3085 3493
rect 3090 3406 3093 3486
rect 3098 3463 3101 3526
rect 3098 3413 3101 3426
rect 3090 3403 3101 3406
rect 3106 3386 3109 3536
rect 3114 3523 3117 3586
rect 3130 3536 3133 3596
rect 3154 3593 3181 3596
rect 3122 3533 3133 3536
rect 3138 3543 3149 3546
rect 3122 3506 3125 3533
rect 3114 3503 3125 3506
rect 3130 3503 3133 3526
rect 3138 3506 3141 3543
rect 3154 3526 3157 3536
rect 3162 3533 3165 3576
rect 3146 3513 3149 3526
rect 3154 3523 3165 3526
rect 3170 3513 3173 3586
rect 3178 3516 3181 3593
rect 3186 3583 3189 3616
rect 3194 3573 3197 3723
rect 3202 3623 3205 3706
rect 3202 3603 3205 3616
rect 3210 3613 3213 3783
rect 3234 3736 3237 3793
rect 3274 3793 3281 3796
rect 3218 3733 3229 3736
rect 3234 3733 3245 3736
rect 3218 3703 3221 3716
rect 3226 3713 3229 3726
rect 3234 3693 3237 3726
rect 3222 3613 3229 3616
rect 3186 3523 3189 3536
rect 3202 3533 3205 3596
rect 3210 3573 3213 3596
rect 3210 3533 3213 3546
rect 3178 3513 3185 3516
rect 3138 3503 3165 3506
rect 3114 3483 3117 3503
rect 3098 3383 3109 3386
rect 3082 3233 3085 3326
rect 3098 3316 3101 3383
rect 3114 3363 3117 3406
rect 3122 3343 3125 3496
rect 3130 3343 3133 3416
rect 3138 3383 3141 3416
rect 3098 3313 3109 3316
rect 3034 3223 3045 3226
rect 3090 3223 3093 3296
rect 3106 3283 3109 3313
rect 3098 3233 3101 3276
rect 3114 3263 3117 3336
rect 3122 3313 3125 3336
rect 3122 3256 3125 3286
rect 3130 3273 3133 3306
rect 3106 3223 3109 3256
rect 3114 3253 3125 3256
rect 3010 3216 3013 3223
rect 2994 3213 3005 3216
rect 3010 3213 3029 3216
rect 2978 3183 2985 3186
rect 2874 3113 2885 3116
rect 2874 3016 2877 3113
rect 2882 3093 2885 3106
rect 2914 3083 2917 3126
rect 2938 3123 2941 3173
rect 2978 3166 2981 3183
rect 2946 3163 2981 3166
rect 2946 3116 2949 3163
rect 3026 3143 3029 3206
rect 3042 3193 3045 3223
rect 3058 3213 3109 3216
rect 2954 3133 3005 3136
rect 2890 3036 2893 3066
rect 2890 3033 2901 3036
rect 2842 3013 2877 3016
rect 2898 3013 2901 3026
rect 2914 3006 2917 3026
rect 2922 3013 2925 3106
rect 2930 3093 2933 3116
rect 2938 3113 2949 3116
rect 2938 3053 2941 3113
rect 2970 3056 2973 3116
rect 2946 3053 2981 3056
rect 2778 2993 2789 2996
rect 2794 2973 2797 3006
rect 2834 3003 2869 3006
rect 2874 3003 2917 3006
rect 2922 2996 2925 3006
rect 2898 2993 2925 2996
rect 2866 2966 2869 2986
rect 2862 2963 2869 2966
rect 2946 2966 2949 3053
rect 2954 3006 2957 3016
rect 2962 3013 2965 3046
rect 2970 3006 2973 3036
rect 2978 3013 2981 3053
rect 2986 3013 2989 3126
rect 3002 3113 3005 3133
rect 3058 3133 3101 3136
rect 2994 3056 2997 3106
rect 2994 3053 3005 3056
rect 2994 3006 2997 3036
rect 2954 3003 2965 3006
rect 2970 3003 2997 3006
rect 3002 3006 3005 3053
rect 3010 3013 3013 3116
rect 3018 3006 3021 3106
rect 3034 3093 3037 3126
rect 3058 3113 3061 3133
rect 3042 3103 3061 3106
rect 3026 3023 3029 3086
rect 3034 3013 3037 3026
rect 3042 3013 3045 3103
rect 3074 3093 3077 3126
rect 3106 3113 3109 3196
rect 3114 3173 3117 3253
rect 3122 3166 3125 3226
rect 3130 3223 3133 3256
rect 3138 3233 3141 3326
rect 3146 3216 3149 3486
rect 3154 3393 3157 3406
rect 3154 3313 3157 3386
rect 3162 3376 3165 3503
rect 3182 3446 3185 3513
rect 3194 3473 3197 3526
rect 3202 3466 3205 3526
rect 3194 3463 3205 3466
rect 3182 3443 3189 3446
rect 3170 3423 3181 3426
rect 3170 3386 3173 3423
rect 3178 3396 3181 3416
rect 3186 3403 3189 3443
rect 3178 3393 3189 3396
rect 3170 3383 3181 3386
rect 3162 3373 3173 3376
rect 3162 3333 3165 3366
rect 3142 3213 3149 3216
rect 3114 3163 3125 3166
rect 3050 3033 3061 3036
rect 3066 3023 3069 3056
rect 3082 3013 3085 3106
rect 3114 3033 3117 3163
rect 3130 3156 3133 3176
rect 3122 3153 3133 3156
rect 3122 3123 3125 3153
rect 3142 3146 3145 3213
rect 3142 3143 3149 3146
rect 3154 3143 3157 3276
rect 3130 3106 3133 3136
rect 3122 3103 3133 3106
rect 3138 3103 3141 3126
rect 3146 3073 3149 3143
rect 3154 3053 3157 3136
rect 3162 3123 3165 3326
rect 3170 3293 3173 3373
rect 3178 3343 3181 3383
rect 3186 3346 3189 3393
rect 3194 3356 3197 3463
rect 3210 3456 3213 3526
rect 3218 3503 3221 3586
rect 3226 3523 3229 3606
rect 3234 3526 3237 3646
rect 3242 3533 3245 3733
rect 3250 3703 3253 3716
rect 3258 3693 3261 3716
rect 3266 3643 3269 3746
rect 3274 3733 3277 3793
rect 3290 3783 3293 3943
rect 3306 3933 3309 3973
rect 3338 3946 3341 3983
rect 3338 3943 3349 3946
rect 3322 3926 3325 3936
rect 3330 3933 3341 3936
rect 3314 3913 3317 3926
rect 3322 3923 3333 3926
rect 3346 3916 3349 3943
rect 3322 3913 3349 3916
rect 3322 3826 3325 3913
rect 3354 3896 3357 3966
rect 3318 3823 3325 3826
rect 3346 3893 3357 3896
rect 3298 3803 3301 3816
rect 3318 3766 3321 3823
rect 3330 3793 3333 3816
rect 3338 3796 3341 3816
rect 3346 3803 3349 3893
rect 3370 3836 3373 3956
rect 3378 3933 3381 4016
rect 3426 4013 3429 4113
rect 3434 4006 3437 4086
rect 3418 4003 3437 4006
rect 3394 3926 3397 3936
rect 3402 3933 3405 3956
rect 3418 3933 3421 4003
rect 3442 3966 3445 4126
rect 3450 4113 3453 4136
rect 3450 4003 3453 4016
rect 3458 4003 3461 4126
rect 3466 4103 3469 4136
rect 3474 4123 3477 4146
rect 3482 4106 3485 4186
rect 3498 4133 3501 4186
rect 3514 4163 3517 4193
rect 3538 4176 3541 4206
rect 3562 4183 3565 4216
rect 3570 4176 3573 4296
rect 3586 4256 3589 4340
rect 3586 4253 3621 4256
rect 3586 4216 3589 4253
rect 3538 4173 3573 4176
rect 3570 4163 3573 4173
rect 3582 4213 3589 4216
rect 3582 4156 3585 4213
rect 3610 4206 3613 4216
rect 3618 4213 3621 4253
rect 3610 4203 3621 4206
rect 3634 4203 3637 4296
rect 3650 4246 3653 4340
rect 3714 4337 3749 4340
rect 3650 4243 3661 4246
rect 3578 4153 3585 4156
rect 3514 4133 3517 4146
rect 3478 4103 3485 4106
rect 3478 4026 3481 4103
rect 3478 4023 3485 4026
rect 3434 3963 3445 3966
rect 3386 3916 3389 3926
rect 3394 3923 3405 3926
rect 3410 3923 3421 3926
rect 3410 3916 3413 3923
rect 3386 3913 3413 3916
rect 3418 3863 3421 3923
rect 3370 3833 3413 3836
rect 3370 3823 3397 3826
rect 3370 3813 3373 3823
rect 3394 3816 3397 3823
rect 3378 3813 3389 3816
rect 3394 3813 3405 3816
rect 3354 3803 3365 3806
rect 3378 3803 3381 3813
rect 3410 3806 3413 3833
rect 3386 3796 3389 3806
rect 3338 3793 3389 3796
rect 3318 3763 3325 3766
rect 3282 3743 3285 3756
rect 3282 3693 3285 3736
rect 3290 3643 3293 3746
rect 3306 3713 3309 3726
rect 3314 3636 3317 3746
rect 3322 3733 3325 3763
rect 3330 3723 3333 3786
rect 3338 3783 3349 3786
rect 3338 3733 3341 3783
rect 3386 3776 3389 3793
rect 3402 3803 3413 3806
rect 3338 3703 3341 3726
rect 3346 3656 3349 3746
rect 3354 3703 3357 3776
rect 3386 3773 3393 3776
rect 3370 3733 3373 3756
rect 3330 3653 3349 3656
rect 3306 3633 3317 3636
rect 3250 3596 3253 3616
rect 3266 3603 3269 3616
rect 3250 3593 3269 3596
rect 3234 3523 3245 3526
rect 3242 3476 3245 3516
rect 3234 3473 3245 3476
rect 3250 3473 3253 3576
rect 3266 3556 3269 3593
rect 3274 3583 3277 3606
rect 3258 3553 3269 3556
rect 3282 3556 3285 3616
rect 3290 3603 3293 3616
rect 3298 3576 3301 3616
rect 3290 3573 3301 3576
rect 3306 3573 3309 3633
rect 3314 3603 3317 3626
rect 3322 3603 3325 3646
rect 3330 3596 3333 3653
rect 3338 3603 3341 3646
rect 3346 3633 3365 3636
rect 3346 3613 3349 3633
rect 3346 3596 3349 3606
rect 3354 3603 3357 3626
rect 3362 3616 3365 3633
rect 3370 3623 3373 3716
rect 3362 3613 3373 3616
rect 3370 3603 3373 3613
rect 3322 3584 3325 3596
rect 3330 3593 3349 3596
rect 3316 3581 3325 3584
rect 3316 3566 3319 3581
rect 3330 3566 3333 3576
rect 3282 3553 3293 3556
rect 3258 3466 3261 3553
rect 3266 3543 3277 3546
rect 3266 3533 3269 3543
rect 3274 3533 3285 3536
rect 3266 3516 3269 3526
rect 3274 3523 3285 3526
rect 3266 3513 3277 3516
rect 3258 3463 3269 3466
rect 3210 3453 3245 3456
rect 3202 3366 3205 3406
rect 3210 3403 3213 3416
rect 3218 3376 3221 3416
rect 3226 3413 3229 3446
rect 3226 3393 3229 3406
rect 3218 3373 3229 3376
rect 3202 3363 3221 3366
rect 3194 3353 3213 3356
rect 3186 3343 3197 3346
rect 3170 3143 3173 3236
rect 3178 3223 3181 3336
rect 3194 3333 3197 3343
rect 3186 3313 3189 3326
rect 3202 3306 3205 3326
rect 3198 3303 3205 3306
rect 3186 3216 3189 3236
rect 3198 3216 3201 3303
rect 3178 3213 3189 3216
rect 3194 3213 3201 3216
rect 3170 3083 3173 3136
rect 3002 3003 3021 3006
rect 2962 2996 2965 3003
rect 3002 2996 3005 3003
rect 2962 2993 3005 2996
rect 2946 2963 2953 2966
rect 2730 2893 2737 2896
rect 2734 2816 2737 2893
rect 2730 2813 2737 2816
rect 2730 2793 2733 2813
rect 2746 2803 2749 2906
rect 2762 2853 2797 2856
rect 2754 2786 2757 2846
rect 2762 2813 2765 2853
rect 2714 2783 2725 2786
rect 2750 2783 2757 2786
rect 2626 2713 2645 2716
rect 2642 2696 2645 2713
rect 2626 2603 2629 2626
rect 2634 2613 2637 2696
rect 2642 2693 2653 2696
rect 2650 2636 2653 2693
rect 2674 2686 2677 2706
rect 2642 2633 2653 2636
rect 2666 2683 2677 2686
rect 2666 2636 2669 2683
rect 2666 2633 2677 2636
rect 2634 2596 2637 2606
rect 2626 2593 2637 2596
rect 2626 2533 2629 2593
rect 2634 2533 2637 2546
rect 2626 2403 2629 2516
rect 2634 2473 2637 2526
rect 2642 2513 2645 2633
rect 2650 2583 2653 2606
rect 2666 2596 2669 2616
rect 2674 2603 2677 2633
rect 2682 2603 2685 2696
rect 2690 2596 2693 2616
rect 2666 2593 2693 2596
rect 2650 2506 2653 2566
rect 2642 2503 2653 2506
rect 2626 2363 2629 2396
rect 2634 2346 2637 2386
rect 2574 2303 2581 2306
rect 2586 2323 2621 2326
rect 2630 2343 2637 2346
rect 2530 2253 2557 2256
rect 2490 2136 2493 2206
rect 2482 2093 2485 2136
rect 2490 2133 2501 2136
rect 2466 2073 2477 2076
rect 2466 1943 2469 2073
rect 2490 2056 2493 2126
rect 2498 2063 2501 2133
rect 2514 2056 2517 2166
rect 2522 2096 2525 2246
rect 2530 2113 2533 2253
rect 2538 2213 2541 2226
rect 2562 2203 2565 2266
rect 2574 2236 2577 2303
rect 2574 2233 2581 2236
rect 2570 2146 2573 2216
rect 2538 2143 2573 2146
rect 2538 2133 2541 2143
rect 2562 2126 2565 2136
rect 2550 2123 2565 2126
rect 2522 2093 2529 2096
rect 2482 2053 2493 2056
rect 2498 2053 2517 2056
rect 2482 2013 2485 2053
rect 2474 1946 2477 2006
rect 2490 1953 2493 2046
rect 2498 1946 2501 2053
rect 2506 1953 2509 2026
rect 2514 1993 2517 2046
rect 2526 2026 2529 2093
rect 2522 2023 2529 2026
rect 2474 1943 2501 1946
rect 2450 1923 2457 1926
rect 2466 1923 2469 1936
rect 2426 1823 2445 1826
rect 2454 1826 2457 1923
rect 2454 1823 2461 1826
rect 2406 1803 2413 1806
rect 2386 1713 2389 1726
rect 2394 1613 2397 1746
rect 2410 1733 2413 1803
rect 2426 1736 2429 1823
rect 2434 1746 2437 1806
rect 2442 1803 2445 1816
rect 2458 1806 2461 1823
rect 2466 1813 2469 1886
rect 2434 1743 2445 1746
rect 2410 1713 2413 1726
rect 2418 1683 2421 1736
rect 2426 1733 2437 1736
rect 2426 1713 2429 1726
rect 2386 1573 2389 1596
rect 2402 1553 2405 1606
rect 2386 1406 2389 1526
rect 2402 1486 2405 1546
rect 2394 1483 2405 1486
rect 2394 1413 2397 1483
rect 2410 1426 2413 1656
rect 2418 1473 2421 1606
rect 2426 1553 2429 1616
rect 2434 1473 2437 1733
rect 2442 1543 2445 1743
rect 2450 1706 2453 1806
rect 2458 1803 2469 1806
rect 2458 1743 2461 1776
rect 2466 1723 2469 1736
rect 2450 1703 2461 1706
rect 2458 1616 2461 1703
rect 2474 1676 2477 1943
rect 2482 1916 2485 1926
rect 2482 1913 2489 1916
rect 2486 1836 2489 1913
rect 2486 1833 2493 1836
rect 2490 1813 2493 1833
rect 2490 1746 2493 1796
rect 2482 1743 2493 1746
rect 2482 1733 2485 1743
rect 2450 1613 2461 1616
rect 2470 1673 2477 1676
rect 2410 1423 2421 1426
rect 2386 1403 2405 1406
rect 2362 1373 2373 1376
rect 2354 1323 2357 1346
rect 2362 1333 2365 1373
rect 2370 1336 2373 1366
rect 2370 1333 2381 1336
rect 2394 1333 2397 1346
rect 2402 1343 2405 1386
rect 2410 1326 2413 1416
rect 2418 1383 2421 1423
rect 2442 1406 2445 1526
rect 2450 1416 2453 1613
rect 2458 1543 2461 1596
rect 2470 1536 2473 1673
rect 2482 1593 2485 1726
rect 2490 1723 2493 1736
rect 2490 1613 2493 1666
rect 2458 1533 2473 1536
rect 2458 1443 2461 1533
rect 2450 1413 2461 1416
rect 2442 1403 2453 1406
rect 2362 1316 2365 1326
rect 2386 1323 2413 1326
rect 2418 1343 2445 1346
rect 2346 1313 2365 1316
rect 2330 1253 2341 1256
rect 2290 1203 2301 1206
rect 2274 1153 2285 1156
rect 2274 1023 2277 1153
rect 2282 1123 2285 1146
rect 2290 1133 2293 1156
rect 2290 1103 2293 1126
rect 2274 993 2277 1016
rect 2298 1013 2301 1203
rect 2306 1133 2309 1196
rect 2322 1133 2325 1146
rect 2314 1123 2325 1126
rect 2330 1106 2333 1253
rect 2362 1223 2365 1313
rect 2418 1306 2421 1343
rect 2410 1303 2421 1306
rect 2326 1103 2333 1106
rect 2306 993 2309 1006
rect 2258 983 2265 986
rect 2262 906 2265 983
rect 2314 946 2317 1056
rect 2326 1036 2329 1103
rect 2326 1033 2333 1036
rect 2274 943 2317 946
rect 2274 933 2277 943
rect 2258 903 2265 906
rect 2274 903 2277 926
rect 2242 803 2245 816
rect 2234 793 2245 796
rect 2226 773 2233 776
rect 2230 696 2233 773
rect 2226 693 2233 696
rect 2242 693 2245 756
rect 2210 603 2221 606
rect 2226 596 2229 693
rect 2154 523 2157 546
rect 2066 483 2077 486
rect 2106 483 2133 486
rect 2050 413 2069 416
rect 2074 386 2077 483
rect 2098 386 2101 406
rect 2130 396 2133 483
rect 2074 383 2101 386
rect 2122 393 2133 396
rect 2146 393 2149 416
rect 2074 366 2077 383
rect 2074 363 2081 366
rect 2066 323 2069 336
rect 2078 296 2081 363
rect 1978 253 1989 256
rect 2018 253 2029 256
rect 2074 293 2081 296
rect 1954 233 1965 236
rect 1962 213 1965 233
rect 1946 203 1957 206
rect 1978 203 1981 253
rect 1938 193 1949 196
rect 2002 193 2005 216
rect 1946 133 1949 193
rect 2018 166 2021 253
rect 2058 203 2061 216
rect 2074 186 2077 293
rect 2098 266 2101 366
rect 2122 363 2125 393
rect 2146 323 2149 346
rect 2090 263 2101 266
rect 2090 203 2093 263
rect 2130 236 2133 256
rect 2126 233 2133 236
rect 2126 186 2129 233
rect 2138 193 2141 216
rect 2074 183 2093 186
rect 2126 183 2133 186
rect 2018 163 2029 166
rect 1978 123 1981 136
rect 2002 123 2005 146
rect 2026 143 2029 163
rect 2058 123 2061 156
rect 2090 123 2093 183
rect 2130 123 2133 183
rect 2178 63 2181 596
rect 2194 593 2229 596
rect 2242 593 2245 676
rect 2250 663 2253 816
rect 2258 793 2261 903
rect 2274 803 2277 856
rect 2282 836 2285 926
rect 2290 873 2293 936
rect 2298 893 2301 926
rect 2282 833 2293 836
rect 2282 786 2285 826
rect 2258 783 2285 786
rect 2194 506 2197 526
rect 2190 503 2197 506
rect 2190 436 2193 503
rect 2190 433 2197 436
rect 2194 413 2197 433
rect 2202 326 2205 556
rect 2210 503 2213 526
rect 2218 473 2221 526
rect 2226 516 2229 593
rect 2250 583 2253 606
rect 2234 523 2245 526
rect 2250 523 2253 576
rect 2242 516 2245 523
rect 2258 516 2261 783
rect 2290 776 2293 833
rect 2306 813 2309 936
rect 2314 933 2317 943
rect 2298 803 2309 806
rect 2314 803 2317 906
rect 2322 806 2325 1016
rect 2330 956 2333 1033
rect 2338 1013 2341 1176
rect 2346 1133 2349 1156
rect 2338 973 2341 996
rect 2330 953 2337 956
rect 2334 886 2337 953
rect 2330 883 2337 886
rect 2330 863 2333 883
rect 2330 813 2333 856
rect 2346 843 2349 1106
rect 2354 1063 2357 1216
rect 2370 1133 2373 1216
rect 2378 1176 2381 1266
rect 2410 1236 2413 1303
rect 2426 1253 2429 1276
rect 2410 1233 2421 1236
rect 2378 1173 2389 1176
rect 2370 1123 2381 1126
rect 2386 1116 2389 1173
rect 2362 1056 2365 1106
rect 2354 1053 2365 1056
rect 2354 996 2357 1053
rect 2370 1013 2373 1116
rect 2378 1113 2389 1116
rect 2378 1103 2381 1113
rect 2394 1106 2397 1206
rect 2386 1103 2397 1106
rect 2386 1013 2389 1103
rect 2402 1086 2405 1216
rect 2398 1083 2405 1086
rect 2398 1016 2401 1083
rect 2398 1013 2405 1016
rect 2378 1002 2389 1005
rect 2354 993 2381 996
rect 2386 993 2389 1002
rect 2402 996 2405 1013
rect 2410 1003 2413 1216
rect 2418 1086 2421 1233
rect 2426 1213 2429 1246
rect 2426 1186 2429 1206
rect 2434 1203 2437 1336
rect 2442 1303 2445 1326
rect 2450 1243 2453 1403
rect 2458 1273 2461 1413
rect 2466 1266 2469 1406
rect 2474 1343 2477 1516
rect 2458 1263 2469 1266
rect 2442 1213 2453 1216
rect 2426 1183 2433 1186
rect 2430 1106 2433 1183
rect 2442 1126 2445 1146
rect 2450 1133 2453 1196
rect 2458 1133 2461 1263
rect 2466 1213 2469 1256
rect 2482 1246 2485 1546
rect 2490 1523 2493 1606
rect 2490 1423 2493 1516
rect 2490 1353 2493 1416
rect 2498 1336 2501 1936
rect 2514 1933 2517 1946
rect 2506 1903 2509 1926
rect 2514 1886 2517 1926
rect 2510 1883 2517 1886
rect 2510 1816 2513 1883
rect 2510 1813 2517 1816
rect 2506 1743 2509 1796
rect 2514 1726 2517 1813
rect 2510 1723 2517 1726
rect 2510 1646 2513 1723
rect 2510 1643 2517 1646
rect 2506 1603 2509 1626
rect 2514 1596 2517 1643
rect 2506 1593 2517 1596
rect 2506 1533 2509 1593
rect 2506 1413 2509 1526
rect 2514 1483 2517 1576
rect 2522 1466 2525 2023
rect 2530 1923 2533 2006
rect 2538 1996 2541 2086
rect 2550 2036 2553 2123
rect 2562 2063 2565 2116
rect 2570 2113 2573 2143
rect 2570 2073 2573 2106
rect 2546 2033 2553 2036
rect 2546 2013 2549 2033
rect 2578 2026 2581 2233
rect 2586 2216 2589 2323
rect 2594 2313 2605 2316
rect 2594 2233 2597 2313
rect 2586 2213 2593 2216
rect 2590 2146 2593 2213
rect 2586 2143 2593 2146
rect 2586 2053 2589 2143
rect 2602 2133 2605 2306
rect 2630 2246 2633 2343
rect 2642 2283 2645 2503
rect 2650 2413 2653 2436
rect 2658 2406 2661 2546
rect 2666 2526 2669 2593
rect 2674 2543 2693 2546
rect 2666 2523 2677 2526
rect 2674 2446 2677 2523
rect 2690 2503 2693 2526
rect 2698 2473 2701 2656
rect 2706 2533 2709 2706
rect 2714 2563 2717 2783
rect 2722 2603 2725 2726
rect 2730 2643 2733 2726
rect 2750 2676 2753 2783
rect 2762 2773 2765 2806
rect 2770 2803 2773 2816
rect 2778 2803 2781 2836
rect 2786 2813 2789 2826
rect 2794 2803 2797 2853
rect 2810 2833 2813 2926
rect 2818 2876 2821 2896
rect 2818 2873 2825 2876
rect 2762 2713 2765 2726
rect 2738 2603 2741 2676
rect 2750 2673 2757 2676
rect 2754 2653 2757 2673
rect 2762 2556 2765 2676
rect 2714 2553 2765 2556
rect 2714 2526 2717 2553
rect 2706 2523 2717 2526
rect 2722 2523 2725 2546
rect 2730 2516 2733 2526
rect 2722 2513 2733 2516
rect 2650 2403 2661 2406
rect 2666 2443 2677 2446
rect 2650 2363 2653 2403
rect 2666 2353 2669 2443
rect 2674 2403 2677 2426
rect 2690 2403 2693 2416
rect 2658 2313 2661 2336
rect 2666 2323 2669 2346
rect 2682 2286 2685 2356
rect 2698 2346 2701 2406
rect 2698 2343 2717 2346
rect 2682 2283 2705 2286
rect 2618 2243 2633 2246
rect 2610 2193 2613 2216
rect 2618 2186 2621 2243
rect 2626 2213 2629 2236
rect 2634 2203 2637 2226
rect 2642 2223 2653 2226
rect 2642 2186 2645 2223
rect 2650 2193 2653 2206
rect 2610 2133 2613 2186
rect 2618 2183 2629 2186
rect 2642 2183 2653 2186
rect 2626 2126 2629 2183
rect 2594 2123 2605 2126
rect 2618 2123 2629 2126
rect 2578 2023 2589 2026
rect 2554 2013 2581 2016
rect 2554 2003 2557 2013
rect 2570 2003 2581 2006
rect 2538 1993 2581 1996
rect 2538 1873 2541 1993
rect 2578 1973 2581 1993
rect 2554 1856 2557 1936
rect 2578 1923 2581 1956
rect 2538 1853 2557 1856
rect 2538 1823 2541 1853
rect 2538 1783 2541 1806
rect 2562 1796 2565 1816
rect 2554 1793 2565 1796
rect 2530 1736 2533 1746
rect 2554 1743 2557 1793
rect 2530 1733 2557 1736
rect 2530 1723 2549 1726
rect 2554 1706 2557 1733
rect 2550 1703 2557 1706
rect 2538 1606 2541 1696
rect 2550 1636 2553 1703
rect 2562 1663 2565 1746
rect 2570 1693 2573 1876
rect 2586 1866 2589 2023
rect 2594 2003 2597 2123
rect 2618 2063 2621 2123
rect 2642 2066 2645 2136
rect 2650 2093 2653 2183
rect 2658 2116 2661 2136
rect 2658 2113 2665 2116
rect 2642 2063 2653 2066
rect 2602 1996 2605 2056
rect 2618 2003 2621 2036
rect 2650 2013 2653 2063
rect 2594 1993 2605 1996
rect 2594 1976 2597 1993
rect 2650 1986 2653 2006
rect 2602 1983 2621 1986
rect 2618 1976 2621 1983
rect 2634 1983 2653 1986
rect 2634 1976 2637 1983
rect 2594 1973 2605 1976
rect 2618 1973 2637 1976
rect 2594 1923 2597 1956
rect 2578 1863 2589 1866
rect 2578 1706 2581 1863
rect 2586 1793 2589 1816
rect 2602 1776 2605 1973
rect 2650 1946 2653 1966
rect 2662 1956 2665 2113
rect 2674 2063 2677 2206
rect 2702 2156 2705 2283
rect 2714 2186 2717 2343
rect 2722 2233 2725 2513
rect 2746 2496 2749 2536
rect 2762 2516 2765 2546
rect 2770 2523 2773 2786
rect 2778 2783 2797 2786
rect 2778 2643 2781 2783
rect 2786 2733 2789 2776
rect 2794 2736 2797 2783
rect 2794 2733 2805 2736
rect 2786 2713 2789 2726
rect 2794 2656 2797 2726
rect 2810 2706 2813 2826
rect 2822 2806 2825 2873
rect 2818 2803 2825 2806
rect 2818 2783 2821 2803
rect 2818 2713 2821 2736
rect 2826 2733 2829 2776
rect 2842 2746 2845 2926
rect 2850 2903 2853 2926
rect 2862 2856 2865 2963
rect 2914 2936 2917 2956
rect 2862 2853 2869 2856
rect 2834 2743 2845 2746
rect 2826 2706 2829 2726
rect 2810 2703 2829 2706
rect 2834 2683 2837 2743
rect 2842 2723 2845 2736
rect 2850 2686 2853 2776
rect 2842 2683 2853 2686
rect 2786 2653 2797 2656
rect 2778 2533 2781 2616
rect 2786 2543 2789 2653
rect 2802 2543 2805 2656
rect 2810 2623 2829 2626
rect 2786 2523 2805 2526
rect 2762 2513 2781 2516
rect 2738 2493 2749 2496
rect 2738 2403 2741 2493
rect 2746 2443 2773 2446
rect 2746 2413 2749 2443
rect 2754 2403 2757 2416
rect 2770 2413 2773 2443
rect 2778 2406 2781 2513
rect 2786 2456 2789 2476
rect 2786 2453 2793 2456
rect 2762 2366 2765 2406
rect 2730 2363 2765 2366
rect 2770 2403 2781 2406
rect 2730 2323 2733 2363
rect 2754 2323 2765 2326
rect 2722 2193 2725 2216
rect 2714 2183 2725 2186
rect 2702 2153 2709 2156
rect 2682 2133 2685 2146
rect 2690 2133 2701 2136
rect 2646 1943 2653 1946
rect 2658 1953 2665 1956
rect 2618 1886 2621 1926
rect 2634 1903 2637 1926
rect 2646 1886 2649 1943
rect 2594 1773 2605 1776
rect 2610 1883 2621 1886
rect 2638 1883 2649 1886
rect 2586 1723 2589 1736
rect 2594 1733 2597 1773
rect 2578 1703 2589 1706
rect 2550 1633 2557 1636
rect 2554 1613 2557 1633
rect 2562 1613 2565 1636
rect 2538 1603 2545 1606
rect 2530 1543 2533 1596
rect 2518 1463 2525 1466
rect 2518 1416 2521 1463
rect 2530 1423 2533 1526
rect 2542 1506 2545 1603
rect 2570 1533 2573 1656
rect 2586 1626 2589 1703
rect 2602 1693 2605 1736
rect 2578 1623 2589 1626
rect 2578 1573 2581 1623
rect 2610 1613 2613 1883
rect 2638 1826 2641 1883
rect 2658 1836 2661 1953
rect 2674 1933 2677 1956
rect 2666 1873 2669 1926
rect 2682 1906 2685 2096
rect 2698 2093 2701 2126
rect 2690 1963 2693 2076
rect 2698 1923 2701 2056
rect 2706 1953 2709 2153
rect 2714 2013 2717 2146
rect 2722 2003 2725 2183
rect 2730 2063 2733 2166
rect 2730 2013 2733 2026
rect 2738 1956 2741 2256
rect 2746 2106 2749 2276
rect 2754 2136 2757 2216
rect 2762 2213 2765 2236
rect 2770 2156 2773 2403
rect 2790 2396 2793 2453
rect 2802 2403 2805 2516
rect 2810 2403 2813 2623
rect 2818 2503 2821 2616
rect 2826 2613 2829 2623
rect 2826 2506 2829 2546
rect 2834 2513 2837 2606
rect 2826 2503 2837 2506
rect 2842 2496 2845 2683
rect 2850 2543 2853 2646
rect 2818 2493 2845 2496
rect 2786 2393 2793 2396
rect 2778 2163 2781 2206
rect 2770 2153 2781 2156
rect 2754 2133 2773 2136
rect 2778 2126 2781 2153
rect 2786 2143 2789 2393
rect 2818 2386 2821 2493
rect 2826 2483 2837 2486
rect 2826 2426 2829 2483
rect 2834 2443 2837 2476
rect 2850 2436 2853 2526
rect 2858 2516 2861 2796
rect 2866 2723 2869 2853
rect 2874 2843 2877 2886
rect 2866 2523 2869 2716
rect 2874 2593 2877 2806
rect 2882 2753 2885 2936
rect 2906 2933 2917 2936
rect 2890 2813 2893 2826
rect 2906 2776 2909 2933
rect 2930 2923 2933 2936
rect 2950 2886 2953 2963
rect 2946 2883 2953 2886
rect 2962 2883 2965 2993
rect 2914 2793 2917 2846
rect 2890 2773 2909 2776
rect 2890 2733 2893 2773
rect 2914 2686 2917 2726
rect 2922 2723 2925 2876
rect 2882 2683 2917 2686
rect 2882 2603 2885 2683
rect 2922 2643 2925 2686
rect 2930 2636 2933 2856
rect 2938 2803 2941 2876
rect 2946 2853 2949 2883
rect 2970 2866 2973 2926
rect 2946 2813 2949 2846
rect 2954 2813 2957 2866
rect 2966 2863 2973 2866
rect 2966 2806 2969 2863
rect 2978 2813 2981 2976
rect 2986 2973 3029 2976
rect 2986 2923 2989 2973
rect 2994 2933 2997 2946
rect 3002 2933 3013 2936
rect 3026 2933 3029 2973
rect 3002 2923 3013 2926
rect 3018 2913 3021 2926
rect 2954 2753 2957 2806
rect 2966 2803 2973 2806
rect 2986 2803 2989 2866
rect 3010 2823 3029 2826
rect 3002 2803 3005 2816
rect 2970 2736 2973 2803
rect 2994 2773 2997 2796
rect 3010 2786 3013 2823
rect 3002 2783 3013 2786
rect 3018 2783 3021 2816
rect 3026 2803 3029 2823
rect 3010 2756 3013 2783
rect 2970 2733 2981 2736
rect 2914 2633 2933 2636
rect 2890 2613 2909 2616
rect 2898 2586 2901 2606
rect 2890 2583 2901 2586
rect 2890 2536 2893 2583
rect 2914 2556 2917 2633
rect 2938 2626 2941 2726
rect 2954 2686 2957 2696
rect 2922 2603 2925 2626
rect 2930 2623 2941 2626
rect 2946 2683 2957 2686
rect 2858 2513 2865 2516
rect 2874 2513 2877 2536
rect 2882 2533 2893 2536
rect 2906 2553 2917 2556
rect 2882 2516 2885 2533
rect 2906 2516 2909 2553
rect 2914 2533 2917 2546
rect 2882 2513 2889 2516
rect 2906 2513 2913 2516
rect 2862 2456 2865 2513
rect 2862 2453 2869 2456
rect 2850 2433 2861 2436
rect 2826 2423 2853 2426
rect 2826 2413 2829 2423
rect 2814 2383 2821 2386
rect 2826 2403 2837 2406
rect 2842 2403 2845 2416
rect 2814 2306 2817 2383
rect 2826 2323 2829 2403
rect 2814 2303 2821 2306
rect 2818 2283 2821 2303
rect 2850 2253 2853 2423
rect 2802 2223 2829 2226
rect 2802 2213 2805 2223
rect 2794 2193 2797 2206
rect 2770 2123 2781 2126
rect 2786 2123 2797 2126
rect 2762 2106 2765 2116
rect 2746 2103 2765 2106
rect 2746 1963 2749 2103
rect 2754 2023 2757 2066
rect 2762 1983 2765 2096
rect 2730 1953 2741 1956
rect 2658 1833 2669 1836
rect 2618 1733 2621 1826
rect 2638 1823 2653 1826
rect 2626 1726 2629 1736
rect 2634 1733 2637 1806
rect 2622 1723 2629 1726
rect 2622 1636 2625 1723
rect 2634 1683 2637 1726
rect 2618 1633 2625 1636
rect 2618 1613 2621 1633
rect 2642 1616 2645 1806
rect 2650 1683 2653 1823
rect 2666 1803 2669 1833
rect 2642 1613 2649 1616
rect 2538 1503 2545 1506
rect 2554 1523 2581 1526
rect 2538 1433 2541 1503
rect 2518 1413 2525 1416
rect 2546 1413 2549 1486
rect 2554 1463 2557 1523
rect 2586 1516 2589 1606
rect 2602 1593 2605 1606
rect 2610 1583 2613 1606
rect 2578 1513 2589 1516
rect 2554 1413 2557 1436
rect 2562 1433 2573 1436
rect 2474 1243 2485 1246
rect 2494 1333 2501 1336
rect 2514 1333 2517 1366
rect 2494 1246 2497 1333
rect 2522 1326 2525 1413
rect 2538 1403 2549 1406
rect 2538 1363 2549 1366
rect 2506 1276 2509 1326
rect 2514 1323 2525 1326
rect 2514 1283 2517 1323
rect 2538 1296 2541 1336
rect 2522 1293 2541 1296
rect 2522 1276 2525 1293
rect 2506 1273 2525 1276
rect 2530 1266 2533 1286
rect 2506 1263 2533 1266
rect 2494 1243 2501 1246
rect 2474 1156 2477 1243
rect 2482 1203 2485 1216
rect 2490 1203 2493 1226
rect 2498 1193 2501 1243
rect 2470 1153 2477 1156
rect 2442 1123 2461 1126
rect 2430 1103 2437 1106
rect 2418 1083 2425 1086
rect 2422 1026 2425 1083
rect 2418 1023 2425 1026
rect 2434 1026 2437 1103
rect 2458 1046 2461 1123
rect 2470 1096 2473 1153
rect 2482 1136 2485 1146
rect 2482 1133 2501 1136
rect 2506 1133 2509 1263
rect 2514 1203 2517 1216
rect 2522 1206 2525 1256
rect 2530 1213 2533 1246
rect 2522 1203 2533 1206
rect 2482 1106 2485 1126
rect 2482 1103 2489 1106
rect 2470 1093 2477 1096
rect 2458 1043 2469 1046
rect 2434 1023 2453 1026
rect 2402 993 2413 996
rect 2354 983 2373 986
rect 2354 933 2357 946
rect 2362 893 2365 966
rect 2338 813 2349 816
rect 2322 803 2333 806
rect 2330 786 2333 803
rect 2338 793 2341 806
rect 2322 783 2333 786
rect 2362 783 2365 816
rect 2282 773 2309 776
rect 2266 723 2269 736
rect 2274 716 2277 726
rect 2282 723 2285 773
rect 2290 733 2293 756
rect 2274 713 2293 716
rect 2282 686 2285 706
rect 2274 683 2285 686
rect 2274 636 2277 683
rect 2274 633 2285 636
rect 2266 603 2269 616
rect 2274 553 2277 616
rect 2282 606 2285 633
rect 2290 613 2293 713
rect 2298 683 2301 726
rect 2306 646 2309 773
rect 2314 723 2317 736
rect 2298 643 2309 646
rect 2282 603 2293 606
rect 2226 513 2237 516
rect 2242 513 2261 516
rect 2218 403 2221 416
rect 2226 403 2229 416
rect 2226 333 2229 366
rect 2202 323 2221 326
rect 2202 213 2205 226
rect 2210 196 2213 323
rect 2226 303 2229 326
rect 2234 236 2237 513
rect 2250 413 2253 426
rect 2242 393 2245 406
rect 2250 403 2261 406
rect 2266 403 2269 526
rect 2242 253 2245 336
rect 2250 323 2253 356
rect 2258 323 2261 336
rect 2266 333 2269 366
rect 2274 306 2277 536
rect 2282 383 2285 596
rect 2290 506 2293 603
rect 2298 593 2301 643
rect 2306 603 2309 636
rect 2314 583 2317 706
rect 2322 696 2325 783
rect 2322 693 2329 696
rect 2326 626 2329 693
rect 2338 686 2341 776
rect 2354 753 2365 756
rect 2362 723 2365 753
rect 2370 693 2373 983
rect 2378 813 2381 993
rect 2394 983 2405 986
rect 2386 823 2389 926
rect 2394 896 2397 983
rect 2410 976 2413 993
rect 2418 983 2421 1023
rect 2426 993 2429 1006
rect 2410 973 2421 976
rect 2402 903 2405 936
rect 2394 893 2401 896
rect 2398 826 2401 893
rect 2410 883 2413 926
rect 2418 913 2421 973
rect 2426 903 2429 926
rect 2434 923 2437 1016
rect 2442 943 2445 1005
rect 2450 923 2453 1023
rect 2434 913 2445 916
rect 2434 886 2437 906
rect 2430 883 2437 886
rect 2398 823 2405 826
rect 2338 683 2365 686
rect 2322 623 2329 626
rect 2322 566 2325 623
rect 2330 583 2333 606
rect 2338 596 2341 616
rect 2346 603 2349 636
rect 2354 613 2357 646
rect 2354 596 2357 606
rect 2338 593 2357 596
rect 2318 563 2325 566
rect 2298 533 2301 546
rect 2290 503 2297 506
rect 2294 376 2297 503
rect 2306 486 2309 526
rect 2318 506 2321 563
rect 2338 546 2341 593
rect 2330 543 2341 546
rect 2318 503 2325 506
rect 2306 483 2317 486
rect 2306 413 2309 476
rect 2314 413 2317 483
rect 2306 393 2309 406
rect 2266 303 2277 306
rect 2290 373 2297 376
rect 2322 373 2325 503
rect 2226 233 2237 236
rect 2266 236 2269 303
rect 2266 233 2277 236
rect 2218 203 2221 216
rect 2202 193 2213 196
rect 2202 146 2205 193
rect 2226 163 2229 233
rect 2242 213 2253 216
rect 2234 203 2245 206
rect 2250 203 2253 213
rect 2242 146 2245 203
rect 2274 153 2277 233
rect 2282 203 2285 216
rect 2290 213 2293 373
rect 2330 366 2333 543
rect 2338 503 2341 536
rect 2346 523 2349 536
rect 2354 533 2357 556
rect 2354 486 2357 526
rect 2338 483 2357 486
rect 2338 403 2341 483
rect 2362 476 2365 683
rect 2378 636 2381 806
rect 2386 803 2397 806
rect 2402 803 2405 823
rect 2410 813 2413 836
rect 2418 786 2421 806
rect 2430 796 2433 883
rect 2430 793 2437 796
rect 2370 633 2381 636
rect 2370 616 2373 633
rect 2370 613 2381 616
rect 2386 613 2389 786
rect 2410 783 2421 786
rect 2410 726 2413 783
rect 2426 733 2429 776
rect 2410 723 2417 726
rect 2402 613 2405 676
rect 2414 626 2417 723
rect 2434 676 2437 793
rect 2410 623 2417 626
rect 2426 673 2437 676
rect 2370 493 2373 536
rect 2378 523 2381 613
rect 2386 506 2389 526
rect 2382 503 2389 506
rect 2354 473 2365 476
rect 2338 383 2349 386
rect 2322 363 2333 366
rect 2306 333 2309 346
rect 2314 323 2317 356
rect 2322 303 2325 363
rect 2338 333 2341 366
rect 2346 323 2349 383
rect 2306 193 2309 206
rect 2314 203 2317 246
rect 2322 203 2325 226
rect 2354 193 2357 473
rect 2382 436 2385 503
rect 2382 433 2389 436
rect 2378 393 2381 416
rect 2386 403 2389 433
rect 2394 386 2397 606
rect 2402 533 2405 606
rect 2410 553 2413 623
rect 2418 593 2421 616
rect 2426 603 2429 673
rect 2434 566 2437 616
rect 2426 563 2437 566
rect 2426 543 2429 563
rect 2410 463 2413 526
rect 2418 523 2421 536
rect 2426 523 2429 536
rect 2434 506 2437 556
rect 2426 503 2437 506
rect 2426 436 2429 503
rect 2426 433 2437 436
rect 2434 413 2437 433
rect 2390 383 2397 386
rect 2370 246 2373 336
rect 2378 323 2381 356
rect 2390 326 2393 383
rect 2402 333 2405 396
rect 2434 343 2437 366
rect 2410 333 2437 336
rect 2390 323 2397 326
rect 2370 243 2381 246
rect 2378 213 2381 243
rect 2394 223 2397 323
rect 2434 316 2437 333
rect 2418 313 2437 316
rect 2418 266 2421 313
rect 2418 263 2429 266
rect 2426 236 2429 263
rect 2426 233 2437 236
rect 2434 213 2437 233
rect 2202 143 2213 146
rect 2242 143 2253 146
rect 2210 123 2213 143
rect 2226 123 2229 136
rect 2250 123 2253 143
rect 2330 123 2333 156
rect 2354 123 2357 136
rect 2402 113 2405 126
rect 2442 123 2445 876
rect 2450 843 2453 916
rect 2458 856 2461 1006
rect 2466 933 2469 1043
rect 2474 943 2477 1093
rect 2486 1026 2489 1103
rect 2482 1023 2489 1026
rect 2482 1003 2485 1023
rect 2466 873 2469 926
rect 2474 856 2477 936
rect 2482 903 2485 926
rect 2458 853 2465 856
rect 2474 853 2485 856
rect 2450 813 2453 826
rect 2450 753 2453 806
rect 2462 746 2465 853
rect 2474 803 2477 846
rect 2482 833 2485 853
rect 2482 783 2485 826
rect 2490 776 2493 1006
rect 2498 996 2501 1133
rect 2514 1126 2517 1176
rect 2530 1166 2533 1203
rect 2538 1173 2541 1276
rect 2546 1186 2549 1363
rect 2554 1313 2557 1346
rect 2546 1183 2557 1186
rect 2530 1163 2549 1166
rect 2546 1133 2549 1163
rect 2506 1123 2517 1126
rect 2506 1013 2509 1123
rect 2514 1003 2517 1106
rect 2522 1096 2525 1126
rect 2522 1093 2529 1096
rect 2526 1026 2529 1093
rect 2526 1023 2533 1026
rect 2498 993 2505 996
rect 2502 936 2505 993
rect 2502 933 2509 936
rect 2514 933 2517 996
rect 2522 956 2525 1016
rect 2530 1003 2533 1023
rect 2522 953 2533 956
rect 2530 943 2533 953
rect 2498 893 2501 926
rect 2506 903 2509 933
rect 2482 773 2493 776
rect 2490 746 2493 766
rect 2498 756 2501 816
rect 2514 813 2517 846
rect 2506 763 2509 806
rect 2522 803 2525 926
rect 2538 906 2541 1126
rect 2554 1123 2557 1183
rect 2562 1146 2565 1433
rect 2578 1413 2581 1513
rect 2602 1433 2605 1536
rect 2618 1533 2621 1596
rect 2610 1473 2613 1526
rect 2626 1483 2629 1606
rect 2634 1583 2637 1606
rect 2646 1566 2649 1613
rect 2642 1563 2649 1566
rect 2642 1546 2645 1563
rect 2638 1543 2645 1546
rect 2638 1446 2641 1543
rect 2650 1473 2653 1536
rect 2658 1496 2661 1776
rect 2666 1653 2669 1786
rect 2674 1693 2677 1906
rect 2682 1903 2693 1906
rect 2714 1903 2717 1936
rect 2690 1846 2693 1903
rect 2682 1843 2693 1846
rect 2682 1803 2685 1843
rect 2730 1836 2733 1953
rect 2746 1933 2749 1956
rect 2730 1833 2741 1836
rect 2690 1823 2725 1826
rect 2690 1813 2693 1823
rect 2698 1736 2701 1816
rect 2706 1793 2709 1806
rect 2714 1803 2717 1816
rect 2722 1803 2725 1823
rect 2730 1803 2733 1826
rect 2682 1683 2685 1716
rect 2690 1646 2693 1736
rect 2698 1733 2717 1736
rect 2722 1733 2725 1796
rect 2738 1746 2741 1833
rect 2746 1793 2749 1826
rect 2682 1643 2693 1646
rect 2682 1613 2685 1643
rect 2690 1613 2693 1626
rect 2698 1616 2701 1726
rect 2714 1633 2717 1733
rect 2730 1726 2733 1746
rect 2738 1743 2749 1746
rect 2738 1733 2741 1743
rect 2754 1736 2757 1866
rect 2746 1733 2757 1736
rect 2762 1733 2765 1796
rect 2722 1623 2725 1726
rect 2730 1723 2741 1726
rect 2698 1613 2733 1616
rect 2658 1493 2669 1496
rect 2638 1443 2645 1446
rect 2570 1316 2573 1406
rect 2594 1393 2597 1406
rect 2578 1333 2581 1376
rect 2586 1323 2589 1366
rect 2570 1313 2577 1316
rect 2574 1256 2577 1313
rect 2574 1253 2581 1256
rect 2578 1243 2581 1253
rect 2562 1143 2573 1146
rect 2562 1113 2565 1136
rect 2546 933 2549 1056
rect 2546 916 2549 926
rect 2554 923 2557 1066
rect 2570 1003 2573 1143
rect 2578 1056 2581 1176
rect 2586 1123 2589 1316
rect 2594 1173 2597 1386
rect 2602 1373 2605 1406
rect 2602 1313 2605 1326
rect 2602 1206 2605 1246
rect 2610 1213 2613 1336
rect 2618 1326 2621 1436
rect 2642 1426 2645 1443
rect 2626 1423 2645 1426
rect 2626 1383 2629 1423
rect 2626 1333 2629 1366
rect 2618 1323 2629 1326
rect 2634 1306 2637 1416
rect 2650 1413 2653 1436
rect 2658 1406 2661 1486
rect 2642 1403 2661 1406
rect 2630 1303 2637 1306
rect 2602 1203 2613 1206
rect 2610 1156 2613 1203
rect 2630 1196 2633 1303
rect 2630 1193 2637 1196
rect 2634 1173 2637 1193
rect 2594 1133 2597 1156
rect 2602 1153 2613 1156
rect 2586 1063 2589 1116
rect 2578 1053 2597 1056
rect 2594 996 2597 1053
rect 2586 993 2597 996
rect 2562 933 2565 946
rect 2570 923 2573 966
rect 2578 916 2581 936
rect 2586 933 2589 993
rect 2602 986 2605 1153
rect 2610 1013 2613 1136
rect 2618 1056 2621 1126
rect 2626 1063 2629 1136
rect 2634 1133 2637 1156
rect 2634 1056 2637 1126
rect 2618 1053 2637 1056
rect 2642 1036 2645 1386
rect 2666 1356 2669 1493
rect 2674 1476 2677 1566
rect 2722 1563 2725 1606
rect 2698 1486 2701 1526
rect 2690 1483 2701 1486
rect 2738 1476 2741 1723
rect 2746 1716 2749 1733
rect 2746 1713 2757 1716
rect 2754 1646 2757 1713
rect 2750 1643 2757 1646
rect 2750 1546 2753 1643
rect 2762 1603 2765 1626
rect 2770 1613 2773 2123
rect 2778 2003 2781 2066
rect 2786 2013 2789 2036
rect 2794 2013 2797 2123
rect 2802 2106 2805 2166
rect 2810 2126 2813 2216
rect 2818 2133 2821 2206
rect 2826 2193 2829 2223
rect 2850 2206 2853 2236
rect 2858 2213 2861 2433
rect 2866 2373 2869 2453
rect 2874 2366 2877 2506
rect 2886 2436 2889 2513
rect 2882 2433 2889 2436
rect 2882 2413 2885 2433
rect 2866 2363 2877 2366
rect 2866 2306 2869 2363
rect 2874 2333 2877 2346
rect 2882 2336 2885 2406
rect 2890 2403 2893 2416
rect 2898 2343 2901 2506
rect 2910 2426 2913 2513
rect 2906 2423 2913 2426
rect 2906 2403 2909 2423
rect 2906 2346 2909 2396
rect 2906 2343 2917 2346
rect 2882 2333 2909 2336
rect 2914 2333 2917 2343
rect 2882 2323 2885 2333
rect 2866 2303 2877 2306
rect 2874 2236 2877 2303
rect 2866 2233 2877 2236
rect 2850 2203 2861 2206
rect 2866 2203 2869 2233
rect 2874 2196 2877 2216
rect 2890 2203 2893 2236
rect 2826 2133 2829 2166
rect 2810 2123 2829 2126
rect 2802 2103 2813 2106
rect 2810 2046 2813 2103
rect 2826 2083 2829 2123
rect 2834 2093 2837 2196
rect 2850 2156 2853 2196
rect 2874 2193 2881 2196
rect 2850 2153 2869 2156
rect 2802 2043 2813 2046
rect 2778 1953 2781 1996
rect 2778 1803 2781 1926
rect 2786 1823 2789 1966
rect 2786 1803 2789 1816
rect 2778 1663 2781 1736
rect 2786 1716 2789 1726
rect 2794 1723 2797 2006
rect 2802 1976 2805 2043
rect 2818 2003 2821 2016
rect 2842 2013 2845 2136
rect 2850 2123 2853 2153
rect 2858 2106 2861 2146
rect 2866 2126 2869 2153
rect 2878 2136 2881 2193
rect 2898 2173 2901 2326
rect 2914 2223 2917 2296
rect 2922 2216 2925 2596
rect 2930 2496 2933 2623
rect 2946 2613 2949 2683
rect 2970 2626 2973 2726
rect 2962 2623 2973 2626
rect 2978 2626 2981 2733
rect 2986 2693 2989 2726
rect 2978 2623 2989 2626
rect 2962 2606 2965 2623
rect 2946 2603 2965 2606
rect 2938 2503 2941 2596
rect 2946 2506 2949 2603
rect 2978 2593 2981 2616
rect 2986 2603 2989 2623
rect 2946 2503 2957 2506
rect 2962 2503 2965 2536
rect 2986 2513 2989 2526
rect 2930 2493 2941 2496
rect 2930 2423 2933 2456
rect 2930 2403 2933 2416
rect 2938 2413 2941 2493
rect 2946 2383 2949 2456
rect 2946 2333 2949 2366
rect 2954 2333 2957 2503
rect 2986 2473 2989 2506
rect 2994 2436 2997 2606
rect 3002 2603 3005 2756
rect 3010 2753 3021 2756
rect 3010 2723 3013 2753
rect 3026 2736 3029 2776
rect 3022 2733 3029 2736
rect 3022 2686 3025 2733
rect 3034 2693 3037 2986
rect 3082 2966 3085 3006
rect 3058 2963 3085 2966
rect 3122 2966 3125 3026
rect 3130 3003 3133 3016
rect 3122 2963 3129 2966
rect 3058 2886 3061 2963
rect 3058 2883 3069 2886
rect 3066 2803 3069 2883
rect 3098 2866 3101 2946
rect 3106 2923 3109 2936
rect 3126 2896 3129 2963
rect 3122 2893 3129 2896
rect 3122 2873 3125 2893
rect 3138 2876 3141 2926
rect 3154 2923 3157 3016
rect 3162 2983 3165 3016
rect 3178 2963 3181 3213
rect 3186 3193 3189 3206
rect 3194 3186 3197 3213
rect 3186 3183 3197 3186
rect 3202 3186 3205 3206
rect 3210 3193 3213 3353
rect 3218 3333 3221 3363
rect 3226 3346 3229 3373
rect 3234 3363 3237 3416
rect 3242 3413 3245 3453
rect 3258 3406 3261 3426
rect 3266 3413 3269 3463
rect 3250 3403 3261 3406
rect 3274 3403 3277 3513
rect 3290 3426 3293 3553
rect 3298 3533 3301 3566
rect 3314 3563 3319 3566
rect 3322 3563 3333 3566
rect 3306 3436 3309 3526
rect 3314 3506 3317 3563
rect 3322 3533 3325 3563
rect 3330 3536 3333 3546
rect 3354 3536 3357 3576
rect 3330 3533 3341 3536
rect 3346 3533 3357 3536
rect 3362 3533 3365 3546
rect 3378 3536 3381 3746
rect 3390 3716 3393 3773
rect 3402 3733 3405 3803
rect 3418 3793 3421 3846
rect 3426 3783 3429 3956
rect 3434 3823 3437 3963
rect 3458 3896 3461 3926
rect 3466 3913 3469 4016
rect 3474 3973 3477 4006
rect 3482 3983 3485 4023
rect 3490 3953 3493 4126
rect 3506 4103 3509 4126
rect 3522 4033 3525 4126
rect 3530 4123 3533 4136
rect 3554 4133 3557 4146
rect 3578 4136 3581 4153
rect 3562 4133 3581 4136
rect 3498 4023 3533 4026
rect 3498 4013 3501 4023
rect 3498 3983 3501 4006
rect 3506 3973 3509 4016
rect 3514 3983 3517 4006
rect 3474 3933 3485 3936
rect 3474 3916 3477 3926
rect 3474 3913 3485 3916
rect 3442 3813 3445 3896
rect 3458 3893 3477 3896
rect 3450 3803 3453 3836
rect 3458 3786 3461 3836
rect 3466 3796 3469 3826
rect 3474 3813 3477 3893
rect 3482 3803 3485 3866
rect 3490 3833 3493 3926
rect 3506 3913 3509 3956
rect 3522 3936 3525 4016
rect 3530 4003 3533 4023
rect 3538 3953 3541 4126
rect 3554 4043 3557 4126
rect 3522 3933 3541 3936
rect 3514 3913 3517 3926
rect 3546 3923 3549 4036
rect 3562 4026 3565 4126
rect 3578 4063 3581 4126
rect 3594 4116 3597 4166
rect 3602 4123 3605 4136
rect 3610 4123 3613 4196
rect 3618 4116 3621 4203
rect 3658 4176 3661 4243
rect 3642 4173 3661 4176
rect 3626 4133 3629 4166
rect 3594 4113 3605 4116
rect 3554 4023 3565 4026
rect 3554 4003 3557 4023
rect 3466 3793 3485 3796
rect 3490 3793 3493 3816
rect 3458 3783 3477 3786
rect 3410 3733 3413 3746
rect 3390 3713 3397 3716
rect 3410 3713 3413 3726
rect 3394 3666 3397 3713
rect 3418 3693 3421 3726
rect 3434 3713 3437 3736
rect 3466 3733 3469 3746
rect 3386 3663 3397 3666
rect 3386 3643 3389 3663
rect 3418 3616 3421 3626
rect 3386 3603 3389 3616
rect 3410 3613 3421 3616
rect 3426 3613 3429 3686
rect 3410 3596 3413 3613
rect 3434 3606 3437 3706
rect 3442 3626 3445 3716
rect 3458 3706 3461 3726
rect 3474 3723 3477 3783
rect 3482 3733 3485 3793
rect 3498 3736 3501 3896
rect 3522 3873 3525 3906
rect 3506 3813 3509 3836
rect 3506 3783 3509 3806
rect 3514 3803 3517 3816
rect 3522 3813 3525 3826
rect 3490 3733 3501 3736
rect 3514 3733 3517 3776
rect 3530 3733 3533 3916
rect 3554 3906 3557 3966
rect 3562 3936 3565 4016
rect 3570 4003 3573 4016
rect 3562 3933 3573 3936
rect 3542 3903 3557 3906
rect 3542 3826 3545 3903
rect 3542 3823 3549 3826
rect 3538 3753 3541 3816
rect 3490 3706 3493 3733
rect 3458 3703 3469 3706
rect 3466 3626 3469 3703
rect 3482 3703 3493 3706
rect 3482 3646 3485 3703
rect 3482 3643 3493 3646
rect 3442 3623 3453 3626
rect 3466 3623 3485 3626
rect 3370 3533 3381 3536
rect 3322 3513 3325 3526
rect 3314 3503 3325 3506
rect 3306 3433 3317 3436
rect 3282 3423 3309 3426
rect 3282 3413 3285 3423
rect 3290 3413 3301 3416
rect 3306 3413 3309 3423
rect 3314 3413 3317 3433
rect 3226 3343 3245 3346
rect 3242 3333 3245 3343
rect 3218 3286 3221 3326
rect 3234 3293 3237 3326
rect 3250 3323 3253 3386
rect 3258 3346 3261 3396
rect 3258 3343 3269 3346
rect 3258 3333 3261 3343
rect 3218 3283 3245 3286
rect 3274 3283 3277 3396
rect 3218 3203 3221 3276
rect 3242 3256 3245 3283
rect 3258 3263 3277 3266
rect 3242 3253 3253 3256
rect 3226 3213 3229 3246
rect 3242 3186 3245 3226
rect 3202 3183 3213 3186
rect 3186 3123 3189 3183
rect 3194 3133 3197 3156
rect 3202 3123 3205 3146
rect 3210 3083 3213 3183
rect 3226 3183 3245 3186
rect 3250 3196 3253 3253
rect 3258 3203 3261 3263
rect 3266 3213 3269 3256
rect 3274 3233 3277 3263
rect 3266 3196 3269 3206
rect 3250 3193 3269 3196
rect 3226 3123 3229 3183
rect 3234 3093 3237 3136
rect 3242 3133 3245 3176
rect 3250 3143 3253 3193
rect 3274 3186 3277 3226
rect 3282 3213 3285 3406
rect 3290 3326 3293 3336
rect 3298 3333 3301 3406
rect 3306 3356 3309 3406
rect 3314 3393 3317 3406
rect 3322 3403 3325 3503
rect 3330 3496 3333 3526
rect 3338 3523 3341 3533
rect 3346 3503 3349 3526
rect 3330 3493 3357 3496
rect 3362 3493 3365 3526
rect 3330 3406 3333 3476
rect 3346 3443 3349 3476
rect 3338 3413 3341 3426
rect 3354 3413 3357 3493
rect 3370 3476 3373 3533
rect 3362 3473 3373 3476
rect 3330 3403 3341 3406
rect 3354 3366 3357 3406
rect 3338 3363 3357 3366
rect 3306 3353 3317 3356
rect 3306 3333 3309 3346
rect 3290 3323 3301 3326
rect 3290 3293 3293 3316
rect 3258 3183 3277 3186
rect 3258 3076 3261 3183
rect 3290 3176 3293 3216
rect 3266 3173 3293 3176
rect 3266 3083 3269 3173
rect 3290 3143 3293 3173
rect 3282 3083 3285 3126
rect 3290 3123 3293 3136
rect 3298 3133 3301 3323
rect 3306 3203 3309 3216
rect 3298 3076 3301 3126
rect 3314 3103 3317 3353
rect 3322 3313 3333 3316
rect 3338 3306 3341 3363
rect 3362 3356 3365 3473
rect 3378 3466 3381 3526
rect 3386 3516 3389 3596
rect 3394 3593 3413 3596
rect 3418 3596 3421 3606
rect 3426 3603 3437 3606
rect 3458 3613 3477 3616
rect 3458 3603 3461 3613
rect 3418 3593 3461 3596
rect 3394 3523 3397 3593
rect 3474 3586 3477 3596
rect 3386 3513 3397 3516
rect 3370 3463 3381 3466
rect 3370 3413 3381 3416
rect 3386 3413 3389 3496
rect 3394 3413 3397 3513
rect 3402 3473 3405 3586
rect 3450 3583 3477 3586
rect 3410 3536 3413 3566
rect 3410 3533 3437 3536
rect 3410 3493 3413 3526
rect 3426 3513 3429 3526
rect 3410 3456 3413 3466
rect 3402 3453 3413 3456
rect 3402 3406 3405 3453
rect 3418 3413 3421 3426
rect 3426 3413 3429 3496
rect 3434 3413 3437 3533
rect 3442 3523 3445 3556
rect 3442 3503 3445 3516
rect 3450 3463 3453 3583
rect 3458 3533 3461 3576
rect 3442 3423 3453 3426
rect 3442 3413 3445 3423
rect 3346 3353 3365 3356
rect 3346 3333 3349 3353
rect 3330 3303 3341 3306
rect 3346 3303 3349 3326
rect 3330 3263 3333 3303
rect 3322 3213 3325 3226
rect 3322 3193 3325 3206
rect 3330 3143 3333 3216
rect 3338 3136 3341 3246
rect 3346 3206 3349 3296
rect 3354 3256 3357 3346
rect 3362 3273 3365 3326
rect 3370 3293 3373 3406
rect 3378 3383 3381 3406
rect 3378 3276 3381 3326
rect 3386 3303 3389 3326
rect 3378 3273 3389 3276
rect 3386 3263 3389 3273
rect 3354 3253 3389 3256
rect 3354 3233 3381 3236
rect 3354 3223 3357 3233
rect 3386 3226 3389 3253
rect 3364 3224 3367 3226
rect 3362 3221 3367 3224
rect 3378 3223 3389 3226
rect 3362 3216 3365 3221
rect 3354 3213 3365 3216
rect 3346 3203 3357 3206
rect 3330 3133 3341 3136
rect 3330 3123 3333 3133
rect 3346 3123 3349 3186
rect 3346 3083 3349 3116
rect 3354 3093 3357 3203
rect 3258 3073 3301 3076
rect 3362 3053 3365 3206
rect 3370 3133 3373 3146
rect 3378 3133 3381 3223
rect 3386 3186 3389 3216
rect 3394 3203 3397 3406
rect 3402 3403 3421 3406
rect 3402 3256 3405 3396
rect 3418 3333 3421 3386
rect 3434 3376 3437 3406
rect 3442 3403 3453 3406
rect 3426 3373 3437 3376
rect 3458 3373 3461 3446
rect 3426 3343 3429 3373
rect 3410 3313 3413 3326
rect 3418 3323 3429 3326
rect 3418 3263 3421 3323
rect 3402 3253 3413 3256
rect 3402 3213 3405 3246
rect 3410 3206 3413 3253
rect 3418 3213 3421 3246
rect 3410 3203 3421 3206
rect 3426 3203 3429 3226
rect 3434 3203 3437 3366
rect 3442 3303 3445 3326
rect 3386 3183 3405 3186
rect 3386 3153 3397 3156
rect 3386 3123 3389 3153
rect 3394 3093 3397 3136
rect 3402 3063 3405 3183
rect 3410 3093 3413 3186
rect 3418 3133 3421 3203
rect 3442 3196 3445 3266
rect 3450 3236 3453 3366
rect 3466 3343 3469 3536
rect 3474 3513 3477 3526
rect 3474 3413 3477 3496
rect 3482 3476 3485 3623
rect 3490 3603 3493 3643
rect 3498 3596 3501 3726
rect 3506 3633 3509 3726
rect 3506 3603 3509 3616
rect 3514 3613 3517 3726
rect 3522 3673 3525 3726
rect 3530 3696 3533 3726
rect 3546 3723 3549 3823
rect 3554 3813 3557 3836
rect 3562 3826 3565 3926
rect 3570 3916 3573 3933
rect 3578 3923 3581 4046
rect 3586 4003 3589 4106
rect 3594 4003 3597 4016
rect 3602 3973 3605 4113
rect 3610 4113 3621 4116
rect 3610 4083 3613 4113
rect 3626 4106 3629 4126
rect 3618 4103 3629 4106
rect 3586 3933 3589 3956
rect 3594 3936 3597 3966
rect 3594 3933 3605 3936
rect 3610 3933 3613 4006
rect 3570 3913 3581 3916
rect 3562 3823 3573 3826
rect 3578 3823 3581 3913
rect 3586 3893 3589 3926
rect 3602 3916 3605 3933
rect 3618 3923 3621 4103
rect 3642 4056 3645 4173
rect 3650 4063 3653 4126
rect 3658 4083 3661 4136
rect 3666 4123 3669 4196
rect 3674 4106 3677 4286
rect 3698 4256 3701 4276
rect 3698 4253 3705 4256
rect 3670 4103 3677 4106
rect 3634 4053 3645 4056
rect 3634 4033 3637 4053
rect 3634 3973 3637 4006
rect 3658 3983 3661 4016
rect 3670 3956 3673 4103
rect 3682 4003 3685 4216
rect 3702 4186 3705 4253
rect 3698 4183 3705 4186
rect 3698 4156 3701 4183
rect 3714 4166 3717 4337
rect 3730 4203 3733 4306
rect 3762 4286 3765 4340
rect 3762 4283 3769 4286
rect 3754 4213 3757 4276
rect 3766 4206 3769 4283
rect 3762 4203 3769 4206
rect 3706 4163 3717 4166
rect 3698 4153 3725 4156
rect 3690 4143 3717 4146
rect 3690 4056 3693 4143
rect 3698 4103 3701 4126
rect 3690 4053 3701 4056
rect 3650 3953 3673 3956
rect 3626 3926 3629 3936
rect 3634 3933 3645 3936
rect 3626 3923 3637 3926
rect 3602 3913 3621 3916
rect 3562 3803 3565 3816
rect 3570 3796 3573 3823
rect 3554 3793 3573 3796
rect 3578 3793 3581 3816
rect 3538 3706 3541 3716
rect 3554 3713 3557 3793
rect 3562 3723 3565 3756
rect 3586 3753 3589 3836
rect 3594 3773 3597 3826
rect 3578 3713 3581 3746
rect 3586 3723 3589 3736
rect 3594 3706 3597 3746
rect 3602 3733 3605 3826
rect 3618 3806 3621 3913
rect 3642 3893 3645 3933
rect 3650 3843 3653 3953
rect 3682 3946 3685 3966
rect 3698 3946 3701 4053
rect 3658 3943 3685 3946
rect 3690 3943 3701 3946
rect 3706 3986 3709 4136
rect 3714 4123 3717 4143
rect 3722 4133 3725 4153
rect 3730 4096 3733 4126
rect 3738 4103 3741 4136
rect 3746 4133 3749 4186
rect 3746 4096 3749 4126
rect 3730 4093 3749 4096
rect 3754 4086 3757 4106
rect 3730 4083 3757 4086
rect 3714 4013 3717 4036
rect 3706 3983 3717 3986
rect 3666 3926 3669 3936
rect 3674 3933 3685 3936
rect 3666 3923 3685 3926
rect 3626 3823 3661 3826
rect 3626 3813 3629 3823
rect 3610 3796 3613 3806
rect 3618 3803 3629 3806
rect 3634 3796 3637 3816
rect 3610 3793 3637 3796
rect 3642 3793 3645 3806
rect 3650 3796 3653 3816
rect 3658 3803 3661 3823
rect 3666 3796 3669 3816
rect 3674 3803 3677 3866
rect 3682 3833 3685 3923
rect 3690 3906 3693 3943
rect 3698 3913 3701 3936
rect 3706 3933 3709 3983
rect 3714 3933 3717 3966
rect 3722 3926 3725 3956
rect 3706 3923 3725 3926
rect 3690 3903 3697 3906
rect 3694 3836 3697 3903
rect 3730 3893 3733 4083
rect 3762 4043 3765 4203
rect 3778 4166 3781 4340
rect 3794 4183 3797 4340
rect 3810 4293 3813 4340
rect 3842 4296 3845 4340
rect 3818 4293 3845 4296
rect 3818 4286 3821 4293
rect 3810 4283 3821 4286
rect 3802 4176 3805 4196
rect 3770 4163 3781 4166
rect 3794 4173 3805 4176
rect 3770 4103 3773 4163
rect 3778 4063 3781 4126
rect 3786 4103 3789 4136
rect 3794 4123 3797 4173
rect 3802 4123 3805 4136
rect 3810 4056 3813 4283
rect 3826 4213 3829 4256
rect 3818 4183 3821 4206
rect 3834 4203 3837 4286
rect 3842 4196 3845 4216
rect 3850 4203 3853 4326
rect 3922 4286 3925 4340
rect 3898 4283 3925 4286
rect 3858 4213 3861 4256
rect 3834 4193 3845 4196
rect 3858 4196 3861 4206
rect 3874 4203 3877 4216
rect 3858 4193 3877 4196
rect 3882 4193 3885 4216
rect 3818 4063 3821 4126
rect 3802 4053 3813 4056
rect 3778 4043 3797 4046
rect 3754 4013 3757 4036
rect 3778 4016 3781 4043
rect 3738 4003 3749 4006
rect 3738 3886 3741 4003
rect 3754 3983 3757 4006
rect 3762 4003 3765 4016
rect 3770 4013 3781 4016
rect 3770 4003 3781 4006
rect 3786 4003 3789 4036
rect 3794 4013 3797 4043
rect 3802 4003 3805 4053
rect 3810 3996 3813 4046
rect 3826 4043 3829 4136
rect 3834 4123 3837 4193
rect 3842 4036 3845 4136
rect 3850 4093 3853 4136
rect 3866 4133 3869 4186
rect 3874 4156 3877 4193
rect 3890 4163 3893 4206
rect 3898 4156 3901 4283
rect 3874 4153 3901 4156
rect 3858 4116 3861 4126
rect 3874 4123 3877 4146
rect 3906 4143 3909 4216
rect 3922 4156 3925 4266
rect 3946 4183 3949 4216
rect 3954 4176 3957 4326
rect 3914 4153 3925 4156
rect 3938 4173 3957 4176
rect 3882 4126 3885 4136
rect 3890 4133 3901 4136
rect 3882 4123 3893 4126
rect 3898 4116 3901 4133
rect 3914 4126 3917 4153
rect 3858 4113 3901 4116
rect 3898 4056 3901 4113
rect 3910 4123 3917 4126
rect 3910 4076 3913 4123
rect 3922 4093 3925 4146
rect 3922 4083 3933 4086
rect 3910 4073 3917 4076
rect 3802 3993 3813 3996
rect 3826 4033 3845 4036
rect 3882 4053 3901 4056
rect 3706 3883 3741 3886
rect 3694 3833 3701 3836
rect 3682 3813 3693 3816
rect 3650 3793 3669 3796
rect 3610 3723 3613 3776
rect 3618 3726 3621 3736
rect 3626 3733 3629 3746
rect 3618 3723 3629 3726
rect 3538 3703 3557 3706
rect 3530 3693 3549 3696
rect 3530 3666 3533 3686
rect 3546 3666 3549 3693
rect 3554 3673 3557 3703
rect 3562 3696 3565 3706
rect 3570 3703 3581 3706
rect 3590 3703 3597 3706
rect 3562 3693 3581 3696
rect 3522 3663 3533 3666
rect 3538 3663 3549 3666
rect 3522 3613 3525 3663
rect 3514 3603 3525 3606
rect 3490 3593 3501 3596
rect 3490 3533 3493 3593
rect 3530 3563 3533 3636
rect 3538 3603 3541 3663
rect 3546 3643 3549 3656
rect 3490 3483 3493 3526
rect 3498 3523 3501 3536
rect 3482 3473 3501 3476
rect 3482 3406 3485 3466
rect 3490 3413 3493 3426
rect 3474 3403 3485 3406
rect 3474 3393 3477 3403
rect 3490 3396 3493 3406
rect 3482 3393 3493 3396
rect 3474 3333 3477 3376
rect 3482 3346 3485 3393
rect 3498 3386 3501 3473
rect 3506 3463 3509 3536
rect 3522 3533 3525 3556
rect 3514 3503 3517 3526
rect 3506 3413 3509 3446
rect 3490 3383 3501 3386
rect 3506 3366 3509 3406
rect 3514 3403 3517 3496
rect 3522 3403 3525 3526
rect 3530 3483 3533 3526
rect 3538 3523 3541 3536
rect 3530 3393 3533 3416
rect 3498 3363 3509 3366
rect 3514 3356 3517 3366
rect 3498 3353 3517 3356
rect 3482 3343 3493 3346
rect 3458 3293 3461 3326
rect 3466 3323 3477 3326
rect 3450 3233 3477 3236
rect 3450 3223 3461 3226
rect 3426 3193 3445 3196
rect 3450 3203 3461 3206
rect 3450 3183 3453 3203
rect 3442 3083 3445 3126
rect 3450 3103 3453 3136
rect 3458 3133 3461 3176
rect 3458 3063 3461 3126
rect 3466 3093 3469 3216
rect 3474 3173 3477 3233
rect 3482 3193 3485 3336
rect 3490 3333 3493 3343
rect 3498 3333 3501 3353
rect 3522 3333 3525 3376
rect 3490 3303 3493 3326
rect 3498 3316 3501 3326
rect 3506 3323 3517 3326
rect 3522 3316 3525 3326
rect 3498 3313 3525 3316
rect 3490 3146 3493 3216
rect 3498 3213 3509 3216
rect 3514 3206 3517 3306
rect 3482 3143 3493 3146
rect 3482 3093 3485 3143
rect 3498 3136 3501 3206
rect 3490 3133 3501 3136
rect 3506 3203 3517 3206
rect 3522 3203 3525 3256
rect 3490 3053 3493 3133
rect 3498 3103 3501 3126
rect 3506 3123 3509 3203
rect 3530 3196 3533 3346
rect 3538 3303 3541 3496
rect 3546 3476 3549 3606
rect 3554 3546 3557 3616
rect 3570 3613 3573 3636
rect 3578 3583 3581 3693
rect 3590 3636 3593 3703
rect 3590 3633 3597 3636
rect 3554 3543 3565 3546
rect 3554 3523 3557 3536
rect 3562 3533 3565 3543
rect 3570 3533 3573 3566
rect 3586 3556 3589 3616
rect 3594 3613 3597 3633
rect 3602 3613 3605 3686
rect 3594 3583 3597 3606
rect 3578 3553 3589 3556
rect 3562 3523 3573 3526
rect 3578 3483 3581 3553
rect 3586 3493 3589 3536
rect 3594 3506 3597 3536
rect 3610 3526 3613 3666
rect 3618 3623 3621 3656
rect 3634 3636 3637 3793
rect 3650 3783 3653 3793
rect 3682 3773 3685 3813
rect 3690 3783 3693 3806
rect 3642 3713 3645 3746
rect 3674 3743 3693 3746
rect 3658 3653 3661 3736
rect 3666 3723 3669 3736
rect 3634 3633 3653 3636
rect 3626 3613 3645 3616
rect 3626 3603 3629 3613
rect 3650 3603 3653 3633
rect 3626 3573 3629 3596
rect 3658 3563 3661 3626
rect 3666 3613 3669 3666
rect 3674 3606 3677 3743
rect 3690 3726 3693 3736
rect 3698 3733 3701 3833
rect 3706 3786 3709 3883
rect 3746 3876 3749 3976
rect 3762 3933 3765 3956
rect 3786 3913 3789 3926
rect 3722 3873 3749 3876
rect 3722 3803 3725 3873
rect 3754 3813 3757 3826
rect 3706 3783 3717 3786
rect 3706 3733 3709 3746
rect 3682 3713 3685 3726
rect 3690 3723 3709 3726
rect 3714 3716 3717 3783
rect 3710 3713 3717 3716
rect 3682 3623 3685 3636
rect 3666 3603 3677 3606
rect 3698 3603 3701 3676
rect 3710 3636 3713 3713
rect 3706 3633 3713 3636
rect 3706 3603 3709 3633
rect 3722 3616 3725 3736
rect 3730 3666 3733 3736
rect 3738 3723 3741 3766
rect 3746 3743 3765 3746
rect 3746 3673 3749 3743
rect 3762 3726 3765 3736
rect 3730 3663 3749 3666
rect 3626 3533 3629 3546
rect 3602 3523 3621 3526
rect 3594 3503 3601 3506
rect 3618 3503 3621 3516
rect 3546 3473 3565 3476
rect 3546 3463 3557 3466
rect 3546 3413 3549 3463
rect 3554 3403 3557 3416
rect 3562 3363 3565 3473
rect 3570 3413 3573 3446
rect 3570 3383 3573 3406
rect 3578 3373 3581 3476
rect 3586 3413 3589 3466
rect 3598 3436 3601 3503
rect 3634 3476 3637 3536
rect 3666 3533 3669 3603
rect 3642 3523 3661 3526
rect 3650 3513 3661 3516
rect 3594 3433 3601 3436
rect 3626 3473 3637 3476
rect 3594 3356 3597 3433
rect 3610 3423 3621 3426
rect 3602 3403 3605 3416
rect 3618 3403 3621 3416
rect 3626 3396 3629 3473
rect 3554 3353 3597 3356
rect 3602 3393 3629 3396
rect 3554 3343 3557 3353
rect 3602 3346 3605 3393
rect 3570 3333 3573 3346
rect 3578 3343 3605 3346
rect 3546 3323 3565 3326
rect 3554 3313 3565 3316
rect 3578 3253 3581 3343
rect 3602 3326 3605 3336
rect 3610 3333 3613 3366
rect 3586 3246 3589 3326
rect 3522 3193 3533 3196
rect 3538 3213 3557 3216
rect 3522 3133 3525 3193
rect 3538 3166 3541 3213
rect 3554 3193 3557 3206
rect 3530 3163 3541 3166
rect 3514 3063 3517 3126
rect 3530 3123 3533 3163
rect 3562 3153 3565 3226
rect 3570 3203 3573 3246
rect 3578 3243 3589 3246
rect 3594 3323 3605 3326
rect 3578 3186 3581 3243
rect 3594 3236 3597 3323
rect 3602 3273 3605 3316
rect 3570 3183 3581 3186
rect 3586 3233 3597 3236
rect 3538 3033 3541 3136
rect 3562 3123 3565 3136
rect 3562 3083 3565 3116
rect 3570 3043 3573 3183
rect 3578 3133 3581 3176
rect 3586 3133 3589 3233
rect 3594 3093 3597 3226
rect 3602 3193 3605 3266
rect 3610 3203 3613 3256
rect 3610 3103 3613 3116
rect 3618 3053 3621 3376
rect 3634 3353 3637 3416
rect 3642 3396 3645 3496
rect 3650 3403 3653 3506
rect 3674 3446 3677 3536
rect 3698 3533 3701 3596
rect 3714 3593 3717 3616
rect 3722 3613 3733 3616
rect 3746 3613 3749 3663
rect 3754 3623 3757 3726
rect 3762 3723 3781 3726
rect 3722 3583 3725 3606
rect 3730 3586 3733 3613
rect 3746 3593 3749 3606
rect 3730 3583 3749 3586
rect 3706 3533 3709 3546
rect 3698 3513 3701 3526
rect 3666 3443 3677 3446
rect 3642 3393 3653 3396
rect 3650 3353 3653 3393
rect 3658 3383 3661 3426
rect 3634 3333 3645 3336
rect 3626 3323 3645 3326
rect 3626 3303 3629 3323
rect 3642 3293 3645 3316
rect 3650 3306 3653 3336
rect 3666 3313 3669 3443
rect 3674 3433 3709 3436
rect 3674 3403 3677 3433
rect 3690 3393 3693 3426
rect 3698 3413 3701 3426
rect 3706 3413 3709 3433
rect 3714 3406 3717 3566
rect 3722 3533 3725 3576
rect 3730 3523 3733 3546
rect 3738 3533 3741 3566
rect 3746 3523 3749 3583
rect 3754 3563 3757 3606
rect 3754 3506 3757 3556
rect 3746 3503 3757 3506
rect 3746 3446 3749 3503
rect 3762 3493 3765 3606
rect 3770 3553 3773 3656
rect 3770 3533 3773 3546
rect 3770 3513 3773 3526
rect 3778 3513 3781 3626
rect 3786 3573 3789 3836
rect 3794 3733 3797 3966
rect 3802 3783 3805 3993
rect 3810 3843 3813 3946
rect 3802 3716 3805 3736
rect 3810 3723 3813 3736
rect 3818 3733 3821 3886
rect 3826 3863 3829 4033
rect 3834 3803 3837 3976
rect 3842 3953 3845 4006
rect 3866 4003 3869 4016
rect 3882 3996 3885 4053
rect 3914 4026 3917 4073
rect 3906 4023 3917 4026
rect 3882 3993 3893 3996
rect 3842 3893 3845 3926
rect 3858 3786 3861 3986
rect 3874 3946 3877 3976
rect 3890 3963 3893 3993
rect 3874 3943 3885 3946
rect 3882 3933 3885 3943
rect 3906 3933 3909 4023
rect 3914 4013 3925 4016
rect 3930 4013 3933 4083
rect 3938 4043 3941 4173
rect 3962 4166 3965 4296
rect 3954 4163 3965 4166
rect 3946 4123 3949 4136
rect 3954 4123 3957 4163
rect 3970 4133 3973 4226
rect 3978 4126 3981 4146
rect 3962 4123 3981 4126
rect 3962 4106 3965 4123
rect 3986 4116 3989 4136
rect 3994 4123 3997 4226
rect 4002 4213 4005 4286
rect 4010 4213 4013 4276
rect 4010 4166 4013 4206
rect 4002 4163 4013 4166
rect 4002 4133 4005 4163
rect 4010 4133 4013 4146
rect 4018 4136 4021 4246
rect 4026 4223 4069 4226
rect 4026 4213 4037 4216
rect 4034 4146 4037 4206
rect 4042 4203 4061 4206
rect 4066 4203 4069 4216
rect 4074 4213 4077 4236
rect 4098 4223 4101 4316
rect 4090 4213 4101 4216
rect 4122 4213 4125 4256
rect 4154 4226 4157 4316
rect 4150 4223 4157 4226
rect 4090 4206 4093 4213
rect 4074 4203 4093 4206
rect 4098 4203 4125 4206
rect 4130 4203 4133 4216
rect 4058 4146 4061 4203
rect 4122 4196 4125 4203
rect 4138 4196 4141 4216
rect 4106 4156 4109 4196
rect 4122 4193 4141 4196
rect 4098 4153 4109 4156
rect 4026 4143 4037 4146
rect 4018 4133 4029 4136
rect 4042 4133 4045 4146
rect 4058 4143 4093 4146
rect 4002 4123 4013 4126
rect 3954 4103 3965 4106
rect 3954 4026 3957 4103
rect 3978 4096 3981 4116
rect 3986 4113 4005 4116
rect 3986 4103 3997 4106
rect 4002 4103 4005 4113
rect 3970 4036 3973 4096
rect 3978 4093 3989 4096
rect 3978 4046 3981 4093
rect 3978 4043 3989 4046
rect 3970 4033 3981 4036
rect 3954 4023 3969 4026
rect 3954 3973 3957 4006
rect 3914 3933 3949 3936
rect 3914 3926 3917 3933
rect 3946 3926 3949 3933
rect 3866 3923 3917 3926
rect 3882 3856 3885 3906
rect 3878 3853 3885 3856
rect 3866 3793 3869 3816
rect 3858 3783 3869 3786
rect 3818 3716 3821 3726
rect 3802 3713 3821 3716
rect 3834 3713 3837 3736
rect 3842 3733 3853 3736
rect 3842 3723 3861 3726
rect 3794 3623 3797 3636
rect 3794 3603 3797 3616
rect 3802 3613 3805 3626
rect 3810 3606 3813 3696
rect 3802 3603 3813 3606
rect 3802 3583 3805 3603
rect 3818 3556 3821 3713
rect 3866 3653 3869 3783
rect 3878 3766 3881 3853
rect 3914 3813 3917 3866
rect 3914 3803 3925 3806
rect 3878 3763 3885 3766
rect 3874 3733 3877 3746
rect 3794 3553 3821 3556
rect 3786 3496 3789 3536
rect 3782 3493 3789 3496
rect 3722 3423 3725 3446
rect 3730 3443 3749 3446
rect 3698 3403 3717 3406
rect 3730 3403 3733 3443
rect 3738 3416 3741 3436
rect 3738 3413 3749 3416
rect 3698 3386 3701 3403
rect 3682 3383 3701 3386
rect 3674 3313 3677 3326
rect 3682 3306 3685 3383
rect 3738 3376 3741 3406
rect 3690 3333 3693 3376
rect 3698 3373 3741 3376
rect 3698 3333 3701 3373
rect 3730 3336 3733 3356
rect 3746 3346 3749 3413
rect 3762 3393 3765 3456
rect 3770 3403 3773 3446
rect 3782 3416 3785 3493
rect 3778 3413 3785 3416
rect 3770 3363 3773 3396
rect 3778 3383 3781 3413
rect 3794 3406 3797 3553
rect 3802 3543 3821 3546
rect 3802 3503 3805 3543
rect 3818 3526 3821 3536
rect 3826 3533 3829 3636
rect 3850 3613 3869 3616
rect 3850 3603 3853 3613
rect 3874 3603 3877 3726
rect 3882 3633 3885 3763
rect 3890 3706 3893 3766
rect 3930 3736 3933 3926
rect 3946 3923 3957 3926
rect 3938 3783 3941 3796
rect 3890 3703 3897 3706
rect 3894 3636 3897 3703
rect 3894 3633 3901 3636
rect 3882 3613 3893 3616
rect 3898 3603 3901 3633
rect 3906 3623 3909 3736
rect 3930 3733 3941 3736
rect 3930 3713 3933 3726
rect 3938 3663 3941 3733
rect 3946 3683 3949 3856
rect 3906 3603 3909 3616
rect 3818 3523 3837 3526
rect 3810 3453 3813 3516
rect 3802 3413 3805 3446
rect 3818 3416 3821 3436
rect 3834 3423 3837 3456
rect 3842 3423 3845 3596
rect 3850 3533 3853 3546
rect 3850 3513 3853 3526
rect 3858 3496 3861 3566
rect 3866 3536 3869 3586
rect 3874 3553 3877 3596
rect 3914 3583 3917 3616
rect 3890 3573 3925 3576
rect 3930 3573 3933 3606
rect 3890 3543 3893 3573
rect 3866 3533 3873 3536
rect 3854 3493 3861 3496
rect 3854 3416 3857 3493
rect 3870 3466 3873 3533
rect 3890 3526 3893 3536
rect 3898 3533 3901 3556
rect 3906 3533 3909 3546
rect 3882 3513 3885 3526
rect 3890 3523 3909 3526
rect 3914 3516 3917 3566
rect 3870 3463 3877 3466
rect 3866 3423 3869 3456
rect 3818 3413 3837 3416
rect 3842 3413 3857 3416
rect 3786 3403 3797 3406
rect 3746 3343 3781 3346
rect 3722 3326 3725 3336
rect 3730 3333 3741 3336
rect 3650 3303 3685 3306
rect 3706 3303 3709 3326
rect 3714 3323 3725 3326
rect 3626 3196 3629 3226
rect 3634 3203 3637 3276
rect 3674 3243 3677 3303
rect 3642 3223 3661 3226
rect 3642 3213 3645 3223
rect 3658 3216 3661 3223
rect 3642 3196 3645 3206
rect 3626 3193 3645 3196
rect 3650 3166 3653 3216
rect 3658 3213 3669 3216
rect 3666 3203 3669 3213
rect 3666 3193 3677 3196
rect 3626 3163 3653 3166
rect 3682 3163 3685 3226
rect 3714 3213 3717 3323
rect 3722 3213 3725 3316
rect 3730 3306 3733 3326
rect 3738 3323 3741 3333
rect 3754 3316 3757 3336
rect 3750 3313 3757 3316
rect 3730 3303 3741 3306
rect 3738 3246 3741 3303
rect 3730 3243 3741 3246
rect 3706 3163 3709 3206
rect 3714 3193 3717 3206
rect 3730 3193 3733 3243
rect 3750 3226 3753 3313
rect 3746 3223 3753 3226
rect 3746 3213 3749 3223
rect 3738 3183 3741 3206
rect 3746 3186 3749 3206
rect 3754 3193 3757 3216
rect 3762 3206 3765 3336
rect 3770 3213 3773 3326
rect 3778 3323 3781 3343
rect 3786 3233 3789 3403
rect 3794 3313 3797 3396
rect 3802 3383 3805 3406
rect 3810 3336 3813 3406
rect 3834 3393 3837 3406
rect 3842 3356 3845 3413
rect 3874 3406 3877 3463
rect 3882 3413 3885 3506
rect 3874 3403 3885 3406
rect 3874 3373 3877 3396
rect 3826 3353 3845 3356
rect 3802 3313 3805 3336
rect 3810 3333 3821 3336
rect 3810 3216 3813 3326
rect 3818 3323 3821 3333
rect 3818 3223 3821 3246
rect 3794 3213 3813 3216
rect 3762 3203 3789 3206
rect 3762 3186 3765 3203
rect 3746 3183 3765 3186
rect 3626 3073 3629 3163
rect 3634 3133 3637 3156
rect 3730 3143 3741 3146
rect 3650 3123 3653 3136
rect 3194 3023 3229 3026
rect 3194 3013 3197 3023
rect 3202 3013 3213 3016
rect 3194 2973 3197 3006
rect 3202 3003 3213 3006
rect 3218 2993 3221 3016
rect 3226 3003 3229 3023
rect 3234 2986 3237 3006
rect 3250 3003 3253 3016
rect 3210 2983 3237 2986
rect 3162 2933 3173 2936
rect 3178 2933 3189 2936
rect 3146 2886 3149 2906
rect 3146 2883 3153 2886
rect 3134 2873 3141 2876
rect 3094 2863 3101 2866
rect 3094 2796 3097 2863
rect 3094 2793 3101 2796
rect 3042 2733 3045 2746
rect 3090 2743 3093 2776
rect 3022 2683 3029 2686
rect 3018 2613 3021 2646
rect 3018 2576 3021 2606
rect 3026 2593 3029 2683
rect 3042 2603 3045 2726
rect 3050 2686 3053 2726
rect 3058 2703 3061 2736
rect 3050 2683 3057 2686
rect 3066 2683 3069 2726
rect 3054 2616 3057 2683
rect 3050 2613 3057 2616
rect 3074 2613 3077 2726
rect 3002 2573 3021 2576
rect 3002 2453 3005 2573
rect 2978 2433 2997 2436
rect 2930 2323 2949 2326
rect 2954 2316 2957 2326
rect 2938 2313 2957 2316
rect 2938 2256 2941 2313
rect 2954 2293 2957 2306
rect 2914 2213 2925 2216
rect 2930 2253 2941 2256
rect 2878 2133 2893 2136
rect 2866 2123 2877 2126
rect 2858 2103 2865 2106
rect 2850 2023 2853 2096
rect 2862 2036 2865 2103
rect 2874 2066 2877 2123
rect 2874 2063 2885 2066
rect 2858 2033 2865 2036
rect 2858 2016 2861 2033
rect 2850 2013 2861 2016
rect 2842 1976 2845 1986
rect 2802 1973 2845 1976
rect 2818 1923 2829 1926
rect 2802 1716 2805 1876
rect 2786 1713 2805 1716
rect 2786 1603 2789 1646
rect 2810 1596 2813 1866
rect 2818 1803 2821 1923
rect 2826 1743 2829 1806
rect 2834 1793 2837 1973
rect 2850 1933 2853 2013
rect 2818 1733 2845 1736
rect 2818 1606 2821 1726
rect 2826 1613 2829 1666
rect 2842 1656 2845 1733
rect 2850 1723 2853 1906
rect 2866 1803 2869 1816
rect 2874 1803 2877 1926
rect 2882 1813 2885 2063
rect 2890 2033 2893 2133
rect 2898 1993 2901 2136
rect 2906 2013 2909 2206
rect 2922 2133 2925 2206
rect 2930 2133 2933 2253
rect 2938 2203 2941 2236
rect 2946 2213 2949 2226
rect 2938 2126 2941 2176
rect 2954 2143 2957 2286
rect 2858 1743 2885 1746
rect 2858 1733 2861 1743
rect 2866 1723 2869 1736
rect 2874 1723 2877 1736
rect 2882 1733 2885 1743
rect 2866 1656 2869 1706
rect 2882 1693 2885 1726
rect 2842 1653 2869 1656
rect 2818 1603 2829 1606
rect 2810 1593 2821 1596
rect 2674 1473 2681 1476
rect 2678 1386 2681 1473
rect 2730 1473 2741 1476
rect 2746 1543 2753 1546
rect 2690 1396 2693 1406
rect 2706 1396 2709 1436
rect 2714 1413 2717 1446
rect 2690 1393 2709 1396
rect 2678 1383 2701 1386
rect 2658 1353 2669 1356
rect 2650 1253 2653 1336
rect 2658 1243 2661 1353
rect 2674 1346 2677 1376
rect 2666 1343 2677 1346
rect 2682 1333 2685 1366
rect 2674 1286 2677 1326
rect 2682 1293 2685 1326
rect 2690 1286 2693 1326
rect 2674 1283 2693 1286
rect 2698 1276 2701 1383
rect 2666 1273 2701 1276
rect 2650 1213 2653 1226
rect 2666 1203 2669 1273
rect 2690 1196 2693 1216
rect 2650 1186 2653 1196
rect 2682 1193 2693 1196
rect 2650 1183 2657 1186
rect 2654 1116 2657 1183
rect 2666 1133 2669 1156
rect 2654 1113 2661 1116
rect 2638 1033 2645 1036
rect 2594 983 2605 986
rect 2546 913 2581 916
rect 2538 903 2549 906
rect 2530 826 2533 866
rect 2538 833 2541 846
rect 2530 823 2541 826
rect 2546 823 2549 903
rect 2530 803 2533 816
rect 2498 753 2509 756
rect 2462 743 2469 746
rect 2490 743 2501 746
rect 2450 723 2453 736
rect 2458 673 2461 736
rect 2466 716 2469 743
rect 2474 733 2485 736
rect 2466 713 2473 716
rect 2470 666 2473 713
rect 2466 663 2473 666
rect 2450 603 2453 616
rect 2466 596 2469 663
rect 2482 626 2485 726
rect 2490 633 2493 736
rect 2498 726 2501 743
rect 2506 736 2509 753
rect 2506 733 2517 736
rect 2498 723 2509 726
rect 2482 623 2493 626
rect 2450 583 2453 596
rect 2458 593 2469 596
rect 2474 613 2485 616
rect 2450 463 2453 536
rect 2458 473 2461 593
rect 2474 586 2477 613
rect 2466 583 2477 586
rect 2466 533 2469 583
rect 2482 563 2485 606
rect 2490 596 2493 623
rect 2498 603 2501 706
rect 2514 626 2517 733
rect 2522 703 2525 786
rect 2538 726 2541 823
rect 2546 733 2549 806
rect 2554 796 2557 896
rect 2562 803 2565 906
rect 2586 903 2589 926
rect 2594 906 2597 983
rect 2638 966 2641 1033
rect 2638 963 2645 966
rect 2626 943 2637 946
rect 2594 903 2605 906
rect 2554 793 2565 796
rect 2554 733 2557 746
rect 2538 723 2557 726
rect 2546 706 2549 716
rect 2530 703 2549 706
rect 2554 703 2557 723
rect 2562 713 2565 793
rect 2570 733 2573 836
rect 2586 833 2589 846
rect 2578 773 2581 826
rect 2586 803 2589 826
rect 2506 623 2517 626
rect 2506 606 2509 623
rect 2514 613 2525 616
rect 2530 613 2533 703
rect 2506 603 2517 606
rect 2490 593 2501 596
rect 2474 503 2477 526
rect 2482 523 2485 536
rect 2490 483 2493 526
rect 2458 383 2461 406
rect 2482 346 2485 416
rect 2498 393 2501 593
rect 2506 463 2509 586
rect 2514 516 2517 603
rect 2522 593 2525 613
rect 2538 586 2541 696
rect 2578 643 2581 736
rect 2586 693 2589 726
rect 2594 636 2597 896
rect 2602 856 2605 903
rect 2610 863 2613 936
rect 2634 923 2637 943
rect 2642 893 2645 963
rect 2650 913 2653 1096
rect 2602 853 2613 856
rect 2602 783 2605 836
rect 2610 813 2613 853
rect 2602 746 2605 756
rect 2618 753 2621 826
rect 2634 816 2637 846
rect 2626 746 2629 816
rect 2634 813 2645 816
rect 2634 763 2637 806
rect 2650 803 2653 876
rect 2658 803 2661 1113
rect 2666 1086 2669 1116
rect 2674 1093 2677 1176
rect 2682 1133 2685 1193
rect 2682 1123 2693 1126
rect 2666 1083 2677 1086
rect 2666 993 2669 1026
rect 2674 1013 2677 1083
rect 2674 913 2677 1006
rect 2682 1003 2685 1116
rect 2690 1063 2693 1123
rect 2698 1086 2701 1273
rect 2706 1243 2709 1393
rect 2730 1366 2733 1473
rect 2746 1456 2749 1543
rect 2742 1453 2749 1456
rect 2742 1396 2745 1453
rect 2754 1433 2757 1526
rect 2770 1506 2773 1526
rect 2770 1503 2781 1506
rect 2778 1436 2781 1503
rect 2802 1486 2805 1536
rect 2818 1533 2821 1593
rect 2810 1516 2813 1526
rect 2826 1523 2829 1603
rect 2858 1563 2861 1646
rect 2866 1613 2869 1653
rect 2874 1603 2877 1616
rect 2834 1516 2837 1556
rect 2882 1533 2885 1616
rect 2890 1553 2893 1926
rect 2914 1876 2917 2126
rect 2926 2123 2941 2126
rect 2926 1986 2929 2123
rect 2946 2096 2949 2136
rect 2954 2123 2957 2136
rect 2910 1873 2917 1876
rect 2922 1983 2929 1986
rect 2938 2093 2949 2096
rect 2910 1826 2913 1873
rect 2898 1603 2901 1826
rect 2906 1823 2913 1826
rect 2906 1733 2909 1823
rect 2922 1816 2925 1983
rect 2938 1933 2941 2093
rect 2946 2013 2949 2086
rect 2954 1956 2957 2006
rect 2946 1953 2957 1956
rect 2914 1813 2925 1816
rect 2906 1663 2909 1716
rect 2914 1556 2917 1813
rect 2930 1806 2933 1926
rect 2946 1866 2949 1953
rect 2954 1893 2957 1946
rect 2922 1803 2933 1806
rect 2942 1863 2949 1866
rect 2942 1796 2945 1863
rect 2962 1813 2965 2406
rect 2970 2093 2973 2416
rect 2978 2413 2981 2433
rect 2986 2423 3005 2426
rect 2986 2413 2989 2423
rect 2978 2403 2989 2406
rect 2978 2273 2981 2326
rect 2994 2323 2997 2416
rect 3002 2413 3005 2423
rect 3010 2403 3013 2566
rect 3042 2516 3045 2546
rect 3026 2513 3045 2516
rect 3050 2513 3053 2613
rect 3058 2563 3061 2596
rect 3058 2523 3061 2536
rect 3066 2533 3069 2606
rect 3082 2546 3085 2736
rect 3090 2703 3093 2736
rect 3098 2723 3101 2793
rect 3106 2786 3109 2856
rect 3114 2793 3117 2816
rect 3106 2783 3117 2786
rect 3090 2593 3093 2616
rect 3098 2603 3101 2686
rect 3106 2636 3109 2726
rect 3114 2683 3117 2783
rect 3122 2686 3125 2776
rect 3134 2766 3137 2873
rect 3150 2826 3153 2883
rect 3162 2866 3165 2933
rect 3170 2916 3173 2926
rect 3178 2923 3189 2926
rect 3194 2923 3197 2936
rect 3202 2916 3205 2936
rect 3210 2933 3213 2983
rect 3274 2946 3277 3016
rect 3234 2943 3277 2946
rect 3170 2913 3205 2916
rect 3210 2896 3213 2926
rect 3194 2893 3213 2896
rect 3162 2863 3189 2866
rect 3150 2823 3165 2826
rect 3146 2803 3149 2816
rect 3134 2763 3141 2766
rect 3130 2733 3133 2746
rect 3138 2706 3141 2763
rect 3146 2723 3149 2786
rect 3162 2733 3165 2823
rect 3178 2803 3181 2816
rect 3186 2803 3189 2863
rect 3194 2813 3197 2893
rect 3218 2886 3221 2936
rect 3234 2933 3237 2943
rect 3250 2926 3253 2936
rect 3258 2933 3269 2936
rect 3282 2933 3285 2976
rect 3298 2933 3301 2986
rect 3314 2976 3317 2996
rect 3306 2973 3317 2976
rect 3210 2883 3221 2886
rect 3202 2803 3205 2826
rect 3210 2813 3213 2883
rect 3226 2776 3229 2926
rect 3242 2913 3245 2926
rect 3250 2923 3261 2926
rect 3266 2923 3269 2933
rect 3274 2893 3277 2926
rect 3306 2923 3309 2973
rect 3314 2926 3317 2936
rect 3322 2933 3325 2946
rect 3314 2923 3325 2926
rect 3330 2916 3333 3016
rect 3362 2976 3365 3016
rect 3386 2983 3389 3016
rect 3362 2973 3373 2976
rect 3310 2913 3333 2916
rect 3234 2803 3237 2826
rect 3242 2783 3245 2806
rect 3194 2773 3229 2776
rect 3138 2703 3145 2706
rect 3122 2683 3133 2686
rect 3106 2633 3117 2636
rect 3106 2596 3109 2616
rect 3114 2603 3117 2633
rect 3130 2623 3133 2683
rect 3142 2626 3145 2703
rect 3154 2653 3181 2656
rect 3154 2633 3157 2653
rect 3142 2623 3157 2626
rect 3122 2603 3125 2616
rect 3146 2596 3149 2616
rect 3106 2593 3149 2596
rect 3074 2543 3085 2546
rect 3026 2486 3029 2513
rect 3018 2483 3029 2486
rect 3034 2486 3037 2506
rect 3034 2483 3041 2486
rect 2994 2293 2997 2316
rect 2978 2133 2981 2206
rect 2986 2186 2989 2286
rect 3002 2266 3005 2386
rect 3010 2323 3013 2336
rect 3018 2333 3021 2483
rect 3026 2383 3029 2456
rect 3038 2396 3041 2483
rect 3074 2446 3077 2543
rect 3090 2536 3093 2546
rect 3082 2533 3093 2536
rect 3090 2503 3093 2526
rect 3074 2443 3085 2446
rect 3058 2403 3061 2416
rect 3034 2393 3041 2396
rect 3034 2373 3037 2393
rect 3082 2386 3085 2443
rect 3090 2403 3093 2416
rect 3034 2323 3053 2326
rect 3026 2273 3045 2276
rect 3050 2273 3053 2316
rect 3002 2263 3037 2266
rect 3002 2203 3005 2216
rect 3026 2213 3029 2236
rect 2986 2183 2997 2186
rect 2978 2003 2981 2126
rect 2986 2123 2989 2166
rect 2994 2156 2997 2183
rect 3034 2156 3037 2263
rect 2994 2153 3005 2156
rect 3002 2123 3005 2153
rect 3010 2153 3037 2156
rect 2986 2023 2989 2116
rect 2970 1923 2973 1966
rect 2978 1933 2981 1986
rect 2986 1963 2989 2016
rect 2978 1923 2989 1926
rect 2978 1856 2981 1923
rect 2978 1853 2989 1856
rect 2938 1793 2945 1796
rect 2954 1793 2957 1806
rect 2922 1696 2925 1736
rect 2930 1703 2933 1726
rect 2938 1723 2941 1793
rect 2946 1723 2949 1746
rect 2954 1696 2957 1736
rect 2922 1693 2957 1696
rect 2922 1623 2925 1686
rect 2970 1633 2973 1826
rect 2986 1813 2989 1853
rect 2994 1823 2997 2096
rect 3002 1966 3005 2116
rect 3010 2086 3013 2153
rect 3018 2096 3021 2136
rect 3034 2133 3037 2146
rect 3018 2093 3037 2096
rect 3010 2083 3021 2086
rect 3010 1983 3013 2016
rect 3002 1963 3009 1966
rect 3006 1906 3009 1963
rect 3018 1923 3021 2083
rect 3026 2013 3029 2056
rect 3034 2003 3037 2093
rect 3042 2013 3045 2273
rect 3058 2266 3061 2376
rect 3066 2293 3069 2336
rect 3074 2333 3077 2386
rect 3082 2383 3089 2386
rect 3074 2286 3077 2326
rect 3050 2263 3061 2266
rect 3066 2283 3077 2286
rect 3026 1906 3029 1936
rect 3006 1903 3013 1906
rect 3010 1816 3013 1903
rect 3022 1903 3029 1906
rect 3022 1836 3025 1903
rect 3022 1833 3029 1836
rect 3002 1813 3013 1816
rect 3026 1813 3029 1833
rect 2978 1793 2981 1806
rect 3002 1746 3005 1813
rect 2986 1743 3005 1746
rect 2978 1723 2981 1736
rect 2898 1553 2917 1556
rect 2810 1513 2837 1516
rect 2802 1483 2829 1486
rect 2770 1433 2781 1436
rect 2742 1393 2749 1396
rect 2746 1373 2749 1393
rect 2730 1363 2741 1366
rect 2706 1093 2709 1226
rect 2714 1146 2717 1336
rect 2738 1333 2741 1363
rect 2722 1266 2725 1326
rect 2754 1283 2757 1426
rect 2762 1316 2765 1396
rect 2770 1386 2773 1433
rect 2802 1426 2805 1476
rect 2802 1423 2809 1426
rect 2778 1413 2797 1416
rect 2778 1403 2781 1413
rect 2786 1386 2789 1406
rect 2770 1383 2789 1386
rect 2770 1333 2773 1366
rect 2794 1363 2797 1406
rect 2806 1356 2809 1423
rect 2818 1393 2821 1416
rect 2802 1353 2809 1356
rect 2762 1313 2769 1316
rect 2722 1263 2757 1266
rect 2754 1203 2757 1263
rect 2714 1143 2725 1146
rect 2714 1123 2717 1136
rect 2698 1083 2717 1086
rect 2698 1013 2701 1076
rect 2706 1013 2709 1036
rect 2714 1013 2717 1083
rect 2722 1033 2725 1143
rect 2698 1003 2717 1006
rect 2666 813 2669 866
rect 2674 846 2677 896
rect 2682 856 2685 996
rect 2690 863 2693 996
rect 2698 873 2701 1003
rect 2706 893 2709 996
rect 2714 923 2717 996
rect 2722 993 2725 1026
rect 2730 1016 2733 1186
rect 2738 1023 2741 1136
rect 2754 1133 2757 1176
rect 2766 1156 2769 1313
rect 2778 1223 2781 1346
rect 2786 1323 2789 1346
rect 2794 1233 2797 1326
rect 2778 1206 2781 1216
rect 2794 1213 2797 1226
rect 2778 1203 2789 1206
rect 2766 1153 2773 1156
rect 2746 1103 2749 1126
rect 2762 1123 2765 1146
rect 2730 1013 2749 1016
rect 2738 1003 2749 1006
rect 2722 906 2725 936
rect 2718 903 2725 906
rect 2682 853 2709 856
rect 2674 843 2685 846
rect 2602 743 2629 746
rect 2562 633 2597 636
rect 2602 633 2605 736
rect 2522 583 2541 586
rect 2522 533 2525 583
rect 2530 533 2541 536
rect 2546 526 2549 606
rect 2530 523 2549 526
rect 2514 513 2541 516
rect 2530 406 2533 446
rect 2538 426 2541 513
rect 2546 436 2549 523
rect 2554 443 2557 616
rect 2562 523 2565 633
rect 2578 623 2597 626
rect 2570 583 2573 616
rect 2578 613 2581 623
rect 2594 606 2597 616
rect 2578 603 2597 606
rect 2570 533 2589 536
rect 2594 533 2597 596
rect 2602 533 2605 616
rect 2586 526 2589 533
rect 2610 526 2613 676
rect 2618 616 2621 743
rect 2626 683 2629 736
rect 2650 726 2653 736
rect 2674 733 2677 786
rect 2682 766 2685 843
rect 2706 783 2709 853
rect 2718 826 2721 903
rect 2718 823 2725 826
rect 2714 776 2717 806
rect 2706 773 2717 776
rect 2682 763 2689 766
rect 2634 633 2637 726
rect 2650 723 2677 726
rect 2626 623 2637 626
rect 2642 623 2645 676
rect 2618 613 2629 616
rect 2546 433 2565 436
rect 2538 423 2557 426
rect 2538 413 2541 423
rect 2530 403 2537 406
rect 2458 343 2485 346
rect 2450 316 2453 336
rect 2458 333 2461 343
rect 2466 323 2469 336
rect 2482 316 2485 326
rect 2450 313 2485 316
rect 2466 193 2469 206
rect 2490 133 2493 366
rect 2498 333 2501 386
rect 2522 376 2525 396
rect 2514 373 2525 376
rect 2498 206 2501 326
rect 2506 213 2509 336
rect 2514 263 2517 373
rect 2534 346 2537 403
rect 2546 383 2549 416
rect 2554 403 2557 423
rect 2562 396 2565 433
rect 2554 393 2565 396
rect 2534 343 2541 346
rect 2522 256 2525 336
rect 2514 253 2525 256
rect 2514 213 2517 253
rect 2530 243 2533 326
rect 2498 203 2517 206
rect 2490 116 2493 126
rect 2498 123 2501 166
rect 2506 123 2509 136
rect 2514 123 2517 203
rect 2538 143 2541 343
rect 2546 193 2549 356
rect 2554 316 2557 393
rect 2562 333 2565 376
rect 2570 316 2573 486
rect 2578 403 2581 526
rect 2586 523 2613 526
rect 2594 503 2597 516
rect 2602 483 2605 516
rect 2618 513 2621 556
rect 2594 403 2597 446
rect 2618 396 2621 416
rect 2610 393 2621 396
rect 2578 333 2581 356
rect 2594 333 2597 366
rect 2610 333 2613 393
rect 2626 353 2629 613
rect 2634 603 2637 616
rect 2650 603 2653 723
rect 2658 713 2669 716
rect 2658 596 2661 713
rect 2674 703 2677 716
rect 2634 593 2661 596
rect 2634 503 2637 593
rect 2666 586 2669 696
rect 2674 593 2677 656
rect 2686 586 2689 763
rect 2698 683 2701 736
rect 2706 716 2709 773
rect 2714 723 2717 746
rect 2722 726 2725 823
rect 2730 813 2733 936
rect 2738 923 2741 1003
rect 2754 973 2757 1096
rect 2770 1093 2773 1153
rect 2762 993 2765 1056
rect 2746 926 2749 936
rect 2754 933 2773 936
rect 2746 923 2757 926
rect 2746 856 2749 916
rect 2746 853 2753 856
rect 2750 786 2753 853
rect 2762 813 2765 933
rect 2778 873 2781 1146
rect 2786 1123 2789 1203
rect 2794 1126 2797 1176
rect 2802 1146 2805 1353
rect 2810 1323 2813 1336
rect 2818 1323 2821 1386
rect 2810 1213 2813 1246
rect 2818 1203 2821 1256
rect 2826 1146 2829 1483
rect 2842 1463 2845 1526
rect 2866 1523 2893 1526
rect 2898 1516 2901 1553
rect 2878 1513 2901 1516
rect 2834 1343 2837 1446
rect 2842 1296 2845 1416
rect 2850 1393 2853 1406
rect 2858 1383 2861 1416
rect 2858 1333 2861 1366
rect 2866 1326 2869 1466
rect 2878 1436 2881 1513
rect 2906 1443 2909 1536
rect 2914 1533 2917 1546
rect 2930 1463 2933 1616
rect 2962 1613 2981 1616
rect 2986 1613 2989 1743
rect 2994 1683 2997 1726
rect 3002 1723 3005 1736
rect 3010 1723 3013 1766
rect 3018 1686 3021 1736
rect 3026 1733 3029 1806
rect 3002 1683 3021 1686
rect 2938 1586 2941 1606
rect 2954 1593 2957 1606
rect 2962 1603 2965 1613
rect 2938 1583 2961 1586
rect 2946 1483 2949 1546
rect 2958 1486 2961 1583
rect 2958 1483 2965 1486
rect 2850 1323 2869 1326
rect 2874 1433 2881 1436
rect 2850 1313 2853 1323
rect 2874 1303 2877 1433
rect 2882 1383 2885 1416
rect 2890 1403 2893 1436
rect 2890 1363 2917 1366
rect 2890 1333 2893 1363
rect 2914 1333 2917 1363
rect 2914 1313 2917 1326
rect 2842 1293 2877 1296
rect 2834 1216 2837 1236
rect 2834 1213 2845 1216
rect 2802 1143 2813 1146
rect 2818 1143 2829 1146
rect 2794 1123 2805 1126
rect 2810 1116 2813 1143
rect 2834 1136 2837 1206
rect 2842 1173 2845 1213
rect 2850 1213 2869 1216
rect 2826 1133 2837 1136
rect 2802 1113 2813 1116
rect 2802 1096 2805 1113
rect 2794 1093 2805 1096
rect 2794 1036 2797 1093
rect 2794 1033 2805 1036
rect 2786 1003 2789 1016
rect 2794 1003 2797 1016
rect 2802 996 2805 1033
rect 2794 993 2805 996
rect 2794 926 2797 993
rect 2810 986 2813 1096
rect 2818 1013 2821 1126
rect 2834 1056 2837 1126
rect 2842 1093 2845 1136
rect 2850 1063 2853 1213
rect 2858 1193 2861 1206
rect 2858 1126 2861 1136
rect 2866 1133 2869 1156
rect 2858 1123 2869 1126
rect 2874 1056 2877 1293
rect 2906 1216 2909 1226
rect 2890 1213 2909 1216
rect 2890 1203 2893 1213
rect 2914 1203 2917 1216
rect 2922 1186 2925 1456
rect 2946 1393 2949 1416
rect 2954 1376 2957 1466
rect 2934 1373 2957 1376
rect 2962 1376 2965 1483
rect 2970 1443 2973 1606
rect 3002 1603 3005 1683
rect 3034 1626 3037 1996
rect 3042 1923 3045 1936
rect 3050 1906 3053 2263
rect 3066 2253 3069 2283
rect 3074 2236 3077 2276
rect 3086 2236 3089 2383
rect 3098 2373 3101 2576
rect 3154 2556 3157 2623
rect 3106 2536 3109 2556
rect 3122 2553 3157 2556
rect 3106 2533 3113 2536
rect 3122 2533 3125 2553
rect 3110 2466 3113 2533
rect 3130 2513 3133 2546
rect 3106 2463 3113 2466
rect 3138 2466 3141 2536
rect 3146 2523 3149 2546
rect 3154 2523 3157 2553
rect 3162 2476 3165 2626
rect 3170 2593 3173 2606
rect 3170 2533 3173 2566
rect 3178 2536 3181 2653
rect 3186 2603 3189 2696
rect 3178 2533 3189 2536
rect 3186 2523 3189 2533
rect 3162 2473 3173 2476
rect 3138 2463 3153 2466
rect 3106 2346 3109 2463
rect 3138 2413 3141 2456
rect 3122 2376 3125 2386
rect 3098 2343 3109 2346
rect 3114 2373 3125 2376
rect 3098 2323 3101 2343
rect 3098 2273 3101 2316
rect 3106 2253 3109 2336
rect 3114 2333 3117 2373
rect 3130 2333 3133 2376
rect 3150 2356 3153 2463
rect 3170 2426 3173 2473
rect 3162 2423 3173 2426
rect 3150 2353 3157 2356
rect 3114 2286 3117 2326
rect 3114 2283 3141 2286
rect 3070 2233 3077 2236
rect 3082 2233 3089 2236
rect 3070 2126 3073 2233
rect 3058 2093 3061 2126
rect 3070 2123 3077 2126
rect 3074 2106 3077 2123
rect 3082 2113 3085 2233
rect 3090 2133 3093 2216
rect 3098 2213 3101 2226
rect 3098 2133 3101 2206
rect 3074 2103 3085 2106
rect 3058 1933 3061 2036
rect 3066 2033 3077 2036
rect 3066 2013 3069 2033
rect 3082 2023 3085 2103
rect 3090 2023 3093 2056
rect 3090 2006 3093 2016
rect 3074 2003 3093 2006
rect 3074 1953 3077 2003
rect 3066 1933 3069 1946
rect 3074 1943 3085 1946
rect 3042 1786 3045 1906
rect 3050 1903 3057 1906
rect 3066 1903 3069 1926
rect 3054 1836 3057 1903
rect 3074 1866 3077 1943
rect 3082 1873 3085 1936
rect 3090 1923 3093 1996
rect 3074 1863 3093 1866
rect 3054 1833 3061 1836
rect 3058 1823 3061 1833
rect 3042 1783 3053 1786
rect 3058 1783 3061 1806
rect 3082 1793 3085 1816
rect 3042 1733 3045 1746
rect 3026 1623 3037 1626
rect 3010 1566 3013 1616
rect 2978 1563 3013 1566
rect 3026 1566 3029 1623
rect 3026 1563 3037 1566
rect 2978 1456 2981 1563
rect 2986 1523 2989 1556
rect 2994 1533 3021 1536
rect 3010 1463 3013 1526
rect 3026 1523 3029 1546
rect 3034 1506 3037 1563
rect 3042 1513 3045 1616
rect 3050 1533 3053 1783
rect 3090 1776 3093 1863
rect 3066 1773 3093 1776
rect 3066 1723 3069 1773
rect 3098 1756 3101 2036
rect 3106 1933 3109 2136
rect 3114 2133 3117 2236
rect 3122 2203 3125 2226
rect 3130 2203 3133 2216
rect 3138 2136 3141 2283
rect 3146 2203 3149 2276
rect 3130 2133 3141 2136
rect 3146 2133 3149 2146
rect 3154 2133 3157 2353
rect 3162 2296 3165 2423
rect 3170 2396 3173 2406
rect 3186 2403 3189 2486
rect 3194 2433 3197 2773
rect 3210 2703 3213 2726
rect 3202 2613 3205 2696
rect 3210 2553 3213 2686
rect 3202 2526 3205 2546
rect 3210 2533 3213 2546
rect 3218 2536 3221 2606
rect 3226 2566 3229 2616
rect 3234 2586 3237 2776
rect 3250 2733 3253 2816
rect 3266 2813 3269 2856
rect 3282 2813 3285 2826
rect 3290 2806 3293 2846
rect 3258 2793 3261 2806
rect 3266 2803 3277 2806
rect 3282 2803 3293 2806
rect 3298 2803 3301 2866
rect 3310 2846 3313 2913
rect 3306 2843 3313 2846
rect 3266 2746 3269 2803
rect 3258 2743 3269 2746
rect 3242 2603 3245 2626
rect 3250 2593 3253 2726
rect 3258 2603 3261 2743
rect 3266 2723 3269 2736
rect 3282 2716 3285 2736
rect 3274 2713 3285 2716
rect 3274 2703 3277 2713
rect 3290 2703 3293 2726
rect 3298 2693 3301 2736
rect 3266 2603 3269 2686
rect 3306 2683 3309 2843
rect 3314 2813 3317 2826
rect 3234 2583 3269 2586
rect 3226 2563 3245 2566
rect 3218 2533 3229 2536
rect 3202 2523 3209 2526
rect 3206 2436 3209 2523
rect 3218 2466 3221 2526
rect 3226 2476 3229 2533
rect 3234 2513 3237 2536
rect 3242 2513 3245 2563
rect 3226 2473 3245 2476
rect 3218 2463 3237 2466
rect 3206 2433 3213 2436
rect 3170 2393 3197 2396
rect 3170 2316 3173 2393
rect 3178 2353 3181 2386
rect 3194 2376 3197 2393
rect 3202 2383 3205 2416
rect 3210 2403 3213 2433
rect 3218 2413 3221 2456
rect 3218 2403 3229 2406
rect 3194 2373 3213 2376
rect 3178 2323 3181 2336
rect 3170 2313 3181 2316
rect 3162 2293 3169 2296
rect 3166 2226 3169 2293
rect 3162 2223 3169 2226
rect 3114 2003 3117 2036
rect 3106 1903 3109 1926
rect 3106 1776 3109 1876
rect 3114 1856 3117 1926
rect 3122 1873 3125 2126
rect 3130 2046 3133 2133
rect 3138 2103 3141 2126
rect 3162 2116 3165 2223
rect 3170 2163 3173 2206
rect 3154 2113 3165 2116
rect 3130 2043 3141 2046
rect 3130 2013 3133 2036
rect 3130 1946 3133 2006
rect 3138 1993 3141 2043
rect 3146 1993 3149 2036
rect 3130 1943 3149 1946
rect 3154 1943 3157 2113
rect 3170 2093 3173 2126
rect 3178 2076 3181 2313
rect 3194 2273 3197 2336
rect 3210 2323 3213 2373
rect 3218 2343 3221 2403
rect 3234 2356 3237 2463
rect 3226 2353 3237 2356
rect 3226 2323 3229 2353
rect 3234 2333 3237 2346
rect 3194 2203 3197 2216
rect 3218 2213 3221 2226
rect 3186 2096 3189 2176
rect 3194 2143 3197 2196
rect 3194 2113 3197 2136
rect 3202 2133 3205 2146
rect 3210 2133 3213 2196
rect 3226 2156 3229 2306
rect 3234 2273 3237 2326
rect 3234 2223 3237 2246
rect 3218 2153 3229 2156
rect 3186 2093 3193 2096
rect 3170 2073 3181 2076
rect 3170 2043 3173 2073
rect 3162 1946 3165 2006
rect 3170 1993 3173 2036
rect 3178 2013 3181 2066
rect 3190 2006 3193 2093
rect 3186 2003 3193 2006
rect 3162 1943 3173 1946
rect 3186 1943 3189 2003
rect 3146 1936 3149 1943
rect 3114 1853 3125 1856
rect 3106 1773 3117 1776
rect 3082 1753 3101 1756
rect 3074 1743 3109 1746
rect 3066 1703 3069 1716
rect 3058 1603 3061 1616
rect 3058 1513 3061 1546
rect 3030 1503 3037 1506
rect 2978 1453 3021 1456
rect 2962 1373 2981 1376
rect 2934 1236 2937 1373
rect 2802 983 2813 986
rect 2802 933 2805 983
rect 2818 973 2821 996
rect 2786 883 2789 926
rect 2794 923 2801 926
rect 2778 806 2781 846
rect 2798 826 2801 923
rect 2810 903 2813 926
rect 2826 913 2829 1056
rect 2834 1053 2877 1056
rect 2874 1036 2877 1053
rect 2890 1183 2925 1186
rect 2930 1233 2937 1236
rect 2890 1046 2893 1183
rect 2914 1093 2917 1126
rect 2890 1043 2897 1046
rect 2874 1033 2885 1036
rect 2834 1003 2837 1016
rect 2810 833 2813 876
rect 2786 813 2789 826
rect 2798 823 2805 826
rect 2778 803 2797 806
rect 2746 783 2753 786
rect 2746 763 2749 783
rect 2746 743 2781 746
rect 2746 733 2749 743
rect 2722 723 2749 726
rect 2706 713 2717 716
rect 2642 533 2645 586
rect 2650 583 2669 586
rect 2682 583 2689 586
rect 2698 596 2701 616
rect 2706 603 2709 626
rect 2714 613 2717 713
rect 2746 666 2749 723
rect 2754 693 2757 736
rect 2762 683 2765 736
rect 2746 663 2757 666
rect 2722 596 2725 616
rect 2698 593 2725 596
rect 2642 423 2645 526
rect 2650 516 2653 583
rect 2658 523 2661 556
rect 2682 546 2685 583
rect 2698 566 2701 593
rect 2730 576 2733 616
rect 2738 613 2741 626
rect 2666 543 2685 546
rect 2690 563 2701 566
rect 2706 573 2733 576
rect 2706 563 2709 573
rect 2666 533 2669 543
rect 2674 526 2677 536
rect 2666 523 2677 526
rect 2650 513 2661 516
rect 2658 453 2661 513
rect 2666 426 2669 523
rect 2674 503 2677 516
rect 2682 493 2685 536
rect 2690 463 2693 563
rect 2730 556 2733 566
rect 2698 553 2733 556
rect 2698 523 2701 553
rect 2706 533 2717 536
rect 2722 533 2725 546
rect 2662 423 2669 426
rect 2554 313 2561 316
rect 2570 313 2581 316
rect 2558 236 2561 313
rect 2578 266 2581 313
rect 2594 303 2597 326
rect 2570 263 2581 266
rect 2570 243 2573 263
rect 2602 253 2605 326
rect 2618 323 2621 336
rect 2626 303 2629 336
rect 2634 323 2637 416
rect 2642 306 2645 366
rect 2662 346 2665 423
rect 2674 353 2677 416
rect 2690 403 2693 426
rect 2698 413 2701 476
rect 2714 436 2717 526
rect 2706 433 2717 436
rect 2638 303 2645 306
rect 2650 343 2665 346
rect 2650 306 2653 343
rect 2658 316 2661 336
rect 2674 333 2685 336
rect 2658 313 2677 316
rect 2650 303 2661 306
rect 2554 233 2561 236
rect 2554 216 2557 233
rect 2554 213 2573 216
rect 2578 203 2581 216
rect 2610 203 2613 216
rect 2626 213 2629 246
rect 2638 236 2641 303
rect 2638 233 2645 236
rect 2642 213 2645 233
rect 2618 166 2621 206
rect 2650 186 2653 286
rect 2658 203 2661 303
rect 2666 206 2669 246
rect 2674 213 2677 313
rect 2682 206 2685 326
rect 2690 276 2693 376
rect 2698 303 2701 336
rect 2706 283 2709 433
rect 2722 353 2725 526
rect 2730 523 2733 553
rect 2738 493 2741 606
rect 2746 523 2749 656
rect 2754 596 2757 663
rect 2762 603 2765 676
rect 2770 613 2773 736
rect 2778 683 2781 743
rect 2786 733 2789 786
rect 2794 706 2797 803
rect 2802 713 2805 823
rect 2810 803 2813 826
rect 2818 733 2821 896
rect 2826 813 2829 846
rect 2826 763 2829 806
rect 2834 746 2837 936
rect 2842 913 2845 1016
rect 2842 813 2845 906
rect 2850 803 2853 1006
rect 2858 916 2861 1026
rect 2866 973 2869 996
rect 2874 923 2877 986
rect 2882 923 2885 1033
rect 2894 986 2897 1043
rect 2922 1026 2925 1176
rect 2930 1083 2933 1233
rect 2906 1023 2933 1026
rect 2906 1013 2909 1023
rect 2890 983 2897 986
rect 2858 913 2877 916
rect 2834 743 2845 746
rect 2794 703 2813 706
rect 2786 613 2789 626
rect 2778 596 2781 606
rect 2794 603 2797 646
rect 2810 616 2813 703
rect 2810 613 2821 616
rect 2754 593 2773 596
rect 2778 593 2805 596
rect 2722 313 2725 336
rect 2746 323 2749 336
rect 2690 273 2709 276
rect 2666 203 2685 206
rect 2690 203 2701 206
rect 2706 203 2709 273
rect 2754 226 2757 586
rect 2762 473 2765 536
rect 2770 463 2773 593
rect 2802 566 2805 586
rect 2778 456 2781 536
rect 2794 533 2797 566
rect 2802 563 2813 566
rect 2802 533 2805 563
rect 2770 453 2781 456
rect 2770 413 2773 453
rect 2786 423 2789 526
rect 2794 406 2797 466
rect 2802 413 2805 526
rect 2810 433 2813 516
rect 2790 403 2797 406
rect 2770 286 2773 356
rect 2770 283 2781 286
rect 2778 236 2781 283
rect 2790 256 2793 403
rect 2790 253 2797 256
rect 2778 233 2785 236
rect 2730 223 2765 226
rect 2730 213 2733 223
rect 2738 203 2741 216
rect 2650 183 2661 186
rect 2602 163 2621 166
rect 2522 116 2525 136
rect 2554 123 2557 136
rect 2602 123 2605 163
rect 2658 123 2661 183
rect 2698 163 2701 203
rect 2746 166 2749 206
rect 2754 193 2757 216
rect 2762 203 2765 223
rect 2770 203 2773 226
rect 2782 166 2785 233
rect 2794 203 2797 253
rect 2802 193 2805 406
rect 2810 373 2813 406
rect 2818 283 2821 613
rect 2826 583 2829 686
rect 2834 646 2837 676
rect 2842 653 2845 743
rect 2850 693 2853 726
rect 2834 643 2845 646
rect 2834 533 2837 616
rect 2842 613 2845 643
rect 2850 556 2853 676
rect 2858 603 2861 906
rect 2866 813 2869 866
rect 2874 786 2877 913
rect 2882 883 2885 916
rect 2890 896 2893 983
rect 2898 956 2901 966
rect 2914 963 2917 1006
rect 2922 956 2925 1016
rect 2898 953 2925 956
rect 2898 903 2901 926
rect 2906 923 2909 936
rect 2914 923 2917 953
rect 2890 893 2909 896
rect 2890 813 2893 866
rect 2882 803 2893 806
rect 2906 803 2909 893
rect 2922 863 2925 936
rect 2866 783 2901 786
rect 2898 723 2901 783
rect 2898 713 2909 716
rect 2866 613 2869 696
rect 2874 613 2877 626
rect 2890 613 2893 656
rect 2882 596 2885 606
rect 2898 603 2901 713
rect 2914 696 2917 736
rect 2906 693 2917 696
rect 2922 693 2925 726
rect 2930 716 2933 1023
rect 2938 1006 2941 1216
rect 2946 1173 2949 1256
rect 2954 1203 2957 1236
rect 2962 1166 2965 1216
rect 2970 1213 2973 1366
rect 2978 1313 2981 1373
rect 2986 1236 2989 1336
rect 2994 1243 2997 1396
rect 3002 1253 3005 1436
rect 3010 1393 3013 1406
rect 3018 1376 3021 1453
rect 3030 1436 3033 1503
rect 3030 1433 3037 1436
rect 3014 1373 3021 1376
rect 3014 1276 3017 1373
rect 3026 1323 3029 1416
rect 3026 1283 3029 1316
rect 3014 1273 3021 1276
rect 2986 1233 2997 1236
rect 2970 1186 2973 1206
rect 2970 1183 2989 1186
rect 2962 1163 2981 1166
rect 2970 1123 2973 1156
rect 2978 1133 2981 1163
rect 2938 1003 2949 1006
rect 2954 1003 2957 1026
rect 2962 983 2965 1096
rect 2986 1063 2989 1183
rect 2994 1046 2997 1233
rect 2978 1043 2997 1046
rect 2970 1003 2973 1026
rect 2978 976 2981 1043
rect 3002 1036 3005 1126
rect 3010 1063 3013 1176
rect 3018 1053 3021 1273
rect 3026 1193 3029 1216
rect 3026 1123 3029 1176
rect 3034 1103 3037 1433
rect 3042 1356 3045 1506
rect 3050 1413 3053 1506
rect 3058 1463 3061 1496
rect 3066 1486 3069 1616
rect 3074 1553 3077 1743
rect 3082 1733 3101 1736
rect 3082 1723 3093 1726
rect 3082 1686 3085 1706
rect 3090 1693 3093 1706
rect 3082 1683 3093 1686
rect 3082 1546 3085 1616
rect 3074 1543 3085 1546
rect 3090 1543 3093 1683
rect 3098 1586 3101 1733
rect 3106 1713 3109 1736
rect 3114 1726 3117 1773
rect 3122 1733 3125 1853
rect 3114 1723 3125 1726
rect 3114 1646 3117 1716
rect 3106 1643 3117 1646
rect 3122 1676 3125 1723
rect 3130 1696 3133 1936
rect 3138 1703 3141 1936
rect 3146 1933 3165 1936
rect 3146 1903 3149 1926
rect 3162 1923 3165 1933
rect 3170 1906 3173 1943
rect 3166 1903 3173 1906
rect 3146 1763 3149 1816
rect 3146 1723 3149 1756
rect 3154 1746 3157 1896
rect 3166 1806 3169 1903
rect 3178 1893 3181 1936
rect 3194 1933 3197 1946
rect 3186 1886 3189 1926
rect 3162 1803 3169 1806
rect 3178 1883 3189 1886
rect 3178 1803 3181 1883
rect 3186 1813 3189 1856
rect 3162 1786 3165 1803
rect 3170 1793 3189 1796
rect 3162 1783 3173 1786
rect 3154 1743 3165 1746
rect 3154 1696 3157 1736
rect 3130 1693 3157 1696
rect 3122 1673 3157 1676
rect 3106 1596 3109 1643
rect 3114 1603 3117 1636
rect 3122 1613 3125 1673
rect 3122 1603 3133 1606
rect 3138 1603 3141 1616
rect 3106 1593 3133 1596
rect 3098 1583 3117 1586
rect 3074 1493 3077 1543
rect 3066 1483 3077 1486
rect 3066 1413 3069 1446
rect 3042 1353 3061 1356
rect 3042 1323 3045 1336
rect 3050 1253 3053 1346
rect 3058 1333 3061 1353
rect 3058 1323 3069 1326
rect 3042 1173 3045 1246
rect 3058 1176 3061 1246
rect 3050 1173 3061 1176
rect 3042 1086 3045 1146
rect 3026 1083 3045 1086
rect 2986 983 2989 1016
rect 2954 973 2981 976
rect 2994 976 2997 1036
rect 3002 1033 3021 1036
rect 3002 993 3005 1026
rect 3010 1003 3013 1026
rect 2994 973 3001 976
rect 2938 896 2941 926
rect 2954 923 2957 973
rect 2938 893 2945 896
rect 2942 836 2945 893
rect 2938 833 2945 836
rect 2938 813 2941 833
rect 2954 783 2957 906
rect 2978 903 2981 936
rect 2986 923 2989 966
rect 2998 916 3001 973
rect 2994 913 3001 916
rect 2938 773 2965 776
rect 2938 733 2941 773
rect 2962 743 2965 773
rect 2930 713 2937 716
rect 2882 593 2909 596
rect 2914 586 2917 646
rect 2842 553 2853 556
rect 2842 533 2845 553
rect 2858 533 2861 546
rect 2834 523 2845 526
rect 2850 516 2853 526
rect 2834 513 2861 516
rect 2834 446 2837 513
rect 2866 473 2869 586
rect 2874 446 2877 526
rect 2826 443 2837 446
rect 2866 443 2877 446
rect 2826 303 2829 443
rect 2834 413 2837 426
rect 2850 386 2853 406
rect 2858 403 2861 416
rect 2866 393 2869 443
rect 2874 403 2877 436
rect 2882 413 2885 586
rect 2890 583 2917 586
rect 2890 523 2893 583
rect 2922 576 2925 656
rect 2934 636 2937 713
rect 2914 573 2925 576
rect 2930 633 2937 636
rect 2898 513 2901 536
rect 2906 533 2909 566
rect 2882 393 2885 406
rect 2850 383 2877 386
rect 2850 313 2853 336
rect 2874 323 2877 383
rect 2882 286 2885 376
rect 2874 283 2885 286
rect 2810 213 2813 226
rect 2826 213 2829 236
rect 2874 226 2877 283
rect 2874 223 2885 226
rect 2738 163 2749 166
rect 2690 123 2693 146
rect 2738 123 2741 163
rect 2770 123 2773 166
rect 2778 163 2785 166
rect 2778 143 2781 163
rect 2794 133 2797 156
rect 2818 123 2821 206
rect 2858 203 2877 206
rect 2882 203 2885 223
rect 2890 213 2893 436
rect 2898 403 2901 446
rect 2906 366 2909 466
rect 2898 363 2909 366
rect 2914 366 2917 573
rect 2922 493 2925 566
rect 2930 463 2933 633
rect 2938 576 2941 616
rect 2946 583 2949 726
rect 2962 713 2965 736
rect 2954 613 2957 686
rect 2954 586 2957 606
rect 2962 603 2965 656
rect 2970 613 2973 866
rect 2978 756 2981 846
rect 2986 763 2989 816
rect 2994 796 2997 913
rect 3018 886 3021 1033
rect 3010 883 3021 886
rect 3010 823 3013 883
rect 3026 876 3029 1083
rect 3034 1013 3037 1046
rect 3034 923 3037 1006
rect 3050 1003 3053 1173
rect 3066 1166 3069 1236
rect 3074 1173 3077 1483
rect 3082 1393 3085 1536
rect 3098 1526 3101 1536
rect 3090 1523 3101 1526
rect 3090 1493 3093 1523
rect 3098 1486 3101 1516
rect 3090 1483 3101 1486
rect 3082 1333 3085 1366
rect 3090 1323 3093 1483
rect 3098 1386 3101 1466
rect 3106 1456 3109 1526
rect 3114 1463 3117 1583
rect 3122 1503 3125 1576
rect 3130 1513 3133 1593
rect 3106 1453 3117 1456
rect 3106 1393 3109 1446
rect 3098 1383 3109 1386
rect 3082 1213 3085 1226
rect 3090 1213 3093 1316
rect 3106 1313 3109 1383
rect 3114 1266 3117 1453
rect 3106 1263 3117 1266
rect 3098 1203 3101 1216
rect 3106 1176 3109 1263
rect 3090 1173 3109 1176
rect 3058 1163 3069 1166
rect 3058 1143 3061 1163
rect 3058 1133 3084 1136
rect 3058 1123 3061 1133
rect 3066 1046 3069 1126
rect 3074 1086 3077 1126
rect 3090 1096 3093 1173
rect 3098 1133 3101 1156
rect 3090 1093 3101 1096
rect 3074 1083 3085 1086
rect 3066 1043 3077 1046
rect 3066 1016 3069 1036
rect 3058 1013 3069 1016
rect 3042 923 3045 986
rect 3066 946 3069 1006
rect 3074 1003 3077 1043
rect 3082 1013 3085 1083
rect 3090 1046 3093 1086
rect 3098 1066 3101 1093
rect 3106 1076 3109 1136
rect 3114 1083 3117 1256
rect 3122 1086 3125 1496
rect 3130 1413 3133 1496
rect 3130 1393 3133 1406
rect 3138 1386 3141 1546
rect 3146 1533 3149 1666
rect 3154 1613 3157 1673
rect 3154 1573 3157 1606
rect 3154 1513 3157 1536
rect 3146 1433 3149 1506
rect 3162 1496 3165 1743
rect 3170 1723 3173 1783
rect 3170 1563 3173 1666
rect 3158 1493 3165 1496
rect 3170 1493 3173 1526
rect 3146 1403 3149 1416
rect 3158 1406 3161 1493
rect 3170 1413 3173 1466
rect 3158 1403 3165 1406
rect 3138 1383 3145 1386
rect 3162 1383 3165 1403
rect 3130 1243 3133 1346
rect 3142 1326 3145 1383
rect 3170 1363 3173 1406
rect 3154 1343 3173 1346
rect 3154 1333 3157 1343
rect 3142 1323 3157 1326
rect 3138 1223 3141 1316
rect 3146 1203 3149 1256
rect 3130 1116 3133 1176
rect 3146 1163 3149 1196
rect 3154 1193 3157 1323
rect 3162 1173 3165 1336
rect 3170 1323 3173 1343
rect 3178 1333 3181 1736
rect 3186 1693 3189 1726
rect 3194 1676 3197 1876
rect 3202 1733 3205 2096
rect 3210 2033 3213 2126
rect 3218 2046 3221 2153
rect 3226 2143 3237 2146
rect 3226 2063 3229 2143
rect 3218 2043 3237 2046
rect 3210 1946 3213 2016
rect 3218 1993 3221 2006
rect 3210 1943 3221 1946
rect 3210 1903 3213 1936
rect 3218 1933 3221 1943
rect 3218 1866 3221 1926
rect 3210 1863 3221 1866
rect 3210 1823 3213 1863
rect 3202 1723 3213 1726
rect 3218 1723 3221 1856
rect 3226 1706 3229 2016
rect 3234 1793 3237 2043
rect 3242 2003 3245 2473
rect 3250 2403 3253 2546
rect 3258 2413 3261 2456
rect 3258 2366 3261 2386
rect 3266 2373 3269 2583
rect 3274 2563 3277 2616
rect 3282 2593 3285 2606
rect 3290 2573 3293 2616
rect 3314 2613 3317 2806
rect 3330 2796 3333 2816
rect 3326 2793 3333 2796
rect 3326 2736 3329 2793
rect 3338 2753 3341 2806
rect 3346 2786 3349 2946
rect 3370 2843 3373 2973
rect 3442 2943 3445 3016
rect 3466 2993 3469 3006
rect 3490 2996 3493 3016
rect 3482 2993 3493 2996
rect 3482 2936 3485 2993
rect 3546 2976 3549 3016
rect 3570 2993 3573 3006
rect 3498 2973 3549 2976
rect 3354 2803 3357 2826
rect 3378 2796 3381 2816
rect 3386 2813 3389 2896
rect 3386 2803 3397 2806
rect 3402 2803 3405 2926
rect 3418 2876 3421 2896
rect 3418 2873 3425 2876
rect 3410 2813 3413 2856
rect 3422 2816 3425 2873
rect 3450 2856 3453 2926
rect 3458 2903 3461 2936
rect 3466 2923 3469 2936
rect 3474 2933 3485 2936
rect 3490 2926 3493 2936
rect 3498 2933 3501 2973
rect 3482 2883 3485 2926
rect 3490 2923 3501 2926
rect 3506 2916 3509 2936
rect 3498 2913 3509 2916
rect 3434 2853 3453 2856
rect 3434 2823 3437 2853
rect 3422 2813 3429 2816
rect 3418 2796 3421 2806
rect 3378 2793 3421 2796
rect 3346 2783 3353 2786
rect 3418 2783 3421 2793
rect 3322 2733 3329 2736
rect 3322 2713 3325 2733
rect 3330 2723 3341 2726
rect 3350 2716 3353 2783
rect 3378 2743 3413 2746
rect 3378 2733 3381 2743
rect 3346 2713 3353 2716
rect 3338 2693 3341 2706
rect 3346 2676 3349 2713
rect 3338 2673 3349 2676
rect 3306 2533 3309 2596
rect 3322 2566 3325 2626
rect 3338 2586 3341 2673
rect 3354 2613 3357 2696
rect 3362 2623 3365 2716
rect 3370 2693 3373 2726
rect 3378 2723 3389 2726
rect 3394 2626 3397 2736
rect 3402 2683 3405 2726
rect 3410 2643 3413 2743
rect 3418 2723 3421 2736
rect 3426 2626 3429 2813
rect 3450 2786 3453 2846
rect 3442 2783 3453 2786
rect 3394 2623 3405 2626
rect 3338 2583 3349 2586
rect 3314 2563 3325 2566
rect 3282 2486 3285 2496
rect 3274 2483 3285 2486
rect 3274 2403 3277 2483
rect 3282 2386 3285 2436
rect 3290 2403 3293 2526
rect 3298 2413 3301 2516
rect 3314 2486 3317 2563
rect 3314 2483 3321 2486
rect 3306 2403 3309 2456
rect 3318 2426 3321 2483
rect 3318 2423 3325 2426
rect 3274 2383 3285 2386
rect 3258 2363 3269 2366
rect 3250 2256 3253 2336
rect 3258 2323 3261 2336
rect 3266 2333 3269 2363
rect 3274 2273 3277 2383
rect 3314 2376 3317 2406
rect 3282 2373 3317 2376
rect 3282 2333 3285 2373
rect 3322 2366 3325 2423
rect 3290 2363 3325 2366
rect 3290 2326 3293 2363
rect 3286 2323 3293 2326
rect 3286 2266 3289 2323
rect 3282 2263 3289 2266
rect 3250 2253 3261 2256
rect 3258 2203 3261 2253
rect 3250 2123 3253 2156
rect 3258 2133 3261 2146
rect 3266 2126 3269 2166
rect 3274 2133 3277 2216
rect 3266 2123 3277 2126
rect 3282 2123 3285 2263
rect 3290 2193 3293 2246
rect 3298 2186 3301 2326
rect 3290 2183 3301 2186
rect 3290 2126 3293 2183
rect 3298 2133 3301 2176
rect 3290 2123 3301 2126
rect 3250 2013 3253 2026
rect 3242 1933 3245 1966
rect 3250 1933 3253 1946
rect 3242 1863 3245 1926
rect 3242 1803 3245 1816
rect 3250 1796 3253 1926
rect 3258 1853 3261 2036
rect 3266 1933 3269 2116
rect 3266 1903 3269 1926
rect 3274 1906 3277 2123
rect 3306 2116 3309 2256
rect 3314 2243 3317 2336
rect 3322 2263 3325 2326
rect 3330 2236 3333 2566
rect 3338 2243 3341 2556
rect 3346 2333 3349 2583
rect 3354 2553 3357 2606
rect 3354 2523 3357 2546
rect 3354 2403 3357 2486
rect 3362 2406 3365 2606
rect 3370 2476 3373 2596
rect 3378 2563 3381 2596
rect 3386 2533 3389 2606
rect 3394 2593 3397 2616
rect 3402 2573 3405 2623
rect 3410 2616 3413 2626
rect 3426 2623 3433 2626
rect 3410 2613 3421 2616
rect 3370 2473 3381 2476
rect 3378 2426 3381 2473
rect 3410 2433 3413 2606
rect 3378 2423 3389 2426
rect 3362 2403 3369 2406
rect 3354 2333 3357 2376
rect 3366 2346 3369 2403
rect 3378 2356 3381 2416
rect 3386 2403 3389 2423
rect 3394 2413 3413 2416
rect 3394 2403 3405 2406
rect 3402 2393 3413 2396
rect 3378 2353 3397 2356
rect 3362 2343 3369 2346
rect 3362 2316 3365 2343
rect 3378 2333 3381 2346
rect 3358 2313 3365 2316
rect 3330 2233 3341 2236
rect 3314 2213 3317 2226
rect 3322 2223 3333 2226
rect 3314 2153 3317 2206
rect 3322 2173 3325 2223
rect 3338 2216 3341 2233
rect 3330 2213 3341 2216
rect 3282 2113 3309 2116
rect 3282 1956 3285 2113
rect 3290 2023 3293 2086
rect 3306 2013 3309 2086
rect 3314 2043 3317 2136
rect 3322 2113 3325 2126
rect 3330 2096 3333 2213
rect 3338 2173 3341 2206
rect 3346 2156 3349 2266
rect 3358 2236 3361 2313
rect 3370 2266 3373 2326
rect 3386 2273 3389 2336
rect 3394 2333 3397 2353
rect 3402 2266 3405 2393
rect 3410 2366 3413 2386
rect 3418 2376 3421 2613
rect 3430 2546 3433 2623
rect 3442 2603 3445 2783
rect 3450 2733 3453 2776
rect 3458 2703 3461 2726
rect 3466 2623 3469 2726
rect 3474 2683 3477 2816
rect 3482 2773 3485 2816
rect 3490 2766 3493 2806
rect 3482 2763 3493 2766
rect 3482 2693 3485 2763
rect 3498 2713 3501 2913
rect 3514 2736 3517 2973
rect 3554 2966 3557 2986
rect 3522 2933 3525 2966
rect 3546 2963 3557 2966
rect 3530 2923 3533 2936
rect 3538 2933 3541 2946
rect 3546 2923 3549 2963
rect 3554 2926 3557 2936
rect 3562 2933 3589 2936
rect 3602 2933 3605 2996
rect 3618 2983 3621 3016
rect 3650 2966 3653 3016
rect 3682 3013 3685 3126
rect 3690 3023 3725 3026
rect 3690 3013 3693 3023
rect 3682 3003 3693 3006
rect 3642 2963 3653 2966
rect 3554 2923 3565 2926
rect 3586 2906 3589 2933
rect 3626 2923 3629 2946
rect 3642 2906 3645 2963
rect 3586 2903 3597 2906
rect 3642 2903 3653 2906
rect 3522 2786 3525 2826
rect 3530 2796 3533 2866
rect 3546 2823 3581 2826
rect 3538 2803 3541 2816
rect 3546 2813 3549 2823
rect 3530 2793 3541 2796
rect 3522 2783 3549 2786
rect 3506 2733 3517 2736
rect 3538 2733 3541 2776
rect 3546 2733 3549 2783
rect 3562 2746 3565 2816
rect 3570 2753 3573 2806
rect 3578 2793 3581 2823
rect 3586 2786 3589 2903
rect 3650 2886 3653 2903
rect 3674 2896 3677 2996
rect 3690 2936 3693 2996
rect 3698 2943 3701 3016
rect 3706 2983 3709 3006
rect 3714 2956 3717 3016
rect 3722 3003 3725 3023
rect 3730 2993 3733 3126
rect 3778 3123 3781 3186
rect 3786 3066 3789 3126
rect 3794 3113 3797 3213
rect 3818 3203 3821 3216
rect 3826 3203 3829 3353
rect 3834 3243 3837 3316
rect 3842 3253 3845 3346
rect 3850 3326 3853 3336
rect 3866 3333 3869 3346
rect 3874 3333 3877 3366
rect 3850 3323 3869 3326
rect 3882 3293 3885 3403
rect 3890 3333 3893 3516
rect 3906 3513 3917 3516
rect 3898 3403 3901 3446
rect 3890 3313 3893 3326
rect 3850 3223 3853 3246
rect 3882 3213 3893 3216
rect 3850 3193 3853 3206
rect 3898 3203 3901 3326
rect 3906 3296 3909 3513
rect 3922 3503 3925 3573
rect 3954 3536 3957 3916
rect 3966 3906 3969 4023
rect 3978 3916 3981 4033
rect 3986 4023 3989 4043
rect 3986 3923 3989 3996
rect 3994 3986 3997 4103
rect 4010 4076 4013 4123
rect 4018 4103 4021 4126
rect 4026 4083 4029 4133
rect 4066 4126 4069 4136
rect 4010 4073 4021 4076
rect 4018 4043 4021 4073
rect 4002 4013 4005 4036
rect 4002 3996 4005 4006
rect 4010 4003 4021 4006
rect 4002 3993 4013 3996
rect 3994 3983 4005 3986
rect 3994 3933 3997 3946
rect 4002 3923 4005 3983
rect 4010 3963 4013 3993
rect 3978 3913 4005 3916
rect 3966 3903 3973 3906
rect 3962 3793 3965 3816
rect 3970 3693 3973 3903
rect 3978 3813 3981 3846
rect 3994 3813 3997 3856
rect 4002 3806 4005 3913
rect 3962 3563 3965 3666
rect 3946 3533 3957 3536
rect 3914 3393 3917 3416
rect 3922 3403 3925 3496
rect 3938 3413 3941 3446
rect 3946 3436 3949 3533
rect 3954 3516 3957 3526
rect 3962 3523 3965 3546
rect 3970 3533 3973 3616
rect 3978 3613 3981 3806
rect 3986 3783 3989 3806
rect 3994 3803 4005 3806
rect 4010 3796 4013 3936
rect 4018 3846 4021 3986
rect 4026 3866 4029 4026
rect 4034 3913 4037 4126
rect 4042 4103 4045 4126
rect 4050 4113 4053 4126
rect 4058 4123 4069 4126
rect 4042 3923 4045 3966
rect 4050 3906 4053 4086
rect 4058 4013 4061 4123
rect 4066 4093 4069 4116
rect 4046 3903 4053 3906
rect 4026 3863 4037 3866
rect 4018 3843 4029 3846
rect 4002 3793 4013 3796
rect 3986 3723 3989 3776
rect 4002 3736 4005 3793
rect 4018 3773 4021 3836
rect 4026 3776 4029 3843
rect 4034 3813 4037 3863
rect 4046 3836 4049 3903
rect 4058 3886 4061 3966
rect 4074 3956 4077 4136
rect 4082 4073 4085 4126
rect 4090 4003 4093 4143
rect 4098 4126 4101 4153
rect 4114 4146 4117 4176
rect 4106 4143 4117 4146
rect 4106 4133 4109 4143
rect 4098 4123 4109 4126
rect 4098 4103 4101 4116
rect 4098 4013 4101 4036
rect 4082 3963 4085 3996
rect 4074 3953 4085 3956
rect 4066 3933 4069 3946
rect 4074 3933 4077 3946
rect 4074 3893 4077 3926
rect 4058 3883 4077 3886
rect 4046 3833 4053 3836
rect 4050 3813 4053 3833
rect 4042 3793 4045 3806
rect 4058 3803 4061 3866
rect 4066 3796 4069 3846
rect 4074 3803 4077 3883
rect 4082 3863 4085 3953
rect 4090 3933 4093 3976
rect 4090 3913 4093 3926
rect 4066 3793 4077 3796
rect 4026 3773 4037 3776
rect 4010 3743 4061 3746
rect 3994 3703 3997 3736
rect 4002 3733 4037 3736
rect 4058 3733 4061 3743
rect 4066 3733 4069 3786
rect 4074 3733 4077 3793
rect 4034 3673 4037 3733
rect 4042 3703 4045 3726
rect 4050 3713 4053 3726
rect 3994 3606 3997 3636
rect 4018 3623 4045 3626
rect 4002 3613 4013 3616
rect 3994 3603 4005 3606
rect 3978 3523 3981 3586
rect 3986 3516 3989 3536
rect 3954 3513 3989 3516
rect 3994 3513 3997 3536
rect 4002 3473 4005 3603
rect 4018 3586 4021 3623
rect 4014 3583 4021 3586
rect 4034 3586 4037 3616
rect 4042 3613 4045 3623
rect 4042 3593 4045 3606
rect 4034 3583 4045 3586
rect 4014 3516 4017 3583
rect 4050 3566 4053 3696
rect 4066 3683 4069 3726
rect 4082 3713 4085 3856
rect 4098 3843 4101 3946
rect 4106 3933 4109 4123
rect 4114 4013 4117 4136
rect 4122 4093 4125 4186
rect 4150 4176 4153 4223
rect 4138 4156 4141 4176
rect 4150 4173 4157 4176
rect 4138 4153 4149 4156
rect 4146 4143 4149 4153
rect 4122 4013 4125 4046
rect 4114 3933 4117 4006
rect 4130 4003 4133 4136
rect 4138 4103 4141 4126
rect 4146 4076 4149 4136
rect 4154 4083 4157 4173
rect 4162 4133 4165 4216
rect 4178 4193 4181 4206
rect 4202 4176 4205 4216
rect 4258 4213 4261 4340
rect 4170 4173 4205 4176
rect 4170 4133 4173 4173
rect 4210 4143 4253 4146
rect 4162 4076 4165 4126
rect 4146 4073 4165 4076
rect 4138 4016 4141 4046
rect 4138 4013 4149 4016
rect 4114 3913 4117 3926
rect 4098 3813 4101 3826
rect 4090 3796 4093 3806
rect 4098 3803 4109 3806
rect 4114 3803 4117 3876
rect 4122 3796 4125 3996
rect 4130 3826 4133 3946
rect 4138 3873 4141 4006
rect 4146 3913 4149 4013
rect 4154 3843 4157 4016
rect 4162 3933 4165 3986
rect 4170 3923 4173 4126
rect 4178 4116 4181 4136
rect 4178 4113 4189 4116
rect 4202 4113 4205 4136
rect 4210 4133 4213 4143
rect 4186 4056 4189 4113
rect 4182 4053 4189 4056
rect 4182 3966 4185 4053
rect 4194 4023 4197 4036
rect 4194 3983 4197 4006
rect 4182 3963 4189 3966
rect 4178 3906 4181 3956
rect 4174 3903 4181 3906
rect 4130 3823 4141 3826
rect 4130 3803 4133 3816
rect 4090 3793 4117 3796
rect 4122 3793 4133 3796
rect 4058 3603 4061 3626
rect 4066 3613 4085 3616
rect 4066 3586 4069 3606
rect 4030 3563 4053 3566
rect 4058 3583 4069 3586
rect 4074 3583 4077 3606
rect 4090 3603 4093 3736
rect 4098 3586 4101 3736
rect 4106 3643 4109 3776
rect 4114 3733 4117 3746
rect 4130 3733 4133 3793
rect 4122 3683 4125 3726
rect 4138 3713 4141 3823
rect 4146 3686 4149 3836
rect 4154 3806 4157 3816
rect 4162 3813 4165 3886
rect 4174 3836 4177 3903
rect 4174 3833 4181 3836
rect 4154 3803 4173 3806
rect 4178 3756 4181 3833
rect 4170 3753 4181 3756
rect 4154 3696 4157 3726
rect 4162 3703 4165 3736
rect 4154 3693 4165 3696
rect 4146 3683 4157 3686
rect 4138 3613 4141 3626
rect 4098 3583 4109 3586
rect 4014 3513 4021 3516
rect 4018 3493 4021 3513
rect 4030 3506 4033 3563
rect 4058 3556 4061 3583
rect 4050 3553 4061 3556
rect 4042 3523 4045 3536
rect 4026 3503 4033 3506
rect 4026 3486 4029 3503
rect 4010 3483 4029 3486
rect 3946 3433 3973 3436
rect 3946 3423 3965 3426
rect 3946 3406 3949 3423
rect 3922 3343 3925 3396
rect 3930 3393 3933 3406
rect 3938 3403 3949 3406
rect 3938 3383 3941 3403
rect 3954 3396 3957 3416
rect 3962 3413 3965 3423
rect 3970 3406 3973 3433
rect 3962 3403 3973 3406
rect 3978 3403 3981 3426
rect 3986 3413 4005 3416
rect 4010 3406 4013 3483
rect 4018 3456 4021 3476
rect 4018 3453 4025 3456
rect 4050 3453 4053 3553
rect 4058 3523 4061 3546
rect 3994 3396 3997 3406
rect 4002 3403 4013 3406
rect 3954 3393 3997 3396
rect 4010 3336 4013 3386
rect 4022 3356 4025 3453
rect 4042 3376 4045 3406
rect 4066 3376 4069 3576
rect 4074 3503 4077 3526
rect 4082 3513 4085 3536
rect 4098 3533 4101 3546
rect 4106 3533 4109 3583
rect 4114 3573 4117 3606
rect 4146 3596 4149 3676
rect 4130 3593 4149 3596
rect 4090 3523 4109 3526
rect 4074 3413 4077 3426
rect 4042 3373 4069 3376
rect 4090 3376 4093 3456
rect 4090 3373 4101 3376
rect 3906 3293 3913 3296
rect 3910 3236 3913 3293
rect 3922 3243 3925 3336
rect 4002 3333 4013 3336
rect 4018 3353 4025 3356
rect 4018 3336 4021 3353
rect 4018 3333 4029 3336
rect 3906 3233 3913 3236
rect 3858 3153 3861 3196
rect 3890 3173 3893 3196
rect 3802 3133 3805 3146
rect 3818 3123 3821 3136
rect 3786 3063 3805 3066
rect 3754 3023 3789 3026
rect 3754 3013 3757 3023
rect 3746 3003 3757 3006
rect 3762 2993 3765 3016
rect 3770 3003 3773 3016
rect 3706 2953 3717 2956
rect 3682 2933 3693 2936
rect 3682 2903 3685 2926
rect 3674 2893 3685 2896
rect 3690 2893 3693 2926
rect 3602 2883 3653 2886
rect 3602 2826 3605 2883
rect 3578 2783 3589 2786
rect 3598 2823 3605 2826
rect 3554 2743 3565 2746
rect 3506 2696 3509 2733
rect 3498 2693 3509 2696
rect 3450 2563 3453 2606
rect 3458 2546 3461 2606
rect 3466 2553 3469 2616
rect 3426 2543 3433 2546
rect 3450 2543 3461 2546
rect 3426 2393 3429 2543
rect 3434 2453 3437 2526
rect 3450 2486 3453 2543
rect 3458 2533 3469 2536
rect 3466 2523 3469 2533
rect 3442 2483 3453 2486
rect 3434 2403 3437 2436
rect 3442 2386 3445 2483
rect 3450 2413 3453 2436
rect 3458 2413 3461 2496
rect 3474 2473 3477 2646
rect 3498 2626 3501 2693
rect 3514 2683 3517 2726
rect 3522 2723 3533 2726
rect 3498 2623 3509 2626
rect 3514 2623 3517 2636
rect 3522 2623 3525 2696
rect 3546 2663 3549 2726
rect 3554 2693 3557 2743
rect 3578 2736 3581 2783
rect 3562 2733 3581 2736
rect 3586 2733 3589 2776
rect 3598 2746 3601 2823
rect 3598 2743 3605 2746
rect 3482 2603 3493 2606
rect 3482 2543 3485 2603
rect 3498 2533 3501 2596
rect 3506 2553 3509 2623
rect 3514 2613 3525 2616
rect 3538 2613 3541 2636
rect 3514 2563 3517 2596
rect 3506 2523 3509 2536
rect 3482 2513 3493 2516
rect 3514 2513 3517 2536
rect 3530 2533 3533 2556
rect 3482 2466 3485 2513
rect 3522 2506 3525 2526
rect 3474 2463 3485 2466
rect 3450 2396 3453 2405
rect 3466 2403 3469 2456
rect 3474 2413 3477 2463
rect 3482 2403 3485 2436
rect 3490 2403 3493 2486
rect 3498 2396 3501 2506
rect 3450 2393 3501 2396
rect 3506 2503 3525 2506
rect 3506 2393 3509 2503
rect 3514 2396 3517 2476
rect 3522 2403 3525 2496
rect 3530 2413 3533 2456
rect 3538 2403 3541 2566
rect 3546 2473 3549 2626
rect 3554 2603 3557 2676
rect 3562 2596 3565 2733
rect 3570 2613 3573 2726
rect 3562 2593 3569 2596
rect 3554 2543 3557 2556
rect 3554 2483 3557 2536
rect 3566 2526 3569 2593
rect 3562 2523 3569 2526
rect 3546 2413 3549 2436
rect 3546 2403 3557 2406
rect 3514 2393 3533 2396
rect 3426 2383 3445 2386
rect 3482 2383 3493 2386
rect 3418 2373 3437 2376
rect 3410 2363 3421 2366
rect 3418 2276 3421 2363
rect 3434 2356 3437 2373
rect 3482 2366 3485 2383
rect 3482 2363 3489 2366
rect 3434 2353 3453 2356
rect 3434 2343 3445 2346
rect 3442 2323 3445 2343
rect 3418 2273 3437 2276
rect 3370 2263 3405 2266
rect 3358 2233 3365 2236
rect 3354 2193 3357 2216
rect 3338 2153 3349 2156
rect 3338 2113 3341 2153
rect 3346 2133 3349 2146
rect 3330 2093 3341 2096
rect 3290 1966 3293 2006
rect 3314 1993 3317 2036
rect 3322 2023 3325 2066
rect 3338 2026 3341 2093
rect 3354 2073 3357 2136
rect 3330 2023 3341 2026
rect 3290 1963 3325 1966
rect 3282 1953 3293 1956
rect 3290 1933 3293 1953
rect 3274 1903 3293 1906
rect 3258 1823 3269 1826
rect 3242 1793 3253 1796
rect 3242 1733 3245 1793
rect 3250 1766 3253 1786
rect 3258 1783 3261 1806
rect 3266 1776 3269 1806
rect 3274 1776 3277 1896
rect 3282 1803 3285 1856
rect 3266 1773 3277 1776
rect 3250 1763 3257 1766
rect 3186 1673 3197 1676
rect 3210 1703 3229 1706
rect 3186 1586 3189 1673
rect 3210 1616 3213 1703
rect 3234 1686 3237 1726
rect 3218 1683 3237 1686
rect 3218 1633 3221 1683
rect 3242 1676 3245 1726
rect 3254 1676 3257 1763
rect 3266 1753 3269 1766
rect 3274 1733 3277 1773
rect 3290 1756 3293 1903
rect 3314 1856 3317 1926
rect 3322 1903 3325 1963
rect 3306 1853 3317 1856
rect 3330 1846 3333 2023
rect 3314 1843 3333 1846
rect 3306 1783 3309 1826
rect 3314 1796 3317 1843
rect 3330 1803 3333 1826
rect 3314 1793 3333 1796
rect 3226 1673 3245 1676
rect 3250 1673 3257 1676
rect 3202 1613 3221 1616
rect 3194 1596 3197 1606
rect 3202 1603 3205 1613
rect 3194 1593 3205 1596
rect 3186 1583 3197 1586
rect 3194 1556 3197 1583
rect 3202 1576 3205 1593
rect 3210 1583 3213 1606
rect 3218 1576 3221 1606
rect 3202 1573 3221 1576
rect 3194 1553 3201 1556
rect 3186 1443 3189 1536
rect 3198 1436 3201 1553
rect 3218 1533 3221 1546
rect 3210 1503 3213 1516
rect 3218 1493 3221 1526
rect 3194 1433 3201 1436
rect 3170 1243 3173 1256
rect 3170 1166 3173 1236
rect 3178 1203 3181 1326
rect 3186 1196 3189 1376
rect 3194 1316 3197 1433
rect 3202 1333 3205 1416
rect 3210 1403 3213 1466
rect 3218 1413 3221 1446
rect 3226 1406 3229 1673
rect 3250 1636 3253 1673
rect 3274 1663 3277 1726
rect 3234 1633 3253 1636
rect 3234 1523 3237 1633
rect 3242 1576 3245 1606
rect 3258 1603 3261 1656
rect 3282 1586 3285 1756
rect 3290 1753 3301 1756
rect 3290 1613 3293 1736
rect 3298 1723 3301 1753
rect 3306 1733 3309 1766
rect 3314 1733 3317 1786
rect 3242 1573 3249 1576
rect 3246 1516 3249 1573
rect 3242 1513 3249 1516
rect 3242 1493 3245 1513
rect 3222 1403 3229 1406
rect 3234 1403 3237 1466
rect 3210 1343 3213 1386
rect 3222 1346 3225 1403
rect 3218 1343 3225 1346
rect 3210 1323 3213 1336
rect 3194 1313 3213 1316
rect 3194 1203 3197 1226
rect 3202 1213 3205 1306
rect 3162 1163 3173 1166
rect 3138 1123 3141 1136
rect 3146 1123 3149 1136
rect 3154 1123 3157 1156
rect 3162 1133 3165 1163
rect 3130 1113 3149 1116
rect 3146 1103 3149 1113
rect 3122 1083 3149 1086
rect 3106 1073 3133 1076
rect 3098 1063 3125 1066
rect 3090 1043 3097 1046
rect 3050 943 3069 946
rect 3018 873 3029 876
rect 3034 913 3045 916
rect 3010 803 3013 816
rect 2994 793 3005 796
rect 2978 753 2989 756
rect 2978 683 2981 746
rect 2986 676 2989 753
rect 2994 733 2997 786
rect 2978 673 2989 676
rect 2994 673 2997 726
rect 2954 583 2965 586
rect 2938 573 2949 576
rect 2978 573 2981 673
rect 2986 613 2989 656
rect 3002 616 3005 793
rect 3010 743 3013 786
rect 3018 776 3021 873
rect 3026 783 3029 826
rect 3034 803 3037 913
rect 3018 773 3037 776
rect 2994 613 3005 616
rect 3010 733 3029 736
rect 3034 733 3037 773
rect 2946 533 2949 573
rect 2986 566 2989 606
rect 2994 583 2997 613
rect 2954 563 2989 566
rect 2954 526 2957 563
rect 3010 556 3013 733
rect 3026 726 3029 733
rect 3042 726 3045 816
rect 3018 696 3021 726
rect 3026 723 3045 726
rect 3018 693 3029 696
rect 3018 603 3021 686
rect 3026 663 3029 693
rect 3034 643 3037 716
rect 2990 553 3013 556
rect 2962 533 2965 546
rect 2938 513 2941 526
rect 2946 523 2957 526
rect 2946 433 2949 523
rect 2922 373 2925 426
rect 2938 403 2941 426
rect 2946 396 2949 416
rect 2954 403 2957 516
rect 2962 396 2965 506
rect 2970 443 2973 536
rect 2914 363 2921 366
rect 2898 213 2901 363
rect 2918 316 2921 363
rect 2930 323 2933 396
rect 2946 393 2965 396
rect 2970 393 2973 406
rect 2978 386 2981 526
rect 2990 446 2993 553
rect 3026 546 3029 616
rect 3042 613 3045 716
rect 3034 583 3037 606
rect 2962 383 2981 386
rect 2986 443 2993 446
rect 2986 386 2989 443
rect 2986 383 2997 386
rect 2918 313 2925 316
rect 2938 313 2941 356
rect 2962 323 2965 383
rect 2970 333 2981 336
rect 2986 326 2989 336
rect 2994 333 2997 383
rect 3002 366 3005 536
rect 3010 533 3013 546
rect 3026 543 3037 546
rect 3018 503 3021 526
rect 3026 523 3029 536
rect 3034 463 3037 543
rect 3042 503 3045 536
rect 3026 413 3029 426
rect 3050 393 3053 943
rect 3074 936 3077 986
rect 3058 933 3077 936
rect 3058 843 3061 933
rect 3066 923 3077 926
rect 3082 906 3085 1006
rect 3094 986 3097 1043
rect 3090 983 3097 986
rect 3090 923 3093 983
rect 3098 923 3101 966
rect 3058 803 3061 816
rect 3066 803 3069 906
rect 3078 903 3085 906
rect 3098 903 3101 916
rect 3078 836 3081 903
rect 3106 896 3109 1006
rect 3114 1003 3117 1026
rect 3122 1013 3125 1063
rect 3114 933 3117 986
rect 3090 893 3109 896
rect 3078 833 3085 836
rect 3074 763 3077 816
rect 3066 743 3077 746
rect 3082 743 3085 833
rect 3090 763 3093 893
rect 3058 713 3061 736
rect 3066 683 3069 736
rect 3058 613 3061 626
rect 3066 603 3069 646
rect 3074 596 3077 743
rect 3082 733 3093 736
rect 3090 676 3093 726
rect 3082 673 3093 676
rect 3098 673 3101 846
rect 3106 813 3109 856
rect 3114 803 3117 926
rect 3122 923 3125 956
rect 3130 856 3133 1073
rect 3138 1013 3141 1066
rect 3138 923 3141 1006
rect 3146 996 3149 1083
rect 3154 1063 3157 1096
rect 3170 1056 3173 1146
rect 3178 1133 3181 1196
rect 3186 1193 3197 1196
rect 3186 1143 3189 1193
rect 3178 1123 3189 1126
rect 3154 1003 3157 1056
rect 3170 1053 3181 1056
rect 3178 1036 3181 1053
rect 3170 1033 3181 1036
rect 3162 1003 3165 1016
rect 3146 993 3165 996
rect 3146 983 3157 986
rect 3146 943 3149 956
rect 3138 863 3141 916
rect 3130 853 3141 856
rect 3122 816 3125 846
rect 3122 813 3133 816
rect 3138 806 3141 853
rect 3146 813 3149 936
rect 3106 693 3109 726
rect 3114 683 3117 766
rect 3122 666 3125 806
rect 3098 663 3125 666
rect 3130 803 3141 806
rect 3058 593 3077 596
rect 3058 513 3061 593
rect 3002 363 3013 366
rect 2970 323 2981 326
rect 2986 323 2997 326
rect 2874 123 2877 203
rect 2906 196 2909 206
rect 2914 203 2917 216
rect 2922 203 2925 313
rect 2962 196 2965 206
rect 2978 203 2981 286
rect 2994 203 2997 316
rect 3010 196 3013 363
rect 3034 303 3037 336
rect 3058 323 3061 336
rect 3074 303 3077 576
rect 3082 566 3085 656
rect 3098 576 3101 663
rect 3130 643 3133 803
rect 3138 783 3141 796
rect 3146 766 3149 806
rect 3154 803 3157 983
rect 3162 903 3165 993
rect 3170 933 3173 1033
rect 3170 863 3173 926
rect 3178 896 3181 1016
rect 3186 933 3189 1106
rect 3194 1053 3197 1166
rect 3202 1003 3205 1176
rect 3194 973 3197 986
rect 3202 963 3205 996
rect 3186 913 3189 926
rect 3178 893 3185 896
rect 3162 803 3165 816
rect 3170 813 3173 856
rect 3182 826 3185 893
rect 3194 883 3197 946
rect 3210 933 3213 1313
rect 3218 1006 3221 1343
rect 3226 1293 3229 1326
rect 3234 1273 3237 1336
rect 3242 1333 3245 1406
rect 3250 1333 3253 1386
rect 3234 1203 3237 1236
rect 3226 1123 3229 1186
rect 3234 1123 3237 1196
rect 3226 1086 3229 1106
rect 3234 1093 3237 1116
rect 3226 1083 3237 1086
rect 3226 1013 3229 1026
rect 3218 1003 3229 1006
rect 3202 876 3205 926
rect 3178 823 3185 826
rect 3194 873 3205 876
rect 3146 763 3173 766
rect 3146 686 3149 736
rect 3170 696 3173 763
rect 3138 683 3149 686
rect 3162 693 3173 696
rect 3122 583 3125 616
rect 3098 573 3117 576
rect 3082 563 3101 566
rect 3098 436 3101 563
rect 3106 523 3109 546
rect 3114 533 3117 573
rect 3094 433 3101 436
rect 3082 393 3085 416
rect 3094 386 3097 433
rect 3094 383 3101 386
rect 3098 366 3101 383
rect 3114 376 3117 406
rect 3138 376 3141 683
rect 3146 486 3149 676
rect 3162 656 3165 693
rect 3162 653 3169 656
rect 3166 596 3169 653
rect 3162 593 3169 596
rect 3162 576 3165 593
rect 3154 573 3165 576
rect 3154 503 3157 573
rect 3178 546 3181 823
rect 3186 783 3189 806
rect 3194 796 3197 873
rect 3218 866 3221 986
rect 3202 863 3221 866
rect 3202 803 3205 863
rect 3210 813 3213 846
rect 3226 813 3229 1003
rect 3194 793 3213 796
rect 3210 776 3213 793
rect 3210 773 3217 776
rect 3186 723 3189 736
rect 3194 716 3197 746
rect 3170 543 3181 546
rect 3186 713 3197 716
rect 3170 506 3173 543
rect 3178 516 3181 536
rect 3186 516 3189 713
rect 3214 706 3217 773
rect 3226 743 3229 806
rect 3210 703 3217 706
rect 3210 686 3213 703
rect 3206 683 3213 686
rect 3226 683 3229 726
rect 3194 613 3197 646
rect 3194 583 3197 606
rect 3206 556 3209 683
rect 3218 583 3221 606
rect 3202 553 3209 556
rect 3194 523 3197 536
rect 3178 513 3197 516
rect 3170 503 3181 506
rect 3146 483 3153 486
rect 3150 406 3153 483
rect 3178 456 3181 503
rect 3178 453 3185 456
rect 3162 413 3165 426
rect 3150 403 3165 406
rect 3114 373 3141 376
rect 3098 363 3105 366
rect 3102 316 3105 363
rect 3114 323 3117 356
rect 3098 313 3105 316
rect 3098 293 3101 313
rect 3026 223 3061 226
rect 3026 213 3029 223
rect 3034 203 3037 216
rect 2906 193 2933 196
rect 2962 193 2989 196
rect 2906 133 2909 156
rect 2930 123 2933 193
rect 2986 123 2989 193
rect 3002 193 3013 196
rect 3002 153 3005 193
rect 3010 133 3013 146
rect 3042 123 3045 206
rect 3050 203 3053 216
rect 3058 203 3061 223
rect 3066 203 3069 216
rect 3074 213 3077 226
rect 3090 123 3093 286
rect 3122 216 3125 326
rect 3138 303 3141 373
rect 3162 296 3165 403
rect 3182 376 3185 453
rect 3194 413 3197 513
rect 3106 213 3125 216
rect 3154 293 3165 296
rect 3178 373 3185 376
rect 3202 373 3205 553
rect 3106 203 3109 213
rect 3114 203 3149 206
rect 3122 133 3125 156
rect 3146 123 3149 203
rect 3154 163 3157 293
rect 3170 193 3173 216
rect 3178 203 3181 373
rect 3186 323 3189 336
rect 3210 326 3213 536
rect 3218 523 3221 566
rect 3226 546 3229 616
rect 3234 593 3237 1083
rect 3242 1003 3245 1136
rect 3250 1093 3253 1146
rect 3258 1073 3261 1586
rect 3278 1583 3285 1586
rect 3266 1483 3269 1536
rect 3278 1486 3281 1583
rect 3298 1576 3301 1696
rect 3314 1656 3317 1726
rect 3290 1573 3301 1576
rect 3306 1653 3317 1656
rect 3290 1513 3293 1573
rect 3298 1526 3301 1566
rect 3306 1543 3309 1653
rect 3322 1583 3325 1786
rect 3330 1563 3333 1793
rect 3338 1766 3341 2006
rect 3346 1786 3349 1876
rect 3354 1863 3357 2016
rect 3362 1873 3365 2233
rect 3370 2213 3373 2263
rect 3402 2243 3413 2246
rect 3378 2213 3397 2216
rect 3370 2123 3373 2206
rect 3378 2163 3381 2213
rect 3386 2203 3397 2206
rect 3402 2193 3405 2206
rect 3402 2136 3405 2156
rect 3378 2076 3381 2136
rect 3398 2133 3405 2136
rect 3386 2113 3389 2126
rect 3378 2073 3385 2076
rect 3370 1856 3373 2066
rect 3382 2026 3385 2073
rect 3398 2056 3401 2133
rect 3398 2053 3405 2056
rect 3382 2023 3389 2026
rect 3378 1883 3381 2016
rect 3386 1953 3389 2023
rect 3394 1933 3397 2036
rect 3402 2013 3405 2053
rect 3410 2003 3413 2243
rect 3418 1986 3421 2246
rect 3434 2153 3437 2273
rect 3450 2243 3453 2353
rect 3486 2286 3489 2363
rect 3498 2323 3501 2386
rect 3506 2343 3525 2346
rect 3530 2336 3533 2393
rect 3562 2383 3565 2523
rect 3570 2483 3573 2506
rect 3570 2413 3573 2456
rect 3570 2366 3573 2406
rect 3482 2283 3489 2286
rect 3458 2193 3461 2216
rect 3426 2113 3429 2136
rect 3434 2076 3437 2126
rect 3442 2093 3445 2136
rect 3450 2083 3453 2126
rect 3434 2073 3445 2076
rect 3442 2003 3445 2073
rect 3458 2056 3461 2136
rect 3466 2123 3469 2226
rect 3474 2133 3477 2236
rect 3482 2176 3485 2283
rect 3506 2246 3509 2266
rect 3502 2243 3509 2246
rect 3482 2173 3493 2176
rect 3454 2053 3461 2056
rect 3402 1983 3421 1986
rect 3362 1853 3373 1856
rect 3362 1803 3365 1853
rect 3346 1783 3365 1786
rect 3338 1763 3345 1766
rect 3342 1646 3345 1763
rect 3354 1723 3357 1766
rect 3342 1643 3349 1646
rect 3338 1613 3341 1636
rect 3346 1596 3349 1643
rect 3354 1603 3357 1706
rect 3346 1593 3357 1596
rect 3338 1583 3349 1586
rect 3314 1533 3333 1536
rect 3298 1523 3317 1526
rect 3298 1493 3301 1516
rect 3278 1483 3285 1486
rect 3282 1463 3285 1483
rect 3266 1423 3277 1426
rect 3266 1373 3269 1416
rect 3274 1333 3277 1406
rect 3266 1233 3269 1296
rect 3266 1173 3269 1226
rect 3274 1193 3277 1216
rect 3250 1003 3253 1016
rect 3258 983 3261 1056
rect 3266 976 3269 1126
rect 3274 1113 3277 1186
rect 3274 1023 3277 1106
rect 3274 1003 3277 1016
rect 3242 973 3269 976
rect 3274 973 3277 996
rect 3242 906 3245 973
rect 3258 933 3261 946
rect 3242 903 3253 906
rect 3242 883 3245 896
rect 3242 753 3245 796
rect 3242 583 3245 746
rect 3250 733 3253 903
rect 3258 806 3261 906
rect 3266 823 3269 866
rect 3274 833 3277 846
rect 3266 813 3277 816
rect 3258 803 3265 806
rect 3262 746 3265 803
rect 3262 743 3269 746
rect 3250 623 3253 706
rect 3258 616 3261 726
rect 3266 713 3269 743
rect 3274 733 3277 766
rect 3282 726 3285 1416
rect 3290 1323 3293 1386
rect 3298 1286 3301 1446
rect 3314 1436 3317 1523
rect 3322 1503 3325 1526
rect 3330 1513 3333 1533
rect 3338 1523 3341 1583
rect 3354 1576 3357 1593
rect 3346 1573 3357 1576
rect 3314 1433 3333 1436
rect 3322 1413 3325 1426
rect 3338 1413 3341 1506
rect 3346 1436 3349 1573
rect 3354 1533 3357 1546
rect 3354 1443 3357 1526
rect 3362 1446 3365 1783
rect 3386 1766 3389 1926
rect 3402 1876 3405 1983
rect 3454 1956 3457 2053
rect 3466 2003 3469 2046
rect 3474 2003 3477 2126
rect 3482 2053 3485 2156
rect 3454 1953 3461 1956
rect 3410 1933 3421 1936
rect 3394 1873 3405 1876
rect 3394 1803 3397 1873
rect 3402 1796 3405 1866
rect 3410 1813 3413 1856
rect 3426 1816 3429 1936
rect 3442 1913 3445 1926
rect 3458 1916 3461 1953
rect 3466 1943 3469 1956
rect 3474 1933 3477 1996
rect 3454 1913 3461 1916
rect 3466 1916 3469 1926
rect 3482 1923 3485 1966
rect 3490 1933 3493 2173
rect 3502 2166 3505 2243
rect 3502 2163 3509 2166
rect 3498 2053 3501 2146
rect 3506 2123 3509 2163
rect 3498 2023 3501 2046
rect 3506 2033 3509 2086
rect 3490 1916 3493 1926
rect 3466 1913 3493 1916
rect 3426 1813 3445 1816
rect 3402 1793 3409 1796
rect 3370 1763 3389 1766
rect 3370 1723 3373 1763
rect 3378 1713 3381 1746
rect 3386 1733 3389 1756
rect 3370 1613 3373 1706
rect 3386 1696 3389 1726
rect 3382 1693 3389 1696
rect 3382 1626 3385 1693
rect 3382 1623 3389 1626
rect 3386 1603 3389 1623
rect 3370 1453 3373 1596
rect 3386 1583 3389 1596
rect 3394 1566 3397 1786
rect 3406 1626 3409 1793
rect 3418 1723 3421 1766
rect 3434 1716 3437 1806
rect 3454 1776 3457 1913
rect 3466 1813 3469 1906
rect 3490 1876 3493 1913
rect 3498 1883 3501 2006
rect 3506 1983 3509 2026
rect 3514 1946 3517 2336
rect 3522 2333 3533 2336
rect 3538 2363 3573 2366
rect 3522 2123 3525 2333
rect 3530 2293 3533 2306
rect 3538 2243 3541 2363
rect 3578 2356 3581 2726
rect 3594 2693 3597 2726
rect 3586 2613 3589 2626
rect 3586 2513 3589 2526
rect 3586 2393 3589 2476
rect 3546 2353 3581 2356
rect 3546 2226 3549 2353
rect 3562 2333 3565 2346
rect 3586 2333 3589 2386
rect 3554 2323 3565 2326
rect 3554 2306 3557 2323
rect 3554 2303 3561 2306
rect 3558 2226 3561 2303
rect 3570 2233 3573 2326
rect 3578 2323 3589 2326
rect 3578 2306 3581 2323
rect 3594 2306 3597 2666
rect 3602 2593 3605 2743
rect 3610 2733 3613 2816
rect 3618 2783 3621 2806
rect 3610 2663 3613 2726
rect 3618 2723 3621 2776
rect 3626 2746 3629 2846
rect 3634 2803 3637 2826
rect 3642 2813 3645 2856
rect 3642 2803 3653 2806
rect 3682 2776 3685 2893
rect 3698 2883 3701 2936
rect 3706 2913 3709 2953
rect 3722 2933 3725 2966
rect 3722 2876 3725 2926
rect 3730 2923 3733 2936
rect 3738 2933 3741 2946
rect 3746 2923 3749 2976
rect 3754 2973 3773 2976
rect 3754 2933 3757 2973
rect 3718 2873 3725 2876
rect 3706 2813 3709 2826
rect 3658 2773 3685 2776
rect 3626 2743 3637 2746
rect 3626 2723 3629 2736
rect 3634 2726 3637 2743
rect 3642 2733 3653 2736
rect 3634 2723 3653 2726
rect 3634 2636 3637 2723
rect 3658 2706 3661 2773
rect 3650 2703 3661 2706
rect 3650 2643 3653 2703
rect 3658 2646 3661 2696
rect 3666 2663 3669 2766
rect 3658 2643 3669 2646
rect 3618 2633 3637 2636
rect 3610 2573 3613 2606
rect 3618 2536 3621 2633
rect 3634 2543 3637 2606
rect 3666 2566 3669 2643
rect 3682 2613 3685 2736
rect 3698 2733 3701 2776
rect 3718 2746 3721 2873
rect 3718 2743 3725 2746
rect 3690 2723 3709 2726
rect 3690 2703 3693 2723
rect 3602 2406 3605 2536
rect 3610 2533 3621 2536
rect 3610 2456 3613 2533
rect 3618 2523 3629 2526
rect 3634 2523 3637 2536
rect 3642 2533 3645 2556
rect 3650 2533 3653 2566
rect 3658 2563 3669 2566
rect 3618 2463 3621 2523
rect 3658 2513 3661 2563
rect 3666 2506 3669 2546
rect 3682 2513 3685 2536
rect 3698 2533 3701 2596
rect 3706 2566 3709 2646
rect 3714 2613 3717 2726
rect 3722 2693 3725 2743
rect 3722 2603 3725 2676
rect 3706 2563 3717 2566
rect 3706 2543 3709 2556
rect 3650 2503 3669 2506
rect 3610 2453 3621 2456
rect 3610 2413 3613 2436
rect 3602 2403 3613 2406
rect 3610 2383 3613 2403
rect 3602 2333 3605 2376
rect 3618 2356 3621 2453
rect 3626 2403 3629 2486
rect 3634 2356 3637 2416
rect 3618 2353 3637 2356
rect 3618 2323 3621 2353
rect 3626 2333 3629 2346
rect 3642 2333 3645 2456
rect 3650 2326 3653 2503
rect 3674 2413 3677 2506
rect 3690 2473 3693 2526
rect 3706 2516 3709 2536
rect 3702 2513 3709 2516
rect 3666 2393 3669 2406
rect 3682 2403 3685 2436
rect 3690 2386 3693 2446
rect 3702 2436 3705 2513
rect 3666 2383 3693 2386
rect 3698 2433 3705 2436
rect 3666 2333 3669 2383
rect 3698 2356 3701 2433
rect 3714 2403 3717 2563
rect 3730 2533 3733 2866
rect 3762 2863 3765 2936
rect 3770 2923 3773 2973
rect 3778 2913 3781 3016
rect 3786 3003 3789 3023
rect 3802 2996 3805 3063
rect 3794 2993 3805 2996
rect 3794 2843 3797 2993
rect 3818 2956 3821 3076
rect 3834 3013 3837 3036
rect 3818 2953 3829 2956
rect 3818 2923 3821 2946
rect 3762 2816 3765 2836
rect 3754 2813 3765 2816
rect 3754 2766 3757 2813
rect 3770 2793 3773 2816
rect 3778 2803 3781 2816
rect 3786 2793 3789 2816
rect 3802 2766 3805 2816
rect 3818 2813 3821 2866
rect 3810 2773 3813 2806
rect 3818 2793 3821 2806
rect 3754 2763 3765 2766
rect 3738 2733 3749 2736
rect 3738 2613 3741 2726
rect 3754 2643 3757 2746
rect 3762 2663 3765 2763
rect 3786 2763 3805 2766
rect 3770 2733 3773 2756
rect 3746 2616 3749 2626
rect 3746 2613 3757 2616
rect 3762 2573 3765 2606
rect 3770 2563 3773 2696
rect 3778 2606 3781 2726
rect 3786 2623 3789 2763
rect 3794 2656 3797 2726
rect 3802 2723 3805 2756
rect 3818 2743 3821 2766
rect 3810 2696 3813 2736
rect 3810 2693 3821 2696
rect 3826 2686 3829 2953
rect 3834 2893 3837 3006
rect 3842 2886 3845 3016
rect 3850 3003 3853 3126
rect 3898 3073 3901 3126
rect 3906 3123 3909 3233
rect 3914 3193 3917 3216
rect 3922 3203 3925 3216
rect 3946 3213 3949 3226
rect 3930 3196 3933 3206
rect 3938 3203 3949 3206
rect 3954 3196 3957 3216
rect 3962 3203 3965 3326
rect 4002 3323 4005 3333
rect 4010 3306 4013 3326
rect 4002 3303 4013 3306
rect 4002 3236 4005 3303
rect 3970 3233 4005 3236
rect 3970 3213 3973 3233
rect 4018 3226 4021 3333
rect 4034 3326 4037 3346
rect 4074 3336 4077 3346
rect 4042 3333 4053 3336
rect 4026 3323 4037 3326
rect 4026 3273 4029 3323
rect 4050 3313 4053 3326
rect 4058 3276 4061 3336
rect 4066 3333 4077 3336
rect 4090 3333 4093 3346
rect 4074 3276 4077 3326
rect 4082 3313 4085 3326
rect 4058 3273 4077 3276
rect 4098 3256 4101 3373
rect 4114 3343 4117 3546
rect 4130 3533 4133 3593
rect 4154 3586 4157 3683
rect 4162 3633 4165 3693
rect 4170 3663 4173 3753
rect 4178 3626 4181 3736
rect 4186 3683 4189 3963
rect 4194 3933 4197 3956
rect 4202 3943 4205 4006
rect 4194 3893 4197 3916
rect 4202 3833 4205 3936
rect 4210 3923 4213 4126
rect 4218 4123 4221 4136
rect 4250 4126 4253 4136
rect 4266 4133 4269 4206
rect 4282 4176 4285 4206
rect 4306 4203 4309 4216
rect 4354 4213 4365 4216
rect 4282 4173 4293 4176
rect 4250 4123 4269 4126
rect 4218 3906 4221 3946
rect 4226 3913 4229 4106
rect 4242 4103 4245 4116
rect 4290 4096 4293 4173
rect 4282 4093 4293 4096
rect 4250 4006 4253 4016
rect 4234 4003 4253 4006
rect 4266 4003 4269 4026
rect 4282 4003 4285 4093
rect 4314 4023 4317 4126
rect 4330 4106 4333 4126
rect 4326 4103 4333 4106
rect 4234 3983 4237 3996
rect 4306 3966 4309 4016
rect 4326 4006 4329 4103
rect 4338 4056 4341 4156
rect 4370 4136 4373 4256
rect 4362 4133 4373 4136
rect 4362 4086 4365 4133
rect 4378 4093 4381 4126
rect 4362 4083 4373 4086
rect 4338 4053 4349 4056
rect 4266 3963 4309 3966
rect 4322 4003 4329 4006
rect 4234 3943 4237 3956
rect 4234 3933 4253 3936
rect 4250 3923 4253 3933
rect 4258 3906 4261 3936
rect 4266 3933 4269 3963
rect 4214 3903 4221 3906
rect 4250 3903 4261 3906
rect 4214 3846 4217 3903
rect 4214 3843 4221 3846
rect 4194 3823 4213 3826
rect 4194 3763 4197 3823
rect 4202 3766 4205 3816
rect 4210 3813 4213 3823
rect 4210 3773 4213 3806
rect 4218 3786 4221 3843
rect 4226 3803 4229 3866
rect 4250 3836 4253 3903
rect 4282 3886 4285 3936
rect 4250 3833 4261 3836
rect 4234 3813 4253 3816
rect 4258 3806 4261 3833
rect 4218 3783 4229 3786
rect 4202 3763 4221 3766
rect 4194 3743 4205 3746
rect 4202 3636 4205 3736
rect 4210 3733 4213 3756
rect 4218 3743 4221 3763
rect 4226 3736 4229 3783
rect 4218 3733 4229 3736
rect 4218 3716 4221 3733
rect 4194 3633 4205 3636
rect 4214 3713 4221 3716
rect 4178 3623 4185 3626
rect 4146 3583 4157 3586
rect 4146 3543 4149 3583
rect 4162 3533 4165 3576
rect 4182 3546 4185 3623
rect 4194 3613 4197 3633
rect 4214 3626 4217 3713
rect 4226 3693 4229 3726
rect 4234 3676 4237 3766
rect 4242 3743 4245 3806
rect 4250 3803 4261 3806
rect 4266 3796 4269 3876
rect 4258 3793 4269 3796
rect 4242 3693 4245 3736
rect 4226 3673 4237 3676
rect 4226 3633 4229 3673
rect 4250 3663 4253 3726
rect 4202 3553 4205 3626
rect 4210 3623 4217 3626
rect 4182 3543 4197 3546
rect 4146 3506 4149 3526
rect 4186 3513 4189 3526
rect 4146 3503 4157 3506
rect 4122 3403 4125 3416
rect 4130 3403 4133 3416
rect 4138 3393 4141 3416
rect 4146 3403 4149 3456
rect 4154 3413 4157 3503
rect 4194 3446 4197 3543
rect 4210 3493 4213 3623
rect 4218 3596 4221 3616
rect 4226 3613 4229 3626
rect 4234 3606 4237 3656
rect 4258 3633 4261 3793
rect 4274 3763 4277 3886
rect 4282 3883 4293 3886
rect 4290 3756 4293 3883
rect 4306 3863 4309 3926
rect 4322 3836 4325 4003
rect 4346 3996 4349 4053
rect 4354 4013 4365 4016
rect 4346 3993 4353 3996
rect 4350 3906 4353 3993
rect 4362 3923 4365 3936
rect 4346 3903 4353 3906
rect 4370 3903 4373 4083
rect 4346 3886 4349 3903
rect 4338 3883 4349 3886
rect 4322 3833 4333 3836
rect 4274 3753 4293 3756
rect 4266 3723 4269 3736
rect 4226 3603 4237 3606
rect 4242 3603 4245 3626
rect 4250 3613 4269 3616
rect 4258 3596 4261 3606
rect 4218 3593 4261 3596
rect 4266 3593 4269 3606
rect 4274 3576 4277 3753
rect 4282 3716 4285 3726
rect 4290 3723 4293 3746
rect 4298 3736 4301 3776
rect 4298 3733 4309 3736
rect 4314 3733 4317 3816
rect 4330 3763 4333 3833
rect 4338 3776 4341 3883
rect 4354 3813 4373 3816
rect 4338 3773 4349 3776
rect 4330 3733 4333 3746
rect 4298 3716 4301 3726
rect 4282 3713 4301 3716
rect 4306 3663 4309 3733
rect 4322 3723 4341 3726
rect 4346 3716 4349 3773
rect 4354 3733 4357 3813
rect 4338 3713 4349 3716
rect 4314 3613 4317 3626
rect 4290 3576 4293 3606
rect 4322 3596 4325 3686
rect 4338 3666 4341 3713
rect 4274 3573 4293 3576
rect 4318 3593 4325 3596
rect 4330 3663 4341 3666
rect 4242 3523 4245 3566
rect 4282 3533 4285 3573
rect 4178 3443 4197 3446
rect 4162 3413 4173 3416
rect 4162 3403 4165 3413
rect 4170 3393 4173 3406
rect 4178 3346 4181 3443
rect 4186 3423 4213 3426
rect 4186 3363 4189 3423
rect 4202 3393 4205 3416
rect 4210 3413 4213 3423
rect 4234 3413 4253 3416
rect 4210 3376 4213 3406
rect 4226 3403 4237 3406
rect 4250 3393 4253 3406
rect 4258 3403 4261 3416
rect 4210 3373 4221 3376
rect 4178 3343 4185 3346
rect 4114 3256 4117 3336
rect 4138 3323 4141 3336
rect 4182 3286 4185 3343
rect 4194 3323 4197 3346
rect 4202 3316 4205 3336
rect 4210 3323 4213 3346
rect 4218 3336 4221 3373
rect 4218 3333 4229 3336
rect 4218 3316 4221 3326
rect 4202 3313 4221 3316
rect 4082 3253 4117 3256
rect 4178 3283 4185 3286
rect 3978 3203 3981 3226
rect 4018 3223 4029 3226
rect 3986 3203 3989 3216
rect 3930 3193 3957 3196
rect 4018 3196 4021 3216
rect 4026 3206 4029 3223
rect 4034 3213 4037 3226
rect 4050 3213 4069 3216
rect 4026 3203 4037 3206
rect 4042 3203 4053 3206
rect 4058 3196 4061 3206
rect 4074 3203 4077 3226
rect 4018 3193 4061 3196
rect 3930 3163 3933 3193
rect 3946 3126 3949 3136
rect 4018 3133 4021 3156
rect 3946 3123 4029 3126
rect 3858 2976 3861 3016
rect 3866 3003 3869 3036
rect 3882 3003 3893 3006
rect 3858 2973 3865 2976
rect 3862 2906 3865 2973
rect 3890 2933 3893 3003
rect 3898 2996 3901 3016
rect 3906 3013 3909 3026
rect 3906 3003 3917 3006
rect 3922 3003 3925 3026
rect 3930 2996 3933 3016
rect 3898 2993 3933 2996
rect 3954 3003 3965 3006
rect 3858 2903 3865 2906
rect 3834 2756 3837 2886
rect 3842 2883 3853 2886
rect 3858 2883 3861 2903
rect 3850 2816 3853 2883
rect 3874 2863 3877 2926
rect 3898 2893 3901 2926
rect 3906 2913 3909 2936
rect 3914 2903 3917 2993
rect 3954 2956 3957 3003
rect 3946 2953 3957 2956
rect 3922 2926 3925 2936
rect 3930 2933 3941 2936
rect 3922 2923 3933 2926
rect 3842 2763 3845 2816
rect 3850 2813 3861 2816
rect 3850 2783 3853 2806
rect 3858 2796 3861 2813
rect 3866 2803 3869 2826
rect 3874 2813 3877 2856
rect 3858 2793 3869 2796
rect 3834 2753 3861 2756
rect 3834 2733 3845 2736
rect 3818 2683 3829 2686
rect 3794 2653 3813 2656
rect 3794 2633 3797 2646
rect 3810 2643 3813 2653
rect 3794 2613 3797 2626
rect 3802 2613 3805 2636
rect 3778 2603 3805 2606
rect 3778 2556 3781 2596
rect 3762 2533 3765 2556
rect 3770 2553 3781 2556
rect 3730 2506 3733 2526
rect 3738 2513 3741 2526
rect 3746 2506 3749 2526
rect 3770 2506 3773 2553
rect 3730 2503 3749 2506
rect 3738 2393 3741 2416
rect 3690 2353 3701 2356
rect 3578 2303 3585 2306
rect 3594 2303 3605 2306
rect 3582 2236 3585 2303
rect 3578 2233 3585 2236
rect 3602 2236 3605 2303
rect 3634 2273 3637 2326
rect 3646 2323 3653 2326
rect 3646 2266 3649 2323
rect 3642 2263 3649 2266
rect 3602 2233 3613 2236
rect 3530 2213 3533 2226
rect 3542 2223 3549 2226
rect 3554 2223 3561 2226
rect 3530 2073 3533 2206
rect 3542 2166 3545 2223
rect 3542 2163 3549 2166
rect 3546 2146 3549 2163
rect 3554 2156 3557 2223
rect 3562 2173 3565 2206
rect 3570 2186 3573 2216
rect 3578 2213 3581 2233
rect 3594 2213 3597 2226
rect 3586 2193 3589 2206
rect 3602 2186 3605 2206
rect 3570 2183 3605 2186
rect 3554 2153 3581 2156
rect 3546 2143 3581 2146
rect 3522 1983 3525 2036
rect 3530 2023 3533 2056
rect 3538 2033 3541 2126
rect 3546 2093 3549 2136
rect 3554 2083 3557 2126
rect 3562 2103 3565 2136
rect 3570 2076 3573 2136
rect 3554 2073 3573 2076
rect 3506 1943 3517 1946
rect 3454 1773 3461 1776
rect 3434 1713 3441 1716
rect 3378 1523 3381 1566
rect 3390 1563 3397 1566
rect 3402 1623 3409 1626
rect 3390 1486 3393 1563
rect 3402 1546 3405 1623
rect 3410 1573 3413 1606
rect 3418 1566 3421 1656
rect 3426 1633 3429 1706
rect 3438 1646 3441 1713
rect 3434 1643 3441 1646
rect 3426 1573 3429 1616
rect 3418 1563 3429 1566
rect 3402 1543 3421 1546
rect 3402 1493 3405 1526
rect 3410 1496 3413 1536
rect 3418 1533 3421 1543
rect 3426 1523 3429 1563
rect 3410 1493 3421 1496
rect 3390 1483 3397 1486
rect 3362 1443 3373 1446
rect 3346 1433 3357 1436
rect 3306 1403 3325 1406
rect 3306 1333 3309 1346
rect 3298 1283 3309 1286
rect 3298 1253 3301 1276
rect 3306 1226 3309 1283
rect 3298 1223 3309 1226
rect 3298 1183 3301 1223
rect 3306 1213 3317 1216
rect 3306 1136 3309 1146
rect 3298 1133 3309 1136
rect 3290 1063 3293 1126
rect 3306 1093 3309 1126
rect 3290 903 3293 1016
rect 3298 1013 3301 1056
rect 3306 1033 3309 1076
rect 3314 1046 3317 1213
rect 3322 1103 3325 1316
rect 3330 1093 3333 1326
rect 3338 1303 3341 1336
rect 3346 1273 3349 1426
rect 3354 1253 3357 1433
rect 3362 1423 3365 1436
rect 3362 1383 3365 1406
rect 3362 1283 3365 1316
rect 3370 1246 3373 1443
rect 3394 1403 3397 1483
rect 3402 1413 3405 1436
rect 3410 1413 3413 1426
rect 3418 1403 3421 1456
rect 3378 1363 3393 1366
rect 3378 1353 3381 1363
rect 3378 1333 3381 1346
rect 3390 1316 3393 1363
rect 3402 1323 3405 1346
rect 3410 1323 3413 1336
rect 3418 1323 3421 1376
rect 3426 1333 3429 1516
rect 3390 1313 3397 1316
rect 3346 1243 3373 1246
rect 3338 1213 3341 1226
rect 3346 1156 3349 1243
rect 3338 1153 3349 1156
rect 3338 1123 3341 1153
rect 3338 1053 3341 1116
rect 3314 1043 3341 1046
rect 3306 1013 3317 1016
rect 3314 983 3317 1013
rect 3322 976 3325 1026
rect 3338 1016 3341 1043
rect 3346 1026 3349 1146
rect 3354 1133 3357 1236
rect 3362 1183 3365 1206
rect 3354 1103 3357 1126
rect 3362 1123 3365 1146
rect 3370 1116 3373 1236
rect 3386 1213 3389 1246
rect 3394 1236 3397 1313
rect 3394 1233 3405 1236
rect 3378 1193 3381 1206
rect 3394 1203 3397 1226
rect 3386 1193 3397 1196
rect 3362 1113 3373 1116
rect 3354 1033 3357 1096
rect 3362 1033 3365 1113
rect 3346 1023 3357 1026
rect 3298 973 3325 976
rect 3290 733 3293 836
rect 3298 753 3301 973
rect 3306 923 3309 946
rect 3322 886 3325 966
rect 3314 883 3325 886
rect 3306 803 3309 826
rect 3314 733 3317 883
rect 3330 863 3333 1016
rect 3338 1013 3349 1016
rect 3338 853 3341 986
rect 3354 963 3357 1023
rect 3322 836 3325 846
rect 3322 833 3341 836
rect 3282 723 3293 726
rect 3290 623 3293 723
rect 3250 613 3261 616
rect 3250 573 3253 613
rect 3226 543 3237 546
rect 3226 493 3229 536
rect 3234 533 3237 543
rect 3234 516 3237 526
rect 3242 523 3245 536
rect 3250 516 3253 526
rect 3234 513 3253 516
rect 3234 503 3237 513
rect 3266 506 3269 616
rect 3274 603 3293 606
rect 3298 593 3301 616
rect 3306 563 3309 716
rect 3322 703 3325 816
rect 3338 813 3341 833
rect 3330 803 3341 806
rect 3322 616 3325 626
rect 3314 613 3325 616
rect 3314 603 3317 613
rect 3322 583 3325 606
rect 3282 543 3309 546
rect 3282 533 3285 543
rect 3290 513 3293 526
rect 3298 506 3301 536
rect 3330 533 3333 736
rect 3346 673 3349 936
rect 3354 873 3357 926
rect 3362 853 3365 936
rect 3370 916 3373 1106
rect 3378 1083 3381 1146
rect 3386 1133 3389 1193
rect 3402 1146 3405 1233
rect 3410 1203 3413 1306
rect 3434 1286 3437 1643
rect 3450 1613 3453 1736
rect 3458 1733 3461 1773
rect 3466 1763 3469 1806
rect 3474 1756 3477 1876
rect 3490 1873 3501 1876
rect 3482 1803 3485 1856
rect 3466 1753 3477 1756
rect 3490 1756 3493 1816
rect 3498 1803 3501 1873
rect 3490 1753 3501 1756
rect 3506 1753 3509 1943
rect 3514 1783 3517 1936
rect 3466 1723 3469 1753
rect 3450 1546 3453 1606
rect 3442 1543 3453 1546
rect 3442 1523 3445 1543
rect 3442 1433 3445 1516
rect 3442 1413 3445 1426
rect 3450 1406 3453 1536
rect 3458 1433 3461 1536
rect 3466 1523 3469 1576
rect 3458 1413 3461 1426
rect 3442 1403 3453 1406
rect 3442 1333 3445 1403
rect 3450 1373 3453 1396
rect 3458 1356 3461 1406
rect 3466 1403 3469 1516
rect 3430 1283 3437 1286
rect 3430 1236 3433 1283
rect 3430 1233 3437 1236
rect 3418 1196 3421 1226
rect 3410 1193 3421 1196
rect 3426 1193 3429 1216
rect 3410 1176 3413 1186
rect 3410 1173 3421 1176
rect 3410 1153 3413 1166
rect 3402 1143 3413 1146
rect 3394 1133 3405 1136
rect 3378 1023 3381 1066
rect 3378 1003 3381 1016
rect 3378 933 3381 986
rect 3386 933 3389 1126
rect 3394 1083 3397 1133
rect 3402 1076 3405 1126
rect 3394 1073 3405 1076
rect 3394 1013 3397 1073
rect 3402 1013 3405 1066
rect 3394 943 3397 1006
rect 3410 983 3413 1143
rect 3418 1103 3421 1173
rect 3426 1073 3429 1176
rect 3418 1003 3421 1026
rect 3426 1003 3429 1016
rect 3434 976 3437 1233
rect 3442 1213 3445 1276
rect 3450 1223 3453 1356
rect 3458 1353 3469 1356
rect 3442 1183 3445 1206
rect 3442 1123 3445 1176
rect 3450 1106 3453 1216
rect 3458 1203 3461 1276
rect 3458 1123 3461 1186
rect 3450 1103 3457 1106
rect 3410 973 3437 976
rect 3442 973 3445 1086
rect 3454 1036 3457 1103
rect 3466 1083 3469 1346
rect 3474 1306 3477 1726
rect 3482 1533 3485 1586
rect 3490 1556 3493 1736
rect 3498 1706 3501 1753
rect 3522 1733 3525 1936
rect 3530 1933 3533 1956
rect 3530 1853 3533 1886
rect 3538 1836 3541 2006
rect 3530 1833 3541 1836
rect 3514 1713 3517 1726
rect 3530 1706 3533 1833
rect 3546 1803 3549 2016
rect 3554 1856 3557 2073
rect 3562 1903 3565 2026
rect 3570 2013 3573 2056
rect 3570 1866 3573 1936
rect 3578 1883 3581 2143
rect 3586 2073 3589 2176
rect 3610 2166 3613 2233
rect 3594 2163 3613 2166
rect 3618 2163 3621 2226
rect 3594 2106 3597 2163
rect 3602 2153 3613 2156
rect 3594 2103 3601 2106
rect 3586 2013 3589 2046
rect 3598 2036 3601 2103
rect 3610 2083 3613 2153
rect 3598 2033 3605 2036
rect 3602 2013 3605 2033
rect 3610 2006 3613 2076
rect 3594 1953 3597 2006
rect 3602 2003 3613 2006
rect 3586 1933 3597 1936
rect 3586 1923 3597 1926
rect 3602 1893 3605 2003
rect 3570 1863 3585 1866
rect 3554 1853 3573 1856
rect 3570 1786 3573 1853
rect 3562 1783 3573 1786
rect 3562 1756 3565 1783
rect 3582 1776 3585 1863
rect 3594 1803 3597 1816
rect 3538 1723 3541 1756
rect 3546 1753 3565 1756
rect 3570 1773 3585 1776
rect 3498 1703 3525 1706
rect 3530 1703 3537 1706
rect 3498 1603 3501 1616
rect 3490 1553 3509 1556
rect 3490 1523 3493 1546
rect 3482 1316 3485 1466
rect 3498 1446 3501 1536
rect 3514 1533 3517 1636
rect 3490 1443 3501 1446
rect 3490 1373 3493 1443
rect 3498 1403 3501 1436
rect 3490 1323 3493 1346
rect 3482 1313 3493 1316
rect 3474 1303 3485 1306
rect 3474 1214 3477 1246
rect 3474 1193 3477 1206
rect 3482 1203 3485 1303
rect 3490 1233 3493 1313
rect 3506 1293 3509 1526
rect 3514 1413 3517 1446
rect 3522 1413 3525 1703
rect 3534 1636 3537 1703
rect 3530 1633 3537 1636
rect 3546 1633 3549 1753
rect 3554 1733 3557 1746
rect 3562 1706 3565 1726
rect 3570 1723 3573 1773
rect 3610 1766 3613 1996
rect 3618 1943 3621 2016
rect 3626 1893 3629 2046
rect 3634 2003 3637 2146
rect 3642 2013 3645 2263
rect 3690 2256 3693 2353
rect 3698 2323 3701 2346
rect 3746 2336 3749 2503
rect 3738 2333 3749 2336
rect 3758 2503 3773 2506
rect 3738 2316 3741 2333
rect 3686 2253 3693 2256
rect 3734 2313 3741 2316
rect 3666 2193 3669 2216
rect 3674 2166 3677 2236
rect 3650 2163 3677 2166
rect 3650 2043 3653 2163
rect 3658 2086 3661 2126
rect 3686 2106 3689 2253
rect 3734 2246 3737 2313
rect 3734 2243 3741 2246
rect 3746 2243 3749 2326
rect 3722 2173 3725 2216
rect 3730 2213 3733 2226
rect 3730 2193 3733 2206
rect 3698 2123 3701 2146
rect 3714 2133 3717 2156
rect 3686 2103 3693 2106
rect 3658 2083 3685 2086
rect 3658 1996 3661 2016
rect 3666 2013 3669 2026
rect 3674 2003 3677 2046
rect 3682 2006 3685 2083
rect 3690 2013 3693 2103
rect 3698 2026 3701 2116
rect 3738 2036 3741 2243
rect 3758 2236 3761 2503
rect 3778 2393 3781 2536
rect 3786 2533 3789 2546
rect 3794 2533 3797 2556
rect 3802 2523 3805 2603
rect 3794 2383 3797 2416
rect 3802 2403 3805 2496
rect 3810 2466 3813 2626
rect 3818 2593 3821 2683
rect 3842 2626 3845 2726
rect 3826 2623 3845 2626
rect 3826 2596 3829 2623
rect 3842 2613 3853 2616
rect 3834 2603 3845 2606
rect 3826 2593 3837 2596
rect 3818 2523 3821 2546
rect 3826 2483 3829 2536
rect 3810 2463 3821 2466
rect 3818 2396 3821 2463
rect 3834 2453 3837 2593
rect 3850 2573 3853 2596
rect 3842 2513 3845 2536
rect 3850 2483 3853 2526
rect 3810 2393 3821 2396
rect 3770 2343 3781 2346
rect 3754 2233 3761 2236
rect 3754 2216 3757 2233
rect 3750 2213 3757 2216
rect 3770 2213 3773 2266
rect 3778 2233 3781 2336
rect 3786 2323 3789 2356
rect 3810 2346 3813 2393
rect 3794 2343 3813 2346
rect 3786 2213 3789 2316
rect 3750 2146 3753 2213
rect 3762 2193 3765 2206
rect 3794 2196 3797 2343
rect 3802 2313 3805 2336
rect 3818 2333 3821 2346
rect 3834 2326 3837 2446
rect 3858 2403 3861 2753
rect 3866 2723 3869 2793
rect 3882 2763 3885 2806
rect 3874 2656 3877 2736
rect 3890 2733 3893 2756
rect 3906 2746 3909 2846
rect 3930 2813 3933 2826
rect 3946 2746 3949 2953
rect 3962 2933 3965 2946
rect 3986 2913 3989 2926
rect 3994 2863 3997 3116
rect 4066 3106 4069 3136
rect 4082 3106 4085 3253
rect 4098 3153 4101 3246
rect 4122 3203 4125 3216
rect 4178 3213 4181 3283
rect 4186 3223 4213 3226
rect 4186 3183 4189 3223
rect 4194 3153 4197 3196
rect 4202 3183 4205 3216
rect 4210 3213 4213 3223
rect 4226 3216 4229 3333
rect 4234 3313 4237 3336
rect 4250 3333 4253 3346
rect 4266 3333 4269 3346
rect 4242 3323 4261 3326
rect 4274 3306 4277 3496
rect 4266 3303 4277 3306
rect 4218 3213 4229 3216
rect 4234 3213 4253 3216
rect 4218 3206 4221 3213
rect 4210 3203 4221 3206
rect 4226 3203 4237 3206
rect 4210 3193 4213 3203
rect 4250 3183 4253 3206
rect 4258 3193 4261 3206
rect 4066 3103 4085 3106
rect 4018 3013 4021 3026
rect 4066 3023 4085 3026
rect 4058 2976 4061 2986
rect 4050 2973 4061 2976
rect 4002 2876 4005 2936
rect 4042 2923 4045 2936
rect 4050 2933 4053 2973
rect 4066 2946 4069 3023
rect 4074 3003 4077 3016
rect 4082 3013 4085 3023
rect 4058 2943 4069 2946
rect 4050 2893 4053 2926
rect 4058 2906 4061 2943
rect 4066 2913 4069 2936
rect 4074 2923 4077 2996
rect 4082 2983 4085 3006
rect 4106 3003 4109 3126
rect 4114 2993 4117 3016
rect 4122 3013 4133 3016
rect 4138 3013 4149 3016
rect 4122 3003 4125 3013
rect 4130 2946 4133 3006
rect 4146 2966 4149 3006
rect 4138 2963 4149 2966
rect 4162 2946 4165 3126
rect 4170 3116 4173 3146
rect 4194 3143 4237 3146
rect 4194 3123 4197 3143
rect 4218 3133 4229 3136
rect 4234 3133 4237 3143
rect 4242 3133 4245 3146
rect 4266 3143 4269 3303
rect 4290 3256 4293 3486
rect 4306 3453 4309 3526
rect 4318 3476 4321 3593
rect 4330 3483 4333 3663
rect 4338 3566 4341 3626
rect 4338 3563 4349 3566
rect 4346 3486 4349 3563
rect 4354 3526 4357 3676
rect 4362 3533 4365 3766
rect 4370 3593 4373 3776
rect 4378 3576 4381 3856
rect 4370 3573 4381 3576
rect 4354 3523 4365 3526
rect 4370 3506 4373 3573
rect 4338 3483 4349 3486
rect 4362 3503 4373 3506
rect 4318 3473 4325 3476
rect 4314 3403 4317 3416
rect 4322 3413 4325 3473
rect 4338 3466 4341 3483
rect 4334 3463 4341 3466
rect 4334 3366 4337 3463
rect 4362 3446 4365 3503
rect 4362 3443 4373 3446
rect 4370 3423 4373 3443
rect 4354 3413 4373 3416
rect 4378 3406 4381 3536
rect 4362 3403 4381 3406
rect 4334 3363 4341 3366
rect 4338 3343 4341 3363
rect 4314 3313 4317 3326
rect 4282 3253 4293 3256
rect 4282 3133 4285 3253
rect 4306 3203 4309 3216
rect 4362 3193 4365 3403
rect 4370 3323 4373 3346
rect 4202 3116 4205 3126
rect 4226 3123 4245 3126
rect 4306 3123 4309 3136
rect 4362 3123 4365 3146
rect 4170 3113 4205 3116
rect 4178 3003 4181 3026
rect 4186 2973 4189 3016
rect 4194 3013 4205 3016
rect 4194 3003 4197 3013
rect 4202 2983 4205 3006
rect 4194 2963 4205 2966
rect 4082 2926 4085 2936
rect 4090 2933 4101 2936
rect 4114 2933 4117 2946
rect 4130 2943 4165 2946
rect 4082 2923 4093 2926
rect 4058 2903 4085 2906
rect 4002 2873 4013 2876
rect 3986 2793 3989 2816
rect 3994 2813 3997 2856
rect 3994 2786 3997 2806
rect 3986 2783 3997 2786
rect 4010 2776 4013 2873
rect 4026 2783 4029 2816
rect 4002 2773 4013 2776
rect 3906 2743 3917 2746
rect 3946 2743 3981 2746
rect 3882 2703 3885 2726
rect 3898 2673 3901 2736
rect 3874 2653 3901 2656
rect 3898 2613 3901 2653
rect 3874 2576 3877 2606
rect 3914 2596 3917 2743
rect 3930 2723 3933 2736
rect 3938 2733 3957 2736
rect 3906 2593 3917 2596
rect 3906 2576 3909 2593
rect 3874 2573 3909 2576
rect 3866 2473 3869 2546
rect 3866 2403 3869 2436
rect 3890 2426 3893 2573
rect 3922 2556 3925 2576
rect 3938 2563 3941 2733
rect 3946 2706 3949 2726
rect 3946 2703 3973 2706
rect 3946 2606 3949 2666
rect 3954 2613 3957 2696
rect 3962 2673 3973 2676
rect 3946 2603 3957 2606
rect 3922 2553 3929 2556
rect 3914 2513 3917 2526
rect 3874 2423 3885 2426
rect 3890 2423 3901 2426
rect 3842 2333 3845 2396
rect 3858 2333 3861 2396
rect 3882 2386 3885 2423
rect 3874 2383 3885 2386
rect 3874 2336 3877 2383
rect 3890 2346 3893 2416
rect 3898 2413 3901 2423
rect 3906 2413 3909 2476
rect 3914 2406 3917 2506
rect 3926 2486 3929 2553
rect 3898 2396 3901 2406
rect 3906 2403 3917 2406
rect 3922 2483 3929 2486
rect 3922 2396 3925 2483
rect 3930 2403 3933 2466
rect 3938 2396 3941 2456
rect 3946 2413 3949 2486
rect 3954 2443 3957 2603
rect 3898 2393 3925 2396
rect 3930 2393 3941 2396
rect 3906 2366 3909 2386
rect 3906 2363 3913 2366
rect 3898 2346 3901 2356
rect 3890 2343 3901 2346
rect 3874 2333 3885 2336
rect 3810 2323 3821 2326
rect 3818 2266 3821 2286
rect 3814 2263 3821 2266
rect 3786 2193 3797 2196
rect 3750 2143 3757 2146
rect 3746 2103 3749 2126
rect 3718 2033 3741 2036
rect 3698 2023 3709 2026
rect 3698 2013 3709 2016
rect 3682 2003 3692 2006
rect 3658 1993 3693 1996
rect 3642 1973 3677 1976
rect 3618 1863 3621 1886
rect 3578 1763 3613 1766
rect 3558 1703 3565 1706
rect 3530 1583 3533 1633
rect 3558 1626 3561 1703
rect 3570 1673 3573 1716
rect 3578 1696 3581 1763
rect 3618 1753 3621 1856
rect 3586 1703 3589 1726
rect 3602 1713 3605 1736
rect 3578 1693 3589 1696
rect 3586 1636 3589 1693
rect 3586 1633 3597 1636
rect 3554 1623 3561 1626
rect 3538 1563 3541 1616
rect 3546 1556 3549 1616
rect 3514 1393 3517 1406
rect 3490 1173 3493 1216
rect 3498 1166 3501 1276
rect 3506 1176 3509 1196
rect 3522 1193 3525 1216
rect 3506 1173 3525 1176
rect 3498 1163 3517 1166
rect 3450 1033 3457 1036
rect 3370 913 3377 916
rect 3374 846 3377 913
rect 3386 893 3389 926
rect 3354 763 3357 816
rect 3362 803 3365 846
rect 3370 843 3377 846
rect 3338 533 3341 616
rect 3346 603 3349 616
rect 3354 586 3357 616
rect 3350 583 3357 586
rect 3362 583 3365 606
rect 3350 526 3353 583
rect 3346 523 3353 526
rect 3362 523 3365 566
rect 3370 523 3373 843
rect 3378 813 3381 826
rect 3378 783 3381 806
rect 3386 803 3389 866
rect 3394 733 3397 936
rect 3402 803 3405 966
rect 3410 823 3413 973
rect 3450 963 3453 1033
rect 3466 1013 3469 1066
rect 3482 1026 3485 1136
rect 3474 1023 3485 1026
rect 3418 896 3421 946
rect 3434 923 3437 936
rect 3458 923 3461 1006
rect 3418 893 3429 896
rect 3426 846 3429 893
rect 3418 843 3429 846
rect 3418 823 3421 843
rect 3426 813 3437 816
rect 3410 736 3413 756
rect 3410 733 3417 736
rect 3378 603 3381 726
rect 3414 686 3417 733
rect 3426 723 3429 746
rect 3410 683 3417 686
rect 3386 613 3389 636
rect 3386 603 3397 606
rect 3386 563 3389 603
rect 3266 503 3301 506
rect 3226 403 3229 456
rect 3242 333 3245 356
rect 3210 323 3237 326
rect 3250 323 3253 416
rect 3274 376 3277 416
rect 3322 403 3325 436
rect 3338 396 3341 516
rect 3346 506 3349 523
rect 3378 516 3381 536
rect 3394 533 3397 596
rect 3354 513 3381 516
rect 3346 503 3357 506
rect 3346 403 3349 416
rect 3354 403 3357 503
rect 3386 443 3389 526
rect 3362 403 3365 426
rect 3338 393 3349 396
rect 3370 393 3373 416
rect 3394 403 3397 526
rect 3402 433 3405 646
rect 3410 493 3413 683
rect 3418 613 3429 616
rect 3434 613 3437 813
rect 3442 803 3445 816
rect 3450 756 3453 836
rect 3458 813 3461 826
rect 3466 793 3469 896
rect 3474 823 3477 1023
rect 3446 753 3453 756
rect 3446 706 3449 753
rect 3446 703 3453 706
rect 3450 626 3453 703
rect 3458 633 3461 656
rect 3418 486 3421 566
rect 3426 513 3429 606
rect 3442 603 3445 626
rect 3450 623 3461 626
rect 3450 556 3453 606
rect 3458 603 3461 623
rect 3442 553 3453 556
rect 3434 533 3437 546
rect 3442 526 3445 553
rect 3458 533 3461 596
rect 3466 563 3469 786
rect 3474 766 3477 816
rect 3482 803 3485 1006
rect 3498 1003 3501 1056
rect 3498 886 3501 966
rect 3490 883 3501 886
rect 3490 776 3493 883
rect 3498 873 3501 883
rect 3498 803 3501 816
rect 3490 773 3501 776
rect 3474 763 3493 766
rect 3490 693 3493 763
rect 3498 736 3501 773
rect 3506 753 3509 1146
rect 3514 1123 3517 1163
rect 3514 923 3517 1056
rect 3514 813 3517 856
rect 3522 783 3525 1173
rect 3530 933 3533 1556
rect 3538 1553 3549 1556
rect 3538 1463 3541 1553
rect 3546 1443 3549 1546
rect 3538 1403 3541 1426
rect 3538 1323 3541 1396
rect 3546 1383 3549 1406
rect 3554 1366 3557 1623
rect 3594 1616 3597 1633
rect 3602 1623 3605 1706
rect 3562 1603 3565 1616
rect 3570 1603 3581 1606
rect 3586 1603 3589 1616
rect 3594 1613 3613 1616
rect 3562 1563 3565 1586
rect 3578 1536 3581 1556
rect 3574 1533 3581 1536
rect 3562 1373 3565 1466
rect 3574 1436 3577 1533
rect 3586 1453 3589 1586
rect 3594 1573 3597 1606
rect 3594 1476 3597 1556
rect 3602 1483 3605 1606
rect 3610 1553 3613 1613
rect 3610 1506 3613 1526
rect 3618 1523 3621 1616
rect 3610 1503 3621 1506
rect 3618 1483 3621 1503
rect 3594 1473 3621 1476
rect 3574 1433 3581 1436
rect 3570 1403 3573 1416
rect 3578 1386 3581 1433
rect 3586 1403 3589 1446
rect 3594 1413 3605 1416
rect 3574 1383 3581 1386
rect 3550 1363 3557 1366
rect 3550 1286 3553 1363
rect 3574 1326 3577 1383
rect 3574 1323 3581 1326
rect 3586 1323 3589 1356
rect 3602 1323 3605 1406
rect 3618 1403 3621 1473
rect 3626 1366 3629 1886
rect 3634 1813 3637 1946
rect 3642 1916 3645 1973
rect 3658 1933 3661 1966
rect 3674 1963 3677 1973
rect 3666 1923 3669 1956
rect 3674 1923 3677 1936
rect 3682 1933 3685 1986
rect 3642 1913 3653 1916
rect 3650 1846 3653 1913
rect 3690 1883 3693 1993
rect 3666 1863 3685 1866
rect 3642 1843 3653 1846
rect 3634 1713 3637 1726
rect 3634 1623 3637 1646
rect 3634 1553 3637 1616
rect 3642 1583 3645 1843
rect 3634 1483 3637 1536
rect 3642 1493 3645 1526
rect 3634 1373 3637 1406
rect 3642 1403 3645 1426
rect 3610 1363 3629 1366
rect 3578 1306 3581 1323
rect 3578 1303 3589 1306
rect 3550 1283 3557 1286
rect 3538 1173 3541 1216
rect 3546 1213 3549 1266
rect 3546 1083 3549 1166
rect 3538 1003 3541 1076
rect 3538 926 3541 946
rect 3546 943 3549 1016
rect 3530 776 3533 926
rect 3538 923 3545 926
rect 3542 816 3545 923
rect 3538 813 3545 816
rect 3538 793 3541 813
rect 3554 803 3557 1283
rect 3562 1223 3565 1286
rect 3586 1246 3589 1303
rect 3578 1243 3589 1246
rect 3562 1193 3565 1206
rect 3570 1203 3573 1216
rect 3578 1186 3581 1243
rect 3610 1226 3613 1363
rect 3650 1346 3653 1826
rect 3658 1763 3661 1806
rect 3674 1796 3677 1816
rect 3682 1813 3685 1826
rect 3698 1823 3701 2006
rect 3706 1993 3709 2006
rect 3718 1966 3721 2033
rect 3730 2003 3733 2026
rect 3714 1963 3721 1966
rect 3706 1853 3709 1946
rect 3714 1906 3717 1963
rect 3722 1923 3725 1946
rect 3730 1933 3733 1986
rect 3738 1923 3741 2016
rect 3714 1903 3721 1906
rect 3690 1813 3701 1816
rect 3682 1803 3693 1806
rect 3706 1796 3709 1806
rect 3674 1793 3709 1796
rect 3718 1786 3721 1903
rect 3730 1893 3741 1896
rect 3746 1893 3749 2096
rect 3754 1956 3757 2143
rect 3762 1973 3765 2146
rect 3786 2136 3789 2193
rect 3802 2143 3805 2216
rect 3814 2186 3817 2263
rect 3826 2243 3829 2326
rect 3834 2323 3845 2326
rect 3834 2306 3837 2323
rect 3834 2303 3841 2306
rect 3882 2303 3885 2333
rect 3890 2313 3893 2336
rect 3898 2323 3901 2343
rect 3814 2183 3821 2186
rect 3818 2163 3821 2183
rect 3786 2133 3813 2136
rect 3794 2113 3797 2126
rect 3770 2003 3773 2046
rect 3778 2003 3781 2016
rect 3786 2003 3789 2106
rect 3802 2093 3805 2126
rect 3794 2013 3797 2026
rect 3802 1993 3805 2006
rect 3754 1953 3765 1956
rect 3754 1933 3757 1946
rect 3762 1926 3765 1953
rect 3754 1923 3765 1926
rect 3770 1923 3773 1936
rect 3778 1933 3781 1976
rect 3786 1926 3789 1966
rect 3778 1923 3789 1926
rect 3714 1783 3721 1786
rect 3666 1686 3669 1716
rect 3658 1683 3669 1686
rect 3658 1603 3661 1683
rect 3666 1603 3669 1656
rect 3658 1403 3661 1526
rect 3666 1463 3669 1586
rect 3674 1523 3677 1766
rect 3682 1703 3685 1726
rect 3682 1613 3685 1636
rect 3682 1573 3685 1606
rect 3690 1603 3693 1736
rect 3690 1556 3693 1596
rect 3698 1573 3701 1726
rect 3706 1603 3709 1716
rect 3690 1553 3701 1556
rect 3650 1343 3657 1346
rect 3626 1243 3629 1336
rect 3654 1256 3657 1343
rect 3666 1293 3669 1416
rect 3690 1413 3693 1536
rect 3682 1366 3685 1406
rect 3698 1396 3701 1553
rect 3706 1503 3709 1536
rect 3714 1496 3717 1783
rect 3730 1733 3733 1886
rect 3722 1613 3725 1726
rect 3730 1626 3733 1686
rect 3738 1643 3741 1893
rect 3746 1783 3749 1886
rect 3746 1733 3749 1746
rect 3746 1633 3749 1706
rect 3730 1623 3749 1626
rect 3730 1613 3741 1616
rect 3722 1593 3725 1606
rect 3674 1363 3685 1366
rect 3694 1393 3701 1396
rect 3706 1493 3717 1496
rect 3674 1323 3677 1363
rect 3694 1306 3697 1393
rect 3574 1183 3581 1186
rect 3586 1223 3613 1226
rect 3562 1013 3565 1126
rect 3574 1116 3577 1183
rect 3586 1163 3589 1223
rect 3594 1193 3597 1216
rect 3602 1183 3605 1206
rect 3594 1163 3605 1166
rect 3594 1133 3597 1163
rect 3610 1143 3613 1216
rect 3626 1213 3629 1226
rect 3618 1123 3621 1206
rect 3634 1193 3637 1206
rect 3642 1176 3645 1256
rect 3638 1173 3645 1176
rect 3650 1253 3657 1256
rect 3574 1113 3581 1116
rect 3570 1003 3573 1096
rect 3530 773 3537 776
rect 3546 773 3549 796
rect 3498 733 3505 736
rect 3474 553 3477 656
rect 3482 583 3485 606
rect 3434 523 3445 526
rect 3410 483 3421 486
rect 3410 403 3413 483
rect 3274 373 3333 376
rect 3266 333 3277 336
rect 3282 306 3285 326
rect 3290 323 3293 336
rect 3274 303 3285 306
rect 3274 246 3277 303
rect 3274 243 3285 246
rect 3226 213 3229 226
rect 3282 223 3285 243
rect 3290 213 3293 276
rect 3218 196 3221 206
rect 3218 193 3261 196
rect 3202 123 3205 166
rect 3234 133 3237 146
rect 3258 123 3261 193
rect 3266 166 3269 206
rect 3298 183 3301 356
rect 3330 333 3333 373
rect 3346 333 3349 393
rect 3354 333 3357 356
rect 3306 253 3309 326
rect 3306 213 3309 236
rect 3322 216 3325 226
rect 3338 216 3341 326
rect 3362 323 3365 346
rect 3386 333 3397 336
rect 3418 333 3421 346
rect 3434 333 3437 523
rect 3450 453 3453 526
rect 3466 513 3469 526
rect 3474 503 3477 536
rect 3490 506 3493 686
rect 3502 676 3505 733
rect 3514 686 3517 726
rect 3534 696 3537 773
rect 3546 723 3549 736
rect 3562 706 3565 936
rect 3570 923 3573 946
rect 3570 813 3573 826
rect 3578 736 3581 1113
rect 3638 1106 3641 1173
rect 3650 1163 3653 1253
rect 3658 1213 3661 1236
rect 3666 1193 3669 1206
rect 3674 1186 3677 1306
rect 3694 1303 3701 1306
rect 3690 1223 3693 1286
rect 3698 1273 3701 1303
rect 3666 1183 3677 1186
rect 3586 973 3589 1106
rect 3638 1103 3645 1106
rect 3594 993 3597 1086
rect 3602 996 3605 1016
rect 3610 1003 3613 1076
rect 3602 993 3613 996
rect 3586 923 3589 936
rect 3594 933 3597 946
rect 3602 923 3605 976
rect 3610 933 3613 993
rect 3618 916 3621 1016
rect 3626 1003 3629 1096
rect 3642 1086 3645 1103
rect 3642 1083 3653 1086
rect 3658 1083 3661 1146
rect 3634 1003 3637 1076
rect 3590 913 3621 916
rect 3590 856 3593 913
rect 3626 906 3629 996
rect 3642 946 3645 1056
rect 3634 943 3645 946
rect 3634 923 3637 943
rect 3642 906 3645 936
rect 3650 923 3653 1083
rect 3666 1053 3669 1183
rect 3674 1036 3677 1176
rect 3682 1053 3685 1206
rect 3690 1106 3693 1196
rect 3698 1166 3701 1256
rect 3706 1173 3709 1493
rect 3714 1403 3717 1426
rect 3714 1323 3717 1376
rect 3714 1203 3717 1236
rect 3722 1203 3725 1576
rect 3698 1163 3709 1166
rect 3714 1163 3717 1196
rect 3706 1133 3709 1163
rect 3722 1143 3725 1176
rect 3690 1103 3701 1106
rect 3658 1033 3677 1036
rect 3658 1013 3661 1033
rect 3666 986 3669 1016
rect 3666 983 3677 986
rect 3658 923 3661 936
rect 3666 923 3669 976
rect 3674 933 3677 983
rect 3626 903 3633 906
rect 3642 903 3653 906
rect 3682 903 3685 1016
rect 3690 1003 3693 1096
rect 3698 1013 3701 1103
rect 3586 853 3593 856
rect 3586 823 3589 853
rect 3586 803 3589 816
rect 3578 733 3585 736
rect 3530 693 3537 696
rect 3554 703 3565 706
rect 3514 683 3525 686
rect 3502 673 3517 676
rect 3498 566 3501 616
rect 3498 563 3509 566
rect 3514 556 3517 673
rect 3522 603 3525 683
rect 3530 673 3533 693
rect 3506 553 3517 556
rect 3506 536 3509 553
rect 3482 503 3493 506
rect 3502 533 3509 536
rect 3482 486 3485 503
rect 3478 483 3485 486
rect 3458 413 3461 426
rect 3478 366 3481 483
rect 3490 413 3493 496
rect 3502 436 3505 533
rect 3514 446 3517 526
rect 3522 463 3525 576
rect 3530 523 3533 636
rect 3530 493 3533 516
rect 3514 443 3525 446
rect 3502 433 3509 436
rect 3474 363 3481 366
rect 3498 366 3501 416
rect 3506 413 3509 433
rect 3498 363 3505 366
rect 3394 313 3397 326
rect 3458 323 3461 336
rect 3378 216 3381 226
rect 3322 213 3341 216
rect 3354 213 3381 216
rect 3314 203 3325 206
rect 3354 203 3357 213
rect 3362 183 3365 206
rect 3266 163 3317 166
rect 3314 123 3317 163
rect 3346 133 3349 156
rect 3370 123 3373 206
rect 3378 166 3381 206
rect 3394 183 3397 206
rect 3402 173 3405 216
rect 3450 213 3453 296
rect 3474 286 3477 363
rect 3474 283 3485 286
rect 3482 263 3485 283
rect 3502 276 3505 363
rect 3514 286 3517 436
rect 3522 383 3525 443
rect 3530 403 3533 426
rect 3530 323 3533 346
rect 3538 326 3541 536
rect 3546 533 3549 596
rect 3554 566 3557 703
rect 3570 613 3573 726
rect 3582 676 3585 733
rect 3594 706 3597 836
rect 3602 823 3605 886
rect 3610 733 3613 816
rect 3618 803 3621 866
rect 3630 816 3633 903
rect 3650 826 3653 903
rect 3690 896 3693 996
rect 3698 933 3701 946
rect 3706 916 3709 1126
rect 3730 1086 3733 1606
rect 3738 1566 3741 1596
rect 3746 1573 3749 1606
rect 3738 1563 3749 1566
rect 3738 1513 3741 1536
rect 3746 1533 3749 1563
rect 3738 1296 3741 1506
rect 3746 1416 3749 1516
rect 3754 1503 3757 1923
rect 3778 1916 3781 1923
rect 3762 1913 3781 1916
rect 3762 1723 3765 1913
rect 3786 1863 3789 1916
rect 3794 1856 3797 1936
rect 3770 1803 3773 1856
rect 3778 1853 3797 1856
rect 3778 1813 3781 1853
rect 3802 1813 3805 1976
rect 3778 1796 3781 1806
rect 3786 1796 3789 1806
rect 3778 1793 3789 1796
rect 3746 1413 3757 1416
rect 3746 1383 3749 1406
rect 3762 1366 3765 1686
rect 3770 1676 3773 1746
rect 3778 1683 3781 1793
rect 3786 1723 3789 1786
rect 3802 1763 3805 1806
rect 3810 1783 3813 2133
rect 3818 2103 3821 2126
rect 3818 1933 3821 2016
rect 3826 1963 3829 2236
rect 3838 2226 3841 2303
rect 3890 2273 3893 2306
rect 3910 2276 3913 2363
rect 3922 2333 3925 2376
rect 3910 2273 3917 2276
rect 3834 2223 3841 2226
rect 3834 2173 3837 2223
rect 3850 2213 3853 2266
rect 3866 2213 3869 2226
rect 3842 2203 3853 2206
rect 3858 2203 3869 2206
rect 3850 2156 3853 2203
rect 3850 2153 3861 2156
rect 3834 2143 3853 2146
rect 3834 2123 3837 2143
rect 3842 2123 3845 2136
rect 3850 2133 3853 2143
rect 3834 2043 3845 2046
rect 3850 2043 3853 2126
rect 3826 1923 3829 1946
rect 3834 1923 3837 1936
rect 3842 1916 3845 2043
rect 3834 1913 3845 1916
rect 3818 1756 3821 1896
rect 3834 1893 3837 1913
rect 3850 1906 3853 2026
rect 3858 2013 3861 2153
rect 3866 2113 3869 2166
rect 3866 2013 3869 2026
rect 3858 2003 3869 2006
rect 3842 1903 3853 1906
rect 3842 1886 3845 1903
rect 3802 1753 3821 1756
rect 3826 1883 3845 1886
rect 3826 1756 3829 1883
rect 3834 1813 3845 1816
rect 3834 1763 3837 1806
rect 3850 1796 3853 1896
rect 3842 1793 3853 1796
rect 3826 1753 3837 1756
rect 3802 1733 3805 1753
rect 3810 1733 3821 1736
rect 3794 1683 3797 1726
rect 3802 1723 3813 1726
rect 3802 1703 3805 1723
rect 3826 1713 3829 1726
rect 3834 1706 3837 1753
rect 3826 1703 3837 1706
rect 3770 1673 3781 1676
rect 3770 1603 3773 1636
rect 3778 1623 3781 1673
rect 3786 1653 3813 1656
rect 3786 1643 3789 1653
rect 3794 1616 3797 1626
rect 3786 1613 3797 1616
rect 3770 1523 3773 1596
rect 3786 1546 3789 1613
rect 3802 1606 3805 1646
rect 3810 1613 3813 1653
rect 3794 1603 3805 1606
rect 3794 1553 3797 1603
rect 3778 1543 3789 1546
rect 3770 1373 3773 1416
rect 3762 1363 3773 1366
rect 3770 1353 3773 1363
rect 3738 1293 3745 1296
rect 3742 1246 3745 1293
rect 3754 1286 3757 1336
rect 3754 1283 3765 1286
rect 3762 1253 3765 1283
rect 3742 1243 3753 1246
rect 3738 1213 3741 1236
rect 3738 1193 3741 1206
rect 3750 1156 3753 1243
rect 3762 1193 3765 1216
rect 3770 1183 3773 1206
rect 3750 1153 3757 1156
rect 3726 1083 3733 1086
rect 3714 993 3717 1006
rect 3726 996 3729 1083
rect 3738 1003 3741 1146
rect 3746 1123 3749 1136
rect 3754 1106 3757 1153
rect 3750 1103 3757 1106
rect 3750 1036 3753 1103
rect 3750 1033 3757 1036
rect 3746 1003 3749 1016
rect 3726 993 3733 996
rect 3730 933 3733 993
rect 3746 983 3749 996
rect 3754 993 3757 1033
rect 3762 986 3765 1056
rect 3754 983 3765 986
rect 3714 923 3725 926
rect 3706 913 3725 916
rect 3674 893 3693 896
rect 3674 836 3677 893
rect 3674 833 3681 836
rect 3650 823 3669 826
rect 3626 813 3633 816
rect 3618 723 3621 736
rect 3626 706 3629 813
rect 3642 803 3645 816
rect 3666 806 3669 823
rect 3634 733 3637 796
rect 3650 753 3653 806
rect 3658 803 3669 806
rect 3594 703 3605 706
rect 3578 673 3585 676
rect 3578 653 3581 673
rect 3602 636 3605 703
rect 3594 633 3605 636
rect 3618 703 3629 706
rect 3618 636 3621 703
rect 3618 633 3629 636
rect 3586 613 3589 626
rect 3594 616 3597 633
rect 3626 616 3629 633
rect 3594 613 3605 616
rect 3618 613 3629 616
rect 3634 613 3637 716
rect 3650 613 3653 686
rect 3562 573 3565 606
rect 3570 603 3581 606
rect 3554 563 3565 566
rect 3570 563 3573 603
rect 3594 593 3597 606
rect 3546 496 3549 526
rect 3546 493 3557 496
rect 3546 403 3549 456
rect 3554 413 3557 493
rect 3562 476 3565 563
rect 3570 523 3573 536
rect 3570 493 3573 516
rect 3562 473 3569 476
rect 3566 406 3569 473
rect 3554 333 3557 406
rect 3562 403 3569 406
rect 3578 403 3581 546
rect 3562 383 3565 403
rect 3578 333 3581 346
rect 3538 323 3553 326
rect 3514 283 3525 286
rect 3502 273 3509 276
rect 3442 196 3445 206
rect 3442 193 3485 196
rect 3378 163 3429 166
rect 3426 123 3429 163
rect 3458 123 3461 136
rect 3482 123 3485 193
rect 3490 166 3493 206
rect 3506 203 3509 273
rect 3522 236 3525 283
rect 3514 233 3525 236
rect 3514 213 3517 233
rect 3538 213 3541 316
rect 3550 236 3553 323
rect 3550 233 3557 236
rect 3554 213 3557 233
rect 3546 166 3549 206
rect 3562 203 3565 326
rect 3586 273 3589 536
rect 3602 506 3605 613
rect 3658 606 3661 803
rect 3610 533 3613 606
rect 3650 603 3661 606
rect 3666 603 3669 796
rect 3678 756 3681 833
rect 3690 803 3693 826
rect 3674 753 3681 756
rect 3698 753 3701 886
rect 3722 856 3725 913
rect 3722 853 3733 856
rect 3714 813 3717 836
rect 3706 783 3709 806
rect 3674 643 3677 753
rect 3618 533 3621 546
rect 3610 513 3613 526
rect 3626 506 3629 556
rect 3650 536 3653 603
rect 3658 543 3661 596
rect 3594 333 3597 506
rect 3602 503 3613 506
rect 3602 423 3605 496
rect 3610 403 3613 503
rect 3622 503 3629 506
rect 3634 503 3637 536
rect 3650 533 3661 536
rect 3642 513 3645 526
rect 3622 436 3625 503
rect 3658 496 3661 526
rect 3650 493 3661 496
rect 3622 433 3629 436
rect 3602 333 3605 386
rect 3610 343 3613 396
rect 3610 283 3613 326
rect 3618 253 3621 416
rect 3626 333 3629 433
rect 3634 403 3637 466
rect 3650 406 3653 493
rect 3666 453 3669 596
rect 3674 506 3677 616
rect 3682 553 3685 736
rect 3690 713 3693 726
rect 3706 683 3709 776
rect 3690 653 3709 656
rect 3690 613 3693 653
rect 3698 613 3701 646
rect 3706 623 3709 653
rect 3722 636 3725 806
rect 3730 796 3733 853
rect 3738 803 3741 836
rect 3746 823 3749 906
rect 3730 793 3741 796
rect 3730 706 3733 726
rect 3738 723 3741 793
rect 3746 733 3749 786
rect 3730 703 3741 706
rect 3738 636 3741 703
rect 3714 633 3725 636
rect 3730 633 3741 636
rect 3754 636 3757 983
rect 3770 973 3773 1166
rect 3778 1123 3781 1543
rect 3810 1533 3813 1606
rect 3818 1603 3821 1626
rect 3826 1613 3829 1703
rect 3842 1643 3845 1793
rect 3858 1733 3861 1996
rect 3874 1963 3877 2246
rect 3890 2203 3893 2236
rect 3914 2216 3917 2273
rect 3930 2243 3933 2393
rect 3938 2333 3941 2346
rect 3954 2333 3957 2356
rect 3946 2283 3949 2326
rect 3962 2276 3965 2673
rect 3978 2626 3981 2743
rect 4002 2736 4005 2773
rect 4034 2743 4037 2816
rect 4042 2736 4045 2816
rect 4002 2733 4025 2736
rect 3986 2703 3989 2716
rect 3970 2623 3981 2626
rect 3970 2586 3973 2623
rect 3978 2593 3981 2616
rect 3986 2603 3989 2686
rect 4002 2683 4005 2706
rect 4010 2673 4013 2716
rect 4022 2676 4025 2733
rect 4034 2733 4045 2736
rect 4050 2736 4053 2806
rect 4058 2793 4061 2806
rect 4066 2786 4069 2836
rect 4074 2813 4077 2886
rect 4082 2813 4085 2903
rect 4098 2893 4101 2933
rect 4146 2926 4149 2943
rect 4138 2913 4141 2926
rect 4146 2923 4153 2926
rect 4098 2813 4101 2856
rect 4090 2793 4093 2806
rect 4066 2783 4093 2786
rect 4050 2733 4069 2736
rect 4022 2673 4029 2676
rect 4002 2653 4021 2656
rect 4002 2616 4005 2653
rect 4018 2633 4021 2653
rect 4026 2626 4029 2673
rect 3994 2613 4005 2616
rect 4010 2623 4029 2626
rect 4034 2623 4037 2733
rect 4042 2696 4045 2726
rect 4058 2703 4061 2726
rect 4074 2723 4077 2766
rect 4082 2696 4085 2776
rect 4042 2693 4085 2696
rect 4090 2686 4093 2783
rect 4106 2766 4109 2806
rect 4114 2783 4117 2806
rect 4122 2786 4125 2826
rect 4130 2796 4133 2816
rect 4138 2813 4141 2906
rect 4150 2856 4153 2923
rect 4146 2853 4153 2856
rect 4146 2833 4149 2853
rect 4162 2813 4165 2856
rect 4138 2803 4149 2806
rect 4154 2803 4165 2806
rect 4170 2796 4173 2806
rect 4130 2793 4173 2796
rect 4122 2783 4141 2786
rect 4098 2763 4133 2766
rect 4098 2723 4101 2763
rect 4114 2733 4117 2756
rect 4130 2733 4133 2763
rect 4138 2733 4141 2783
rect 4074 2683 4093 2686
rect 4050 2633 4069 2636
rect 3970 2583 3981 2586
rect 3970 2523 3973 2556
rect 3978 2533 3981 2583
rect 3986 2546 3989 2576
rect 4002 2563 4005 2606
rect 4010 2573 4013 2623
rect 3986 2543 3997 2546
rect 3978 2426 3981 2526
rect 3994 2446 3997 2543
rect 4018 2536 4021 2566
rect 4010 2533 4021 2536
rect 4018 2456 4021 2526
rect 4026 2506 4029 2576
rect 4034 2526 4037 2586
rect 4042 2533 4045 2546
rect 4034 2523 4045 2526
rect 4026 2503 4033 2506
rect 3970 2423 3981 2426
rect 3986 2443 3997 2446
rect 4010 2453 4021 2456
rect 3970 2383 3973 2423
rect 3938 2273 3965 2276
rect 3978 2273 3981 2416
rect 3986 2403 3989 2443
rect 4002 2403 4005 2426
rect 4010 2416 4013 2453
rect 4030 2426 4033 2503
rect 4030 2423 4037 2426
rect 4010 2413 4029 2416
rect 4002 2323 4005 2346
rect 4010 2316 4013 2406
rect 4002 2313 4013 2316
rect 3914 2213 3925 2216
rect 3938 2213 3941 2273
rect 4002 2256 4005 2313
rect 3998 2253 4005 2256
rect 3898 2203 3909 2206
rect 3898 2193 3901 2203
rect 3906 2156 3909 2196
rect 3922 2166 3925 2213
rect 3954 2203 3957 2216
rect 3978 2203 3981 2216
rect 3882 2153 3909 2156
rect 3914 2163 3925 2166
rect 3882 2136 3885 2153
rect 3914 2146 3917 2163
rect 3898 2143 3917 2146
rect 3882 2133 3901 2136
rect 3906 2133 3917 2136
rect 3898 2113 3901 2133
rect 3882 2086 3885 2106
rect 3882 2083 3889 2086
rect 3886 2006 3889 2083
rect 3882 2003 3889 2006
rect 3898 2003 3901 2016
rect 3866 1893 3869 1916
rect 3874 1896 3877 1946
rect 3882 1933 3885 2003
rect 3890 1936 3893 1986
rect 3906 1946 3909 2126
rect 3914 1993 3917 2133
rect 3922 2113 3925 2136
rect 3930 2133 3941 2136
rect 3930 2093 3933 2126
rect 3946 2073 3949 2136
rect 3954 2066 3957 2186
rect 3962 2143 3965 2166
rect 3946 2063 3957 2066
rect 3922 2003 3925 2046
rect 3946 2013 3949 2063
rect 3962 2013 3965 2136
rect 3970 2096 3973 2176
rect 3978 2113 3981 2126
rect 3970 2093 3977 2096
rect 3974 2006 3977 2093
rect 3898 1943 3909 1946
rect 3890 1933 3909 1936
rect 3890 1923 3901 1926
rect 3906 1916 3909 1926
rect 3914 1923 3917 1986
rect 3922 1923 3925 1936
rect 3938 1933 3941 1946
rect 3930 1923 3941 1926
rect 3906 1913 3917 1916
rect 3946 1913 3949 1966
rect 3954 1913 3957 2006
rect 3970 2003 3977 2006
rect 3962 1933 3965 1986
rect 3874 1893 3889 1896
rect 3866 1813 3869 1856
rect 3874 1803 3877 1886
rect 3886 1836 3889 1893
rect 3886 1833 3893 1836
rect 3866 1726 3869 1756
rect 3882 1753 3885 1816
rect 3890 1803 3893 1833
rect 3898 1813 3901 1856
rect 3898 1803 3909 1806
rect 3914 1796 3917 1913
rect 3962 1906 3965 1926
rect 3970 1923 3973 2003
rect 3978 1936 3981 1986
rect 3986 1946 3989 2196
rect 3998 2186 4001 2253
rect 3998 2183 4005 2186
rect 3994 2143 3997 2166
rect 3994 2103 3997 2136
rect 4002 2043 4005 2183
rect 4018 2156 4021 2386
rect 4026 2223 4029 2413
rect 4034 2383 4037 2423
rect 4034 2186 4037 2236
rect 4010 2153 4021 2156
rect 4026 2183 4037 2186
rect 4042 2186 4045 2523
rect 4050 2506 4053 2626
rect 4058 2613 4061 2626
rect 4058 2533 4061 2606
rect 4066 2536 4069 2633
rect 4074 2543 4077 2683
rect 4098 2613 4101 2686
rect 4106 2606 4109 2726
rect 4122 2723 4133 2726
rect 4082 2603 4093 2606
rect 4098 2603 4109 2606
rect 4098 2583 4101 2603
rect 4106 2573 4109 2596
rect 4114 2583 4117 2606
rect 4082 2543 4093 2546
rect 4066 2533 4077 2536
rect 4074 2523 4077 2533
rect 4082 2523 4085 2536
rect 4050 2503 4061 2506
rect 4058 2446 4061 2503
rect 4050 2443 4061 2446
rect 4050 2403 4053 2443
rect 4082 2433 4085 2516
rect 4090 2506 4093 2536
rect 4098 2523 4101 2566
rect 4114 2533 4117 2566
rect 4090 2503 4097 2506
rect 4094 2446 4097 2503
rect 4090 2443 4097 2446
rect 4090 2426 4093 2443
rect 4066 2413 4069 2426
rect 4082 2423 4093 2426
rect 4050 2383 4053 2396
rect 4050 2296 4053 2366
rect 4058 2313 4061 2326
rect 4066 2323 4069 2406
rect 4074 2393 4077 2406
rect 4074 2343 4077 2356
rect 4050 2293 4061 2296
rect 4058 2236 4061 2293
rect 4074 2243 4077 2336
rect 4082 2306 4085 2423
rect 4106 2416 4109 2526
rect 4122 2516 4125 2706
rect 4130 2626 4133 2723
rect 4138 2686 4141 2726
rect 4146 2723 4149 2756
rect 4154 2723 4157 2736
rect 4138 2683 4149 2686
rect 4130 2623 4141 2626
rect 4118 2513 4125 2516
rect 4118 2436 4121 2513
rect 4130 2466 4133 2616
rect 4138 2513 4141 2623
rect 4146 2553 4149 2683
rect 4154 2583 4157 2616
rect 4162 2603 4165 2793
rect 4186 2743 4189 2956
rect 4202 2936 4205 2963
rect 4202 2933 4221 2936
rect 4202 2846 4205 2926
rect 4210 2896 4213 2926
rect 4218 2903 4221 2926
rect 4234 2913 4237 2936
rect 4242 2896 4245 2976
rect 4250 2953 4253 3106
rect 4274 3013 4277 3026
rect 4250 2926 4253 2936
rect 4258 2933 4269 2936
rect 4250 2923 4261 2926
rect 4210 2893 4245 2896
rect 4202 2843 4221 2846
rect 4210 2793 4213 2816
rect 4178 2646 4181 2736
rect 4186 2663 4189 2736
rect 4194 2733 4205 2736
rect 4210 2733 4213 2756
rect 4178 2643 4189 2646
rect 4170 2593 4173 2626
rect 4186 2603 4189 2643
rect 4146 2533 4149 2546
rect 4170 2533 4173 2576
rect 4194 2543 4197 2716
rect 4202 2656 4205 2726
rect 4202 2653 4213 2656
rect 4210 2613 4213 2653
rect 4218 2633 4221 2843
rect 4226 2703 4229 2886
rect 4266 2883 4269 2933
rect 4234 2776 4237 2866
rect 4234 2773 4245 2776
rect 4266 2773 4269 2816
rect 4202 2593 4205 2606
rect 4218 2583 4221 2606
rect 4226 2556 4229 2666
rect 4242 2636 4245 2773
rect 4266 2723 4269 2736
rect 4274 2713 4277 2906
rect 4234 2633 4245 2636
rect 4234 2576 4237 2633
rect 4250 2583 4253 2606
rect 4274 2593 4277 2616
rect 4234 2573 4257 2576
rect 4210 2553 4229 2556
rect 4210 2536 4213 2553
rect 4146 2513 4149 2526
rect 4130 2463 4141 2466
rect 4118 2433 4125 2436
rect 4122 2416 4125 2433
rect 4138 2426 4141 2463
rect 4130 2423 4141 2426
rect 4090 2413 4109 2416
rect 4090 2403 4093 2413
rect 4106 2383 4109 2406
rect 4114 2366 4117 2416
rect 4122 2413 4129 2416
rect 4090 2323 4093 2336
rect 4098 2333 4101 2366
rect 4106 2363 4117 2366
rect 4082 2303 4089 2306
rect 4058 2233 4077 2236
rect 4074 2213 4077 2233
rect 4086 2226 4089 2303
rect 4082 2223 4089 2226
rect 4050 2193 4053 2206
rect 4058 2193 4069 2196
rect 4042 2183 4077 2186
rect 4010 2126 4013 2153
rect 4018 2133 4021 2146
rect 4010 2123 4021 2126
rect 4026 2123 4029 2183
rect 4034 2173 4061 2176
rect 4018 2053 4021 2123
rect 4034 2113 4037 2173
rect 4042 2083 4045 2126
rect 4050 2066 4053 2136
rect 4058 2123 4061 2173
rect 4066 2083 4069 2136
rect 4074 2123 4077 2183
rect 4082 2076 4085 2223
rect 4090 2173 4093 2206
rect 4098 2183 4101 2326
rect 4106 2293 4109 2363
rect 4114 2333 4117 2356
rect 4126 2346 4129 2413
rect 4138 2403 4141 2416
rect 4146 2396 4149 2506
rect 4154 2403 4157 2526
rect 4162 2433 4165 2526
rect 4178 2513 4181 2526
rect 4186 2503 4189 2536
rect 4194 2533 4213 2536
rect 4218 2533 4221 2546
rect 4162 2413 4181 2416
rect 4170 2396 4173 2406
rect 4146 2393 4173 2396
rect 4126 2343 4133 2346
rect 4114 2323 4125 2326
rect 4106 2193 4109 2206
rect 4114 2143 4117 2323
rect 4130 2316 4133 2343
rect 4138 2323 4141 2376
rect 4146 2333 4149 2356
rect 4122 2313 4133 2316
rect 4122 2203 4125 2313
rect 4130 2213 4133 2296
rect 4130 2173 4133 2206
rect 4098 2123 4101 2136
rect 4046 2063 4053 2066
rect 4058 2073 4085 2076
rect 3994 2003 3997 2016
rect 4010 2003 4013 2026
rect 4034 2003 4037 2016
rect 4046 2006 4049 2063
rect 4042 2003 4049 2006
rect 3994 1973 4037 1976
rect 3994 1956 3997 1973
rect 3994 1953 4005 1956
rect 3986 1943 3997 1946
rect 3978 1933 3989 1936
rect 3978 1923 3989 1926
rect 3978 1916 3981 1923
rect 3930 1903 3965 1906
rect 3970 1913 3981 1916
rect 3930 1836 3933 1903
rect 3930 1833 3941 1836
rect 3938 1813 3941 1833
rect 3922 1803 3941 1806
rect 3858 1723 3869 1726
rect 3874 1723 3877 1746
rect 3794 1483 3797 1516
rect 3810 1506 3813 1526
rect 3818 1513 3821 1546
rect 3826 1516 3829 1606
rect 3834 1533 3837 1606
rect 3842 1573 3845 1606
rect 3826 1513 3833 1516
rect 3810 1503 3821 1506
rect 3786 1403 3789 1426
rect 3794 1403 3797 1436
rect 3818 1413 3821 1503
rect 3830 1406 3833 1513
rect 3842 1453 3845 1536
rect 3850 1533 3853 1616
rect 3858 1526 3861 1723
rect 3882 1713 3885 1736
rect 3890 1723 3893 1776
rect 3898 1656 3901 1796
rect 3874 1653 3901 1656
rect 3906 1793 3917 1796
rect 3922 1793 3941 1796
rect 3874 1603 3877 1653
rect 3898 1613 3901 1626
rect 3850 1523 3861 1526
rect 3850 1496 3853 1523
rect 3866 1516 3869 1526
rect 3874 1523 3877 1536
rect 3882 1516 3885 1536
rect 3898 1533 3901 1586
rect 3890 1523 3901 1526
rect 3866 1513 3885 1516
rect 3890 1496 3893 1516
rect 3850 1493 3861 1496
rect 3858 1426 3861 1493
rect 3850 1423 3861 1426
rect 3882 1493 3893 1496
rect 3882 1426 3885 1493
rect 3882 1423 3893 1426
rect 3898 1423 3901 1523
rect 3906 1486 3909 1793
rect 3914 1753 3917 1786
rect 3914 1723 3917 1736
rect 3914 1503 3917 1686
rect 3922 1583 3925 1793
rect 3930 1706 3933 1786
rect 3946 1743 3949 1896
rect 3970 1883 3973 1913
rect 3986 1906 3989 1916
rect 3978 1903 3989 1906
rect 3978 1893 3981 1903
rect 3962 1746 3965 1806
rect 3986 1773 3989 1816
rect 3994 1753 3997 1943
rect 4002 1866 4005 1953
rect 4010 1886 4013 1966
rect 4026 1923 4029 1936
rect 4034 1933 4037 1973
rect 4026 1893 4029 1916
rect 4010 1883 4029 1886
rect 4002 1863 4009 1866
rect 4006 1806 4009 1863
rect 4002 1803 4009 1806
rect 4002 1783 4005 1803
rect 3962 1743 3981 1746
rect 3930 1703 3941 1706
rect 3938 1576 3941 1703
rect 3946 1653 3949 1736
rect 3970 1713 3973 1726
rect 3978 1703 3981 1743
rect 3922 1573 3941 1576
rect 3954 1573 3957 1616
rect 3906 1483 3913 1486
rect 3810 1366 3813 1406
rect 3826 1403 3833 1406
rect 3826 1376 3829 1403
rect 3802 1363 3813 1366
rect 3822 1373 3829 1376
rect 3786 1323 3789 1356
rect 3802 1323 3805 1363
rect 3794 1216 3797 1226
rect 3794 1213 3813 1216
rect 3786 1133 3789 1206
rect 3802 1193 3805 1206
rect 3810 1183 3813 1206
rect 3822 1146 3825 1373
rect 3842 1366 3845 1406
rect 3834 1363 3845 1366
rect 3834 1323 3837 1363
rect 3834 1173 3837 1276
rect 3794 1143 3825 1146
rect 3786 1103 3789 1126
rect 3794 1053 3797 1143
rect 3778 983 3781 1026
rect 3786 993 3789 1016
rect 3802 986 3805 1126
rect 3810 1103 3813 1126
rect 3818 1073 3821 1136
rect 3818 1013 3821 1066
rect 3826 1026 3829 1126
rect 3834 1093 3837 1136
rect 3842 1123 3845 1336
rect 3850 1296 3853 1423
rect 3858 1393 3861 1406
rect 3890 1403 3893 1423
rect 3898 1383 3901 1416
rect 3910 1376 3913 1483
rect 3906 1373 3913 1376
rect 3858 1323 3893 1326
rect 3858 1313 3861 1323
rect 3850 1293 3857 1296
rect 3854 1226 3857 1293
rect 3898 1283 3901 1316
rect 3850 1223 3857 1226
rect 3866 1243 3901 1246
rect 3850 1143 3853 1223
rect 3866 1213 3869 1243
rect 3858 1183 3861 1206
rect 3850 1123 3853 1136
rect 3858 1116 3861 1176
rect 3874 1143 3877 1216
rect 3890 1213 3893 1226
rect 3882 1183 3885 1206
rect 3898 1203 3901 1243
rect 3906 1196 3909 1373
rect 3922 1353 3925 1573
rect 3962 1566 3965 1586
rect 3946 1563 3965 1566
rect 3930 1533 3941 1536
rect 3930 1423 3933 1533
rect 3938 1513 3941 1526
rect 3946 1523 3949 1563
rect 3962 1483 3965 1536
rect 3970 1413 3973 1606
rect 3986 1603 3989 1656
rect 3978 1533 3981 1576
rect 3978 1463 3981 1526
rect 3986 1446 3989 1596
rect 4010 1576 4013 1616
rect 3994 1573 4013 1576
rect 3994 1533 3997 1573
rect 4002 1523 4005 1566
rect 4010 1513 4013 1536
rect 3982 1443 3989 1446
rect 3914 1303 3917 1336
rect 3914 1213 3917 1296
rect 3922 1233 3925 1336
rect 3930 1323 3933 1406
rect 3946 1326 3949 1406
rect 3946 1323 3957 1326
rect 3946 1283 3949 1316
rect 3954 1266 3957 1323
rect 3962 1306 3965 1376
rect 3982 1366 3985 1443
rect 3982 1363 3989 1366
rect 3970 1323 3973 1336
rect 3962 1303 3969 1306
rect 3950 1263 3957 1266
rect 3938 1213 3941 1226
rect 3898 1193 3909 1196
rect 3914 1193 3917 1206
rect 3930 1193 3933 1206
rect 3866 1123 3869 1136
rect 3842 1113 3861 1116
rect 3826 1023 3837 1026
rect 3790 983 3805 986
rect 3762 793 3765 836
rect 3770 813 3773 826
rect 3778 733 3781 936
rect 3790 846 3793 983
rect 3810 966 3813 1006
rect 3826 993 3829 1006
rect 3802 963 3813 966
rect 3802 923 3805 963
rect 3786 843 3793 846
rect 3762 713 3773 716
rect 3786 666 3789 843
rect 3802 826 3805 906
rect 3794 823 3805 826
rect 3794 753 3797 823
rect 3802 793 3805 806
rect 3818 803 3821 976
rect 3826 973 3837 976
rect 3826 813 3829 973
rect 3834 923 3837 966
rect 3842 903 3845 1113
rect 3874 1073 3877 1136
rect 3834 736 3837 806
rect 3842 783 3845 816
rect 3850 766 3853 1036
rect 3858 973 3861 1056
rect 3866 1013 3869 1026
rect 3882 936 3885 1126
rect 3890 1123 3893 1136
rect 3898 1113 3901 1193
rect 3950 1186 3953 1263
rect 3966 1246 3969 1303
rect 3966 1243 3973 1246
rect 3906 1183 3953 1186
rect 3890 1003 3893 1026
rect 3858 933 3885 936
rect 3858 913 3861 933
rect 3866 923 3877 926
rect 3874 913 3885 916
rect 3858 803 3861 866
rect 3866 773 3869 906
rect 3874 903 3893 906
rect 3898 903 3901 1076
rect 3906 1013 3909 1183
rect 3962 1176 3965 1236
rect 3914 1073 3917 1176
rect 3922 1173 3965 1176
rect 3970 1173 3973 1243
rect 3922 1123 3925 1173
rect 3978 1166 3981 1346
rect 3986 1263 3989 1363
rect 3994 1333 3997 1446
rect 3994 1303 3997 1326
rect 4010 1283 4013 1346
rect 4018 1306 4021 1776
rect 4026 1613 4029 1883
rect 4026 1503 4029 1536
rect 4034 1443 4037 1926
rect 4042 1763 4045 2003
rect 4050 1803 4053 1996
rect 4058 1976 4061 2073
rect 4058 1973 4069 1976
rect 4066 1933 4069 1973
rect 4058 1843 4061 1926
rect 4074 1893 4077 2046
rect 4082 2013 4093 2016
rect 4098 2003 4101 2116
rect 4106 2066 4109 2086
rect 4106 2063 4113 2066
rect 4082 1923 4085 1996
rect 4110 1986 4113 2063
rect 4122 1996 4125 2126
rect 4138 2043 4141 2306
rect 4154 2283 4157 2336
rect 4146 2176 4149 2246
rect 4162 2203 4165 2336
rect 4178 2323 4181 2406
rect 4186 2393 4189 2406
rect 4194 2356 4197 2533
rect 4202 2403 4205 2526
rect 4210 2523 4213 2533
rect 4234 2526 4237 2536
rect 4242 2533 4245 2566
rect 4218 2506 4221 2526
rect 4214 2503 4221 2506
rect 4214 2436 4217 2503
rect 4226 2446 4229 2526
rect 4234 2523 4245 2526
rect 4242 2513 4245 2523
rect 4254 2496 4257 2573
rect 4266 2506 4269 2586
rect 4266 2503 4273 2506
rect 4254 2493 4261 2496
rect 4226 2443 4237 2446
rect 4214 2433 4221 2436
rect 4210 2396 4213 2416
rect 4218 2403 4221 2433
rect 4226 2403 4229 2426
rect 4234 2413 4237 2443
rect 4242 2396 4245 2406
rect 4210 2393 4245 2396
rect 4194 2353 4213 2356
rect 4186 2213 4189 2336
rect 4194 2283 4197 2326
rect 4202 2293 4205 2336
rect 4210 2263 4213 2353
rect 4218 2333 4221 2376
rect 4234 2333 4237 2346
rect 4250 2326 4253 2436
rect 4258 2386 4261 2493
rect 4270 2446 4273 2503
rect 4282 2466 4285 2746
rect 4290 2676 4293 2946
rect 4314 2913 4317 2926
rect 4314 2803 4317 2816
rect 4330 2766 4333 3016
rect 4370 2883 4373 2926
rect 4370 2783 4373 2816
rect 4322 2763 4333 2766
rect 4322 2746 4325 2763
rect 4314 2743 4325 2746
rect 4290 2673 4297 2676
rect 4294 2606 4297 2673
rect 4314 2656 4317 2743
rect 4338 2713 4341 2726
rect 4314 2653 4325 2656
rect 4290 2603 4297 2606
rect 4290 2583 4293 2603
rect 4306 2523 4309 2546
rect 4322 2516 4325 2653
rect 4338 2613 4341 2626
rect 4362 2576 4365 2646
rect 4318 2513 4325 2516
rect 4354 2573 4365 2576
rect 4354 2516 4357 2573
rect 4370 2523 4373 2566
rect 4354 2513 4365 2516
rect 4282 2463 4309 2466
rect 4270 2443 4277 2446
rect 4258 2383 4269 2386
rect 4258 2333 4261 2366
rect 4242 2286 4245 2326
rect 4250 2323 4261 2326
rect 4266 2306 4269 2383
rect 4274 2333 4277 2443
rect 4298 2413 4301 2426
rect 4306 2396 4309 2463
rect 4290 2393 4309 2396
rect 4290 2333 4293 2393
rect 4318 2376 4321 2513
rect 4354 2393 4357 2416
rect 4314 2373 4321 2376
rect 4314 2356 4317 2373
rect 4306 2353 4317 2356
rect 4314 2323 4317 2346
rect 4266 2303 4285 2306
rect 4234 2283 4245 2286
rect 4146 2173 4169 2176
rect 4146 2063 4149 2096
rect 4166 2046 4169 2173
rect 4178 2113 4181 2126
rect 4166 2043 4173 2046
rect 4130 2023 4165 2026
rect 4130 2013 4133 2023
rect 4138 2013 4149 2016
rect 4130 2003 4141 2006
rect 4146 1996 4149 2006
rect 4122 1993 4149 1996
rect 4106 1983 4113 1986
rect 4154 1983 4157 2016
rect 4162 2003 4165 2023
rect 4170 1993 4173 2043
rect 4178 2003 4181 2096
rect 4090 1923 4093 1936
rect 4098 1923 4101 1956
rect 4106 1943 4109 1983
rect 4114 1963 4149 1966
rect 4114 1936 4117 1963
rect 4106 1933 4117 1936
rect 4058 1786 4061 1836
rect 4074 1803 4077 1856
rect 4058 1783 4069 1786
rect 4042 1713 4045 1726
rect 4050 1553 4053 1726
rect 4042 1523 4045 1546
rect 4042 1513 4053 1516
rect 4042 1473 4045 1513
rect 4026 1413 4029 1426
rect 4034 1333 4037 1416
rect 4042 1393 4045 1406
rect 4026 1323 4037 1326
rect 4018 1303 4025 1306
rect 3994 1203 3997 1246
rect 4022 1236 4025 1303
rect 4018 1233 4025 1236
rect 3962 1163 3981 1166
rect 3930 1036 3933 1136
rect 3938 1113 3941 1126
rect 3946 1123 3949 1136
rect 3954 1106 3957 1156
rect 3962 1146 3965 1163
rect 3962 1143 3973 1146
rect 3946 1103 3957 1106
rect 3962 1103 3965 1136
rect 3970 1106 3973 1143
rect 3978 1113 3981 1126
rect 3994 1113 3997 1136
rect 4002 1133 4013 1136
rect 3970 1103 3997 1106
rect 3946 1053 3949 1103
rect 3922 1033 3933 1036
rect 3874 803 3877 816
rect 3882 803 3885 846
rect 3850 763 3885 766
rect 3802 733 3837 736
rect 3778 663 3789 666
rect 3754 633 3765 636
rect 3690 573 3693 606
rect 3698 566 3701 606
rect 3690 563 3701 566
rect 3690 533 3693 563
rect 3674 503 3685 506
rect 3682 446 3685 503
rect 3682 443 3693 446
rect 3666 423 3685 426
rect 3666 413 3669 423
rect 3650 403 3661 406
rect 3634 333 3637 346
rect 3626 313 3629 326
rect 3642 296 3645 386
rect 3634 293 3645 296
rect 3634 206 3637 293
rect 3650 213 3653 336
rect 3658 323 3661 403
rect 3674 343 3677 416
rect 3682 403 3685 423
rect 3682 316 3685 386
rect 3674 313 3685 316
rect 3674 236 3677 313
rect 3674 233 3685 236
rect 3682 213 3685 233
rect 3690 213 3693 443
rect 3698 403 3701 456
rect 3706 403 3709 416
rect 3714 396 3717 633
rect 3722 603 3725 626
rect 3706 393 3717 396
rect 3706 383 3709 393
rect 3722 386 3725 586
rect 3730 463 3733 633
rect 3738 593 3741 606
rect 3746 583 3749 606
rect 3738 486 3741 526
rect 3738 483 3749 486
rect 3738 413 3741 436
rect 3746 403 3749 483
rect 3754 433 3757 616
rect 3762 613 3765 633
rect 3778 613 3781 663
rect 3786 593 3789 606
rect 3770 573 3781 576
rect 3770 523 3773 536
rect 3762 496 3765 516
rect 3778 506 3781 573
rect 3794 523 3797 616
rect 3802 603 3805 726
rect 3834 713 3837 733
rect 3810 596 3813 656
rect 3802 593 3813 596
rect 3778 503 3789 506
rect 3762 493 3769 496
rect 3766 426 3769 493
rect 3762 423 3769 426
rect 3754 393 3757 416
rect 3762 403 3765 423
rect 3714 383 3725 386
rect 3698 333 3709 336
rect 3714 323 3717 383
rect 3722 333 3725 366
rect 3730 316 3733 386
rect 3770 363 3773 406
rect 3770 333 3773 346
rect 3714 313 3733 316
rect 3722 213 3725 313
rect 3762 263 3765 326
rect 3762 213 3765 256
rect 3490 163 3541 166
rect 3546 163 3597 166
rect 3538 123 3541 163
rect 3570 133 3573 146
rect 3594 123 3597 163
rect 3602 143 3605 206
rect 3634 203 3653 206
rect 3650 123 3653 203
rect 3706 153 3709 206
rect 3738 203 3749 206
rect 3754 196 3757 206
rect 3770 203 3773 236
rect 3778 223 3781 496
rect 3786 363 3789 503
rect 3802 433 3805 593
rect 3818 533 3821 606
rect 3842 603 3845 686
rect 3858 643 3861 736
rect 3866 593 3869 616
rect 3818 483 3821 516
rect 3786 333 3789 356
rect 3730 193 3757 196
rect 3794 193 3797 416
rect 3802 316 3805 396
rect 3810 346 3813 416
rect 3826 413 3829 536
rect 3842 416 3845 526
rect 3858 523 3869 526
rect 3874 523 3877 666
rect 3866 513 3869 523
rect 3882 506 3885 763
rect 3878 503 3885 506
rect 3878 436 3881 503
rect 3866 416 3869 436
rect 3878 433 3885 436
rect 3842 413 3861 416
rect 3866 413 3873 416
rect 3818 396 3821 406
rect 3818 393 3845 396
rect 3850 353 3853 406
rect 3858 373 3861 413
rect 3870 366 3873 413
rect 3866 363 3873 366
rect 3810 343 3837 346
rect 3802 313 3813 316
rect 3810 246 3813 313
rect 3826 303 3829 336
rect 3802 243 3813 246
rect 3802 226 3805 243
rect 3802 223 3829 226
rect 3810 213 3821 216
rect 3826 213 3829 223
rect 3682 133 3685 146
rect 3730 123 3733 193
rect 3762 123 3765 156
rect 3818 146 3821 206
rect 3834 203 3837 343
rect 3850 333 3853 346
rect 3866 316 3869 363
rect 3882 333 3885 433
rect 3890 403 3893 903
rect 3906 863 3909 1006
rect 3914 973 3917 1016
rect 3922 933 3925 1033
rect 3930 1013 3933 1026
rect 3914 913 3917 926
rect 3922 923 3933 926
rect 3898 763 3901 816
rect 3906 746 3909 836
rect 3914 766 3917 856
rect 3930 803 3933 896
rect 3938 843 3941 1006
rect 3938 803 3941 816
rect 3914 763 3941 766
rect 3898 743 3909 746
rect 3898 716 3901 743
rect 3906 723 3909 736
rect 3898 713 3909 716
rect 3906 656 3909 713
rect 3906 653 3913 656
rect 3910 596 3913 653
rect 3922 613 3925 716
rect 3930 606 3933 746
rect 3938 723 3941 763
rect 3946 706 3949 976
rect 3942 703 3949 706
rect 3942 636 3945 703
rect 3906 593 3913 596
rect 3922 603 3933 606
rect 3938 633 3945 636
rect 3906 576 3909 593
rect 3898 573 3909 576
rect 3898 513 3901 573
rect 3906 533 3909 546
rect 3906 473 3909 526
rect 3914 493 3917 536
rect 3922 523 3925 603
rect 3938 553 3941 633
rect 3954 613 3957 1096
rect 3970 1076 3973 1096
rect 3966 1073 3973 1076
rect 3966 976 3969 1073
rect 3978 1003 3981 1076
rect 3986 1013 3989 1046
rect 3994 1003 3997 1103
rect 4002 1053 4005 1126
rect 4018 1093 4021 1233
rect 4026 1193 4029 1216
rect 4026 1086 4029 1146
rect 4034 1106 4037 1286
rect 4042 1133 4045 1356
rect 4050 1333 4053 1456
rect 4058 1133 4061 1736
rect 4066 1723 4069 1783
rect 4082 1723 4085 1756
rect 4090 1733 4093 1786
rect 4098 1726 4101 1756
rect 4090 1723 4101 1726
rect 4090 1716 4093 1723
rect 4082 1713 4093 1716
rect 4106 1713 4109 1846
rect 4114 1773 4117 1926
rect 4122 1813 4125 1936
rect 4130 1923 4133 1936
rect 4138 1933 4141 1956
rect 4146 1933 4149 1963
rect 4146 1843 4149 1926
rect 4146 1786 4149 1836
rect 4154 1813 4157 1926
rect 4162 1896 4165 1936
rect 4170 1916 4173 1936
rect 4178 1923 4181 1976
rect 4186 1933 4189 2106
rect 4194 2023 4197 2216
rect 4210 2176 4213 2226
rect 4242 2176 4245 2216
rect 4258 2193 4261 2206
rect 4210 2173 4221 2176
rect 4234 2173 4245 2176
rect 4218 2063 4221 2173
rect 4226 2106 4229 2126
rect 4226 2103 4237 2106
rect 4234 2046 4237 2103
rect 4226 2043 4237 2046
rect 4194 1953 4197 2016
rect 4210 2013 4213 2026
rect 4202 2003 4213 2006
rect 4218 1973 4221 2016
rect 4226 2003 4229 2043
rect 4234 2023 4245 2026
rect 4194 1923 4197 1936
rect 4202 1933 4205 1946
rect 4210 1916 4213 1936
rect 4170 1913 4213 1916
rect 4162 1893 4169 1896
rect 4166 1826 4169 1893
rect 4162 1823 4169 1826
rect 4162 1806 4165 1823
rect 4178 1813 4181 1846
rect 4186 1816 4189 1913
rect 4218 1826 4221 1966
rect 4234 1946 4237 2016
rect 4242 2003 4245 2023
rect 4250 1963 4253 2016
rect 4234 1943 4253 1946
rect 4226 1913 4229 1936
rect 4234 1923 4237 1936
rect 4242 1863 4245 1936
rect 4250 1833 4253 1943
rect 4258 1853 4261 2126
rect 4266 2083 4269 2216
rect 4282 2203 4285 2303
rect 4354 2276 4357 2326
rect 4350 2273 4357 2276
rect 4274 2093 4277 2126
rect 4266 2003 4277 2006
rect 4266 1893 4269 1936
rect 4266 1846 4269 1886
rect 4258 1843 4269 1846
rect 4258 1826 4261 1843
rect 4274 1836 4277 2003
rect 4282 1983 4285 2066
rect 4290 1856 4293 2156
rect 4314 2086 4317 2126
rect 4322 2103 4325 2216
rect 4350 2176 4353 2273
rect 4350 2173 4357 2176
rect 4298 2083 4317 2086
rect 4298 2003 4301 2083
rect 4322 2026 4325 2056
rect 4338 2036 4341 2146
rect 4338 2033 4345 2036
rect 4322 2023 4333 2026
rect 4306 1993 4309 2016
rect 4314 2013 4325 2016
rect 4314 2003 4317 2013
rect 4322 1993 4325 2006
rect 4314 1913 4317 1926
rect 4202 1823 4221 1826
rect 4250 1823 4261 1826
rect 4266 1833 4277 1836
rect 4282 1853 4293 1856
rect 4186 1813 4197 1816
rect 4202 1813 4205 1823
rect 4162 1803 4189 1806
rect 4162 1786 4165 1796
rect 4146 1783 4165 1786
rect 4114 1733 4117 1746
rect 4130 1733 4133 1766
rect 4138 1733 4141 1756
rect 4122 1723 4141 1726
rect 4066 1613 4069 1686
rect 4074 1593 4077 1616
rect 4082 1546 4085 1713
rect 4122 1706 4125 1723
rect 4118 1703 4125 1706
rect 4118 1636 4121 1703
rect 4118 1633 4125 1636
rect 4122 1616 4125 1633
rect 4106 1613 4125 1616
rect 4090 1603 4101 1606
rect 4106 1556 4109 1613
rect 4114 1583 4117 1606
rect 4130 1603 4133 1696
rect 4122 1576 4125 1596
rect 4098 1553 4109 1556
rect 4114 1573 4125 1576
rect 4066 1543 4085 1546
rect 4066 1533 4069 1543
rect 4074 1534 4085 1537
rect 4090 1533 4093 1546
rect 4066 1423 4069 1526
rect 4074 1343 4077 1486
rect 4082 1443 4085 1526
rect 4098 1413 4101 1553
rect 4114 1416 4117 1573
rect 4138 1556 4141 1716
rect 4146 1563 4149 1783
rect 4186 1773 4189 1803
rect 4162 1703 4165 1736
rect 4186 1723 4189 1746
rect 4154 1613 4157 1626
rect 4154 1573 4157 1606
rect 4138 1553 4149 1556
rect 4138 1523 4141 1536
rect 4114 1413 4125 1416
rect 4130 1413 4133 1466
rect 4090 1356 4093 1406
rect 4090 1353 4101 1356
rect 4074 1323 4077 1336
rect 4098 1323 4101 1353
rect 4106 1333 4109 1406
rect 4114 1343 4117 1406
rect 4122 1323 4125 1413
rect 4066 1186 4069 1216
rect 4074 1213 4077 1236
rect 4066 1183 4077 1186
rect 4050 1123 4061 1126
rect 4034 1103 4045 1106
rect 4018 1083 4029 1086
rect 4018 1036 4021 1083
rect 4042 1046 4045 1103
rect 4002 1003 4005 1036
rect 4014 1033 4021 1036
rect 4034 1043 4045 1046
rect 4014 976 4017 1033
rect 4026 1013 4029 1026
rect 4034 1013 4037 1043
rect 4066 1026 4069 1146
rect 4074 1096 4077 1183
rect 4090 1173 4093 1206
rect 4114 1183 4117 1216
rect 4122 1176 4125 1266
rect 4106 1173 4125 1176
rect 4082 1113 4085 1126
rect 4090 1103 4093 1136
rect 4074 1093 4093 1096
rect 4050 1023 4069 1026
rect 3966 973 3973 976
rect 4014 973 4021 976
rect 3970 956 3973 973
rect 3962 916 3965 956
rect 3970 953 4013 956
rect 3978 923 3981 946
rect 3986 923 4005 926
rect 3986 916 3989 923
rect 3962 913 3989 916
rect 4002 896 4005 916
rect 3994 893 4005 896
rect 3970 813 3973 846
rect 3994 826 3997 893
rect 3994 823 4001 826
rect 3962 733 3965 806
rect 3970 803 3981 806
rect 3986 753 3989 806
rect 3998 776 4001 823
rect 3998 773 4005 776
rect 4002 743 4005 773
rect 3986 673 3989 736
rect 4010 656 4013 953
rect 4018 933 4021 973
rect 3994 653 4013 656
rect 3954 593 3957 606
rect 3930 436 3933 536
rect 3938 523 3941 536
rect 3946 506 3949 546
rect 3898 433 3933 436
rect 3942 503 3949 506
rect 3890 333 3893 396
rect 3898 386 3901 433
rect 3942 426 3945 503
rect 3906 423 3925 426
rect 3906 413 3909 423
rect 3914 396 3917 416
rect 3922 403 3925 423
rect 3930 423 3945 426
rect 3930 413 3933 423
rect 3938 413 3941 423
rect 3946 396 3949 416
rect 3914 393 3949 396
rect 3898 383 3933 386
rect 3858 313 3869 316
rect 3906 316 3909 326
rect 3914 323 3917 336
rect 3922 316 3925 336
rect 3906 313 3925 316
rect 3858 226 3861 313
rect 3858 223 3869 226
rect 3842 193 3845 206
rect 3866 166 3869 223
rect 3874 206 3877 306
rect 3882 213 3885 256
rect 3898 213 3901 226
rect 3874 203 3885 206
rect 3866 163 3873 166
rect 3818 143 3829 146
rect 3802 123 3805 136
rect 3826 123 3829 143
rect 2490 113 2525 116
rect 3870 106 3873 163
rect 3882 123 3885 203
rect 3890 166 3893 206
rect 3906 203 3909 266
rect 3930 243 3933 383
rect 3938 383 3949 386
rect 3938 333 3941 383
rect 3946 306 3949 336
rect 3942 303 3949 306
rect 3954 303 3957 586
rect 3962 513 3965 536
rect 3962 403 3965 506
rect 3970 486 3973 576
rect 3978 493 3981 636
rect 3986 576 3989 646
rect 3994 583 3997 653
rect 4002 593 4005 616
rect 3986 573 3997 576
rect 4018 573 4021 926
rect 4026 596 4029 1006
rect 4034 943 4037 1006
rect 4050 996 4053 1023
rect 4058 1003 4061 1016
rect 4066 1003 4069 1016
rect 4082 1013 4085 1066
rect 4050 993 4061 996
rect 4034 913 4037 936
rect 4034 803 4037 816
rect 4042 803 4045 896
rect 4050 826 4053 976
rect 4058 933 4061 993
rect 4074 986 4077 1006
rect 4070 983 4077 986
rect 4082 983 4085 1006
rect 4058 833 4061 916
rect 4070 906 4073 983
rect 4070 903 4077 906
rect 4050 823 4061 826
rect 4058 796 4061 823
rect 4066 816 4069 846
rect 4074 826 4077 903
rect 4090 863 4093 1093
rect 4098 973 4101 1156
rect 4106 946 4109 1173
rect 4114 1133 4125 1136
rect 4114 1096 4117 1133
rect 4122 1116 4125 1126
rect 4130 1123 4133 1276
rect 4138 1153 4141 1516
rect 4146 1273 4149 1553
rect 4154 1453 4157 1556
rect 4162 1513 4165 1616
rect 4170 1613 4181 1616
rect 4170 1603 4181 1606
rect 4186 1603 4189 1626
rect 4194 1556 4197 1813
rect 4202 1753 4205 1806
rect 4226 1793 4229 1806
rect 4234 1723 4237 1816
rect 4242 1803 4245 1816
rect 4250 1796 4253 1823
rect 4258 1803 4261 1816
rect 4242 1793 4253 1796
rect 4242 1716 4245 1793
rect 4266 1776 4269 1833
rect 4282 1803 4285 1853
rect 4306 1793 4309 1816
rect 4314 1803 4317 1906
rect 4234 1713 4245 1716
rect 4250 1716 4253 1776
rect 4266 1773 4273 1776
rect 4258 1723 4261 1766
rect 4250 1713 4257 1716
rect 4210 1593 4213 1606
rect 4234 1566 4237 1713
rect 4254 1636 4257 1713
rect 4270 1706 4273 1773
rect 4290 1706 4293 1736
rect 4266 1703 4273 1706
rect 4282 1703 4293 1706
rect 4266 1656 4269 1703
rect 4266 1653 4277 1656
rect 4210 1563 4237 1566
rect 4194 1553 4205 1556
rect 4194 1503 4197 1526
rect 4170 1463 4181 1466
rect 4162 1413 4165 1426
rect 4178 1413 4181 1463
rect 4154 1403 4165 1406
rect 4154 1323 4157 1396
rect 4162 1386 4165 1403
rect 4178 1396 4181 1406
rect 4202 1403 4205 1553
rect 4210 1503 4213 1563
rect 4218 1416 4221 1556
rect 4242 1553 4245 1636
rect 4254 1633 4261 1636
rect 4250 1603 4253 1616
rect 4226 1513 4229 1536
rect 4258 1526 4261 1633
rect 4274 1573 4277 1653
rect 4282 1606 4285 1703
rect 4290 1613 4293 1696
rect 4314 1676 4317 1726
rect 4306 1673 4317 1676
rect 4306 1626 4309 1673
rect 4298 1623 4309 1626
rect 4282 1603 4293 1606
rect 4234 1523 4261 1526
rect 4266 1523 4269 1536
rect 4210 1413 4221 1416
rect 4226 1413 4229 1446
rect 4178 1393 4197 1396
rect 4162 1383 4189 1386
rect 4170 1283 4173 1336
rect 4178 1306 4181 1356
rect 4186 1316 4189 1383
rect 4194 1323 4197 1393
rect 4202 1333 4205 1346
rect 4210 1326 4213 1413
rect 4218 1393 4221 1406
rect 4218 1333 4221 1346
rect 4210 1323 4221 1326
rect 4226 1323 4229 1406
rect 4234 1396 4237 1506
rect 4242 1443 4245 1523
rect 4274 1493 4277 1526
rect 4290 1456 4293 1603
rect 4298 1593 4301 1623
rect 4322 1616 4325 1986
rect 4330 1633 4333 2023
rect 4342 1976 4345 2033
rect 4338 1973 4345 1976
rect 4338 1856 4341 1973
rect 4338 1853 4349 1856
rect 4346 1833 4349 1853
rect 4354 1826 4357 2173
rect 4346 1823 4357 1826
rect 4362 1826 4365 2513
rect 4370 2323 4373 2366
rect 4370 2193 4373 2216
rect 4370 2033 4373 2126
rect 4370 1883 4373 2026
rect 4378 1923 4381 2276
rect 4378 1893 4381 1916
rect 4362 1823 4373 1826
rect 4346 1783 4349 1823
rect 4354 1813 4365 1816
rect 4354 1776 4357 1806
rect 4338 1773 4357 1776
rect 4338 1676 4341 1773
rect 4370 1733 4373 1823
rect 4354 1723 4373 1726
rect 4338 1673 4345 1676
rect 4298 1573 4301 1586
rect 4306 1553 4309 1616
rect 4314 1613 4325 1616
rect 4330 1613 4333 1626
rect 4314 1586 4317 1613
rect 4322 1593 4325 1606
rect 4314 1583 4325 1586
rect 4314 1513 4317 1526
rect 4290 1453 4317 1456
rect 4242 1413 4245 1436
rect 4250 1403 4261 1406
rect 4234 1393 4241 1396
rect 4238 1316 4241 1393
rect 4250 1333 4261 1336
rect 4266 1323 4269 1386
rect 4282 1353 4285 1406
rect 4306 1393 4309 1416
rect 4186 1313 4213 1316
rect 4178 1303 4189 1306
rect 4162 1213 4173 1216
rect 4162 1163 4165 1213
rect 4186 1203 4189 1303
rect 4210 1266 4213 1313
rect 4234 1313 4241 1316
rect 4210 1263 4221 1266
rect 4218 1213 4221 1263
rect 4234 1256 4237 1313
rect 4230 1253 4237 1256
rect 4250 1256 4253 1296
rect 4282 1286 4285 1336
rect 4306 1323 4309 1346
rect 4314 1286 4317 1453
rect 4250 1253 4257 1256
rect 4230 1196 4233 1253
rect 4230 1193 4237 1196
rect 4146 1143 4165 1146
rect 4138 1123 4141 1136
rect 4146 1123 4149 1143
rect 4154 1116 4157 1136
rect 4122 1113 4157 1116
rect 4114 1093 4125 1096
rect 4122 1036 4125 1093
rect 4114 1033 4125 1036
rect 4114 983 4117 1033
rect 4146 1016 4149 1086
rect 4162 1016 4165 1143
rect 4186 1133 4189 1176
rect 4234 1173 4237 1193
rect 4218 1113 4221 1126
rect 4106 943 4117 946
rect 4114 886 4117 943
rect 4122 933 4125 1006
rect 4138 993 4141 1016
rect 4146 1013 4157 1016
rect 4162 1013 4173 1016
rect 4146 983 4149 1006
rect 4154 973 4157 1013
rect 4162 966 4165 1006
rect 4178 993 4181 1006
rect 4186 983 4189 1006
rect 4218 996 4221 1016
rect 4226 1003 4229 1166
rect 4254 1156 4257 1253
rect 4266 1213 4269 1286
rect 4282 1283 4317 1286
rect 4290 1183 4293 1283
rect 4250 1153 4257 1156
rect 4250 1076 4253 1153
rect 4246 1073 4253 1076
rect 4234 1013 4237 1056
rect 4246 996 4249 1073
rect 4258 1003 4261 1136
rect 4282 1133 4285 1176
rect 4314 1163 4317 1216
rect 4266 1103 4269 1126
rect 4218 993 4249 996
rect 4138 963 4165 966
rect 4138 923 4141 963
rect 4178 933 4181 946
rect 4186 926 4189 936
rect 4194 933 4213 936
rect 4178 923 4189 926
rect 4194 913 4197 926
rect 4110 883 4117 886
rect 4074 823 4101 826
rect 4066 813 4077 816
rect 4034 723 4037 796
rect 4054 793 4061 796
rect 4066 793 4069 806
rect 4082 803 4085 816
rect 4054 716 4057 793
rect 4090 763 4093 806
rect 4066 723 4069 756
rect 4098 746 4101 823
rect 4110 796 4113 883
rect 4122 803 4125 886
rect 4130 803 4133 816
rect 4110 793 4117 796
rect 4146 793 4149 816
rect 4162 813 4165 846
rect 4202 843 4205 926
rect 4210 886 4213 933
rect 4218 903 4221 993
rect 4226 956 4229 976
rect 4226 953 4237 956
rect 4210 883 4221 886
rect 4090 743 4101 746
rect 4054 713 4061 716
rect 4034 613 4037 696
rect 4058 643 4061 713
rect 4074 703 4077 736
rect 4090 636 4093 743
rect 4114 736 4117 793
rect 4106 733 4117 736
rect 4106 653 4109 733
rect 4114 666 4117 726
rect 4130 683 4133 736
rect 4154 723 4157 806
rect 4178 803 4181 816
rect 4186 803 4189 826
rect 4210 796 4213 816
rect 4218 803 4221 883
rect 4234 866 4237 953
rect 4250 933 4253 946
rect 4226 863 4237 866
rect 4226 803 4229 863
rect 4258 846 4261 966
rect 4266 913 4269 936
rect 4274 883 4277 1006
rect 4306 956 4309 1146
rect 4314 1003 4317 1126
rect 4322 1043 4325 1583
rect 4330 1076 4333 1606
rect 4342 1576 4345 1673
rect 4354 1603 4357 1723
rect 4362 1696 4365 1716
rect 4362 1693 4369 1696
rect 4366 1616 4369 1693
rect 4362 1613 4369 1616
rect 4362 1596 4365 1613
rect 4338 1573 4345 1576
rect 4354 1593 4365 1596
rect 4338 1486 4341 1573
rect 4354 1506 4357 1593
rect 4362 1523 4373 1526
rect 4354 1503 4365 1506
rect 4338 1483 4349 1486
rect 4346 1286 4349 1483
rect 4362 1436 4365 1503
rect 4354 1433 4365 1436
rect 4354 1373 4357 1433
rect 4362 1403 4365 1416
rect 4362 1323 4365 1336
rect 4378 1306 4381 1826
rect 4338 1283 4349 1286
rect 4370 1303 4381 1306
rect 4338 1176 4341 1283
rect 4370 1236 4373 1303
rect 4370 1233 4381 1236
rect 4338 1173 4349 1176
rect 4330 1073 4337 1076
rect 4322 963 4325 1016
rect 4334 976 4337 1073
rect 4346 1003 4349 1173
rect 4354 996 4357 1186
rect 4370 1136 4373 1216
rect 4362 1133 4373 1136
rect 4362 1103 4365 1126
rect 4370 1006 4373 1036
rect 4362 1003 4373 1006
rect 4354 993 4365 996
rect 4330 973 4337 976
rect 4306 953 4325 956
rect 4330 953 4333 973
rect 4242 843 4261 846
rect 4234 803 4237 816
rect 4242 813 4245 843
rect 4250 796 4253 806
rect 4178 766 4181 796
rect 4210 793 4253 796
rect 4170 763 4181 766
rect 4170 686 4173 763
rect 4210 723 4213 766
rect 4258 756 4261 786
rect 4250 753 4261 756
rect 4226 723 4229 736
rect 4250 706 4253 753
rect 4282 733 4285 866
rect 4290 853 4293 936
rect 4314 923 4317 946
rect 4306 813 4309 826
rect 4306 746 4309 806
rect 4306 743 4313 746
rect 4266 713 4269 726
rect 4250 703 4269 706
rect 4170 683 4189 686
rect 4114 663 4173 666
rect 4066 633 4093 636
rect 4026 593 4037 596
rect 3994 533 3997 573
rect 3970 483 3981 486
rect 3970 373 3973 406
rect 3978 366 3981 483
rect 3974 363 3981 366
rect 3942 226 3945 303
rect 3942 223 3949 226
rect 3946 206 3949 223
rect 3954 213 3957 256
rect 3962 213 3965 326
rect 3974 216 3977 363
rect 3970 213 3977 216
rect 3938 196 3941 206
rect 3946 203 3957 206
rect 3970 196 3973 213
rect 3986 203 3989 406
rect 3994 376 3997 416
rect 4002 413 4005 436
rect 4010 396 4013 496
rect 4018 403 4021 526
rect 4034 486 4037 593
rect 4034 483 4045 486
rect 4042 426 4045 483
rect 4058 433 4061 616
rect 4026 413 4029 426
rect 4042 423 4053 426
rect 4034 396 4037 406
rect 4010 393 4037 396
rect 4042 393 4045 406
rect 4050 386 4053 423
rect 4058 403 4061 416
rect 4034 383 4053 386
rect 3994 373 4013 376
rect 3994 333 3997 346
rect 4010 333 4013 373
rect 4034 366 4037 383
rect 4066 373 4069 633
rect 4074 413 4077 626
rect 4082 623 4117 626
rect 4082 613 4085 623
rect 4090 613 4101 616
rect 4082 586 4085 606
rect 4098 593 4101 606
rect 4106 603 4109 616
rect 4114 603 4117 623
rect 4122 613 4125 646
rect 4122 586 4125 606
rect 4154 593 4157 606
rect 4082 583 4125 586
rect 4090 533 4093 546
rect 4114 533 4117 576
rect 4122 563 4125 583
rect 4082 513 4085 526
rect 4082 403 4085 506
rect 4030 363 4037 366
rect 4002 213 4005 326
rect 3938 193 3981 196
rect 3890 163 3941 166
rect 3914 133 3917 156
rect 3938 123 3941 163
rect 3978 126 3981 193
rect 3994 143 3997 206
rect 4018 203 4021 336
rect 4030 306 4033 363
rect 4030 303 4037 306
rect 4034 183 4037 303
rect 4050 196 4053 336
rect 4074 323 4077 346
rect 4090 296 4093 426
rect 4098 403 4101 526
rect 4114 333 4117 526
rect 4138 503 4141 526
rect 4146 496 4149 566
rect 4138 493 4149 496
rect 4138 403 4141 493
rect 4146 413 4149 436
rect 4154 386 4157 556
rect 4162 486 4165 616
rect 4170 603 4173 663
rect 4186 636 4189 683
rect 4182 633 4189 636
rect 4182 536 4185 633
rect 4202 576 4205 676
rect 4266 656 4269 703
rect 4266 653 4273 656
rect 4226 593 4229 616
rect 4194 573 4205 576
rect 4182 533 4189 536
rect 4186 516 4189 533
rect 4194 523 4197 546
rect 4202 533 4205 566
rect 4226 533 4229 546
rect 4202 516 4205 526
rect 4234 523 4237 606
rect 4270 596 4273 653
rect 4282 613 4285 706
rect 4310 696 4313 743
rect 4306 693 4313 696
rect 4290 666 4293 686
rect 4290 663 4297 666
rect 4294 606 4297 663
rect 4306 613 4309 693
rect 4322 626 4325 953
rect 4354 876 4357 906
rect 4350 873 4357 876
rect 4350 736 4353 873
rect 4350 733 4357 736
rect 4314 623 4325 626
rect 4266 593 4273 596
rect 4290 603 4297 606
rect 4266 576 4269 593
rect 4258 573 4269 576
rect 4186 513 4205 516
rect 4162 483 4173 486
rect 4162 396 4165 406
rect 4170 403 4173 483
rect 4178 403 4181 436
rect 4186 413 4189 513
rect 4194 396 4197 416
rect 4234 413 4237 426
rect 4162 393 4189 396
rect 4194 393 4201 396
rect 4122 383 4157 386
rect 4074 293 4093 296
rect 4066 203 4069 216
rect 4074 203 4077 293
rect 4098 213 4101 246
rect 4122 213 4125 383
rect 4130 323 4133 376
rect 4162 306 4165 336
rect 4186 323 4189 393
rect 4198 316 4201 393
rect 4138 303 4165 306
rect 4194 313 4201 316
rect 4050 193 4069 196
rect 4034 133 4037 156
rect 3978 123 3997 126
rect 4058 123 4061 146
rect 4066 123 4069 193
rect 4106 143 4109 206
rect 4114 203 4125 206
rect 4114 123 4117 186
rect 4138 133 4141 303
rect 4194 253 4197 313
rect 4162 213 4165 236
rect 4154 146 4157 206
rect 4170 203 4173 246
rect 4178 213 4181 226
rect 4210 206 4213 406
rect 4226 393 4229 406
rect 4242 403 4245 466
rect 4242 323 4245 336
rect 4250 323 4253 566
rect 4258 513 4261 573
rect 4290 456 4293 603
rect 4306 563 4309 606
rect 4314 553 4317 623
rect 4322 586 4325 616
rect 4330 603 4333 726
rect 4338 603 4341 616
rect 4346 603 4349 716
rect 4322 583 4333 586
rect 4314 523 4317 546
rect 4282 453 4293 456
rect 4258 403 4261 426
rect 4266 313 4269 406
rect 4282 403 4285 453
rect 4306 393 4309 416
rect 4314 386 4317 506
rect 4330 466 4333 583
rect 4354 503 4357 733
rect 4362 696 4365 993
rect 4378 973 4381 1233
rect 4370 923 4373 936
rect 4370 813 4373 836
rect 4370 713 4373 726
rect 4362 693 4369 696
rect 4366 546 4369 693
rect 4362 543 4369 546
rect 4326 463 4333 466
rect 4326 406 4329 463
rect 4306 383 4317 386
rect 4322 403 4329 406
rect 4322 383 4325 403
rect 4234 213 4237 236
rect 4210 203 4221 206
rect 4226 193 4229 206
rect 4242 156 4245 256
rect 4282 166 4285 376
rect 4306 223 4309 383
rect 4362 373 4365 543
rect 4370 513 4373 526
rect 4370 413 4373 426
rect 4378 336 4381 926
rect 4314 296 4317 336
rect 4362 333 4381 336
rect 4322 313 4325 326
rect 4314 293 4325 296
rect 4322 236 4325 293
rect 4314 233 4325 236
rect 4314 213 4317 233
rect 4362 213 4365 333
rect 4274 163 4285 166
rect 4242 153 4253 156
rect 4154 143 4165 146
rect 4162 123 4165 143
rect 4218 123 4221 146
rect 4242 133 4245 146
rect 4250 123 4253 153
rect 4274 123 4277 163
rect 4298 123 4301 196
rect 4354 123 4357 146
rect 3866 103 3873 106
rect 3866 83 3869 103
rect 4390 37 4410 4303
rect 4414 13 4434 4327
rect 4442 1873 4445 2616
<< metal3 >>
rect 2113 4332 2766 4337
rect 2113 4327 2118 4332
rect 2089 4322 2118 4327
rect 2761 4327 2766 4332
rect 2977 4332 3958 4337
rect 2977 4327 2982 4332
rect 2761 4322 2790 4327
rect 2929 4322 2982 4327
rect 3369 4322 3854 4327
rect 3953 4322 3958 4332
rect 2233 4317 2326 4322
rect 3001 4317 3206 4322
rect 2033 4312 2238 4317
rect 2321 4312 2766 4317
rect 2905 4312 3006 4317
rect 3201 4312 4158 4317
rect 2161 4302 2438 4307
rect 2777 4302 2870 4307
rect 2881 4302 3190 4307
rect 3305 4302 3334 4307
rect 3361 4302 3734 4307
rect 2625 4297 2782 4302
rect 2881 4297 2886 4302
rect 3185 4297 3310 4302
rect 2153 4292 2246 4297
rect 2273 4292 2310 4297
rect 2329 4292 2478 4297
rect 2497 4292 2630 4297
rect 2817 4292 2886 4297
rect 3025 4292 3166 4297
rect 2305 4287 2310 4292
rect 2497 4287 2502 4292
rect 2905 4287 3006 4292
rect 3361 4287 3366 4302
rect 3833 4297 3942 4302
rect 3393 4292 3638 4297
rect 3809 4292 3838 4297
rect 3937 4292 3966 4297
rect 529 4282 638 4287
rect 1769 4282 1838 4287
rect 1857 4282 1958 4287
rect 1977 4282 2102 4287
rect 2121 4282 2294 4287
rect 2305 4282 2502 4287
rect 2641 4282 2694 4287
rect 2705 4282 2750 4287
rect 2761 4282 2910 4287
rect 3001 4282 3078 4287
rect 1769 4277 1774 4282
rect 1529 4272 1774 4277
rect 1833 4277 1838 4282
rect 1977 4277 1982 4282
rect 1833 4272 1910 4277
rect 1921 4272 1982 4277
rect 2097 4277 2102 4282
rect 2641 4277 2646 4282
rect 3073 4277 3078 4282
rect 3169 4282 3366 4287
rect 3457 4282 3486 4287
rect 3649 4282 3678 4287
rect 3833 4282 3910 4287
rect 3921 4282 4006 4287
rect 3169 4277 3174 4282
rect 3481 4277 3654 4282
rect 3905 4277 3910 4282
rect 2097 4272 2182 4277
rect 2193 4272 2286 4277
rect 2297 4272 2526 4277
rect 2585 4272 2646 4277
rect 2657 4272 2822 4277
rect 2833 4272 2878 4277
rect 2889 4272 3054 4277
rect 3073 4272 3174 4277
rect 3697 4272 3758 4277
rect 3905 4272 4014 4277
rect 3777 4267 3886 4272
rect 377 4262 510 4267
rect 1793 4262 1854 4267
rect 1937 4262 2910 4267
rect 2945 4262 2998 4267
rect 3353 4262 3422 4267
rect 3441 4262 3526 4267
rect 3545 4262 3678 4267
rect 3729 4262 3782 4267
rect 3881 4262 3926 4267
rect 129 4252 222 4257
rect 129 4247 134 4252
rect 105 4242 134 4247
rect 217 4247 222 4252
rect 377 4247 382 4262
rect 217 4242 382 4247
rect 505 4247 510 4262
rect 3353 4257 3358 4262
rect 553 4252 606 4257
rect 1785 4252 2838 4257
rect 2849 4252 2998 4257
rect 3057 4252 3150 4257
rect 3169 4252 3310 4257
rect 3329 4252 3358 4257
rect 3417 4257 3422 4262
rect 3545 4257 3550 4262
rect 3417 4252 3550 4257
rect 3673 4257 3678 4262
rect 3673 4252 3862 4257
rect 3953 4252 4126 4257
rect 3169 4247 3174 4252
rect 505 4242 710 4247
rect 745 4242 806 4247
rect 1569 4242 1598 4247
rect 1801 4242 1942 4247
rect 1985 4242 2086 4247
rect 2105 4242 3174 4247
rect 3305 4247 3310 4252
rect 3305 4242 4022 4247
rect 2081 4237 2086 4242
rect 393 4232 726 4237
rect 1689 4232 2070 4237
rect 2081 4232 2934 4237
rect 3465 4232 4078 4237
rect 2961 4227 3190 4232
rect 3249 4227 3446 4232
rect 121 4222 206 4227
rect 465 4222 590 4227
rect 609 4222 686 4227
rect 1441 4222 1494 4227
rect 1721 4222 2822 4227
rect 2945 4222 2966 4227
rect 3185 4222 3254 4227
rect 3441 4222 3974 4227
rect 3993 4222 4030 4227
rect 2817 4217 2950 4222
rect 569 4212 614 4217
rect 825 4212 958 4217
rect 977 4212 1406 4217
rect 1529 4212 1782 4217
rect 1825 4212 2534 4217
rect 2545 4212 2670 4217
rect 2721 4212 2798 4217
rect 2977 4212 3014 4217
rect 3033 4212 3174 4217
rect 3265 4212 3366 4217
rect 3425 4212 3510 4217
rect 3537 4212 3614 4217
rect 3873 4212 4030 4217
rect 4065 4212 4134 4217
rect 4353 4212 4448 4217
rect 609 4207 614 4212
rect 977 4207 982 4212
rect 3633 4207 3862 4212
rect 513 4202 598 4207
rect 609 4202 718 4207
rect 881 4202 982 4207
rect 1065 4202 1142 4207
rect 1521 4202 1598 4207
rect 2081 4202 2166 4207
rect 2321 4202 2526 4207
rect 2537 4202 2606 4207
rect 2649 4202 2822 4207
rect 2865 4202 3414 4207
rect 3497 4202 3638 4207
rect 3857 4202 3910 4207
rect 4265 4202 4310 4207
rect 881 4197 886 4202
rect 1833 4197 2062 4202
rect 73 4192 142 4197
rect 241 4192 358 4197
rect 577 4192 622 4197
rect 729 4192 886 4197
rect 905 4192 1118 4197
rect 1553 4192 1654 4197
rect 1673 4192 1750 4197
rect 1809 4192 1838 4197
rect 2057 4192 2142 4197
rect 2161 4192 2166 4202
rect 2217 4197 2326 4202
rect 3409 4197 3502 4202
rect 3905 4197 3990 4202
rect 2193 4192 2222 4197
rect 2345 4192 2430 4197
rect 2441 4192 2558 4197
rect 2601 4192 2854 4197
rect 2945 4192 2998 4197
rect 3041 4192 3086 4197
rect 3097 4192 3390 4197
rect 3521 4192 3886 4197
rect 3985 4187 3990 4197
rect 4177 4192 4286 4197
rect 873 4182 926 4187
rect 1465 4182 1534 4187
rect 1737 4182 1814 4187
rect 1825 4182 1870 4187
rect 1897 4182 2014 4187
rect 2025 4182 2646 4187
rect 2657 4182 2758 4187
rect 2769 4182 2910 4187
rect 3025 4182 3118 4187
rect 3185 4182 3222 4187
rect 3241 4182 3318 4187
rect 3377 4182 3486 4187
rect 3497 4182 3566 4187
rect 3745 4182 3822 4187
rect 3865 4182 3950 4187
rect 3985 4182 4126 4187
rect 1465 4177 1470 4182
rect 1409 4172 1470 4177
rect 1529 4177 1534 4182
rect 3585 4177 3726 4182
rect 1529 4172 1990 4177
rect 2065 4172 3590 4177
rect 3721 4172 3998 4177
rect 4113 4172 4142 4177
rect 361 4162 462 4167
rect 633 4162 782 4167
rect 945 4162 1062 4167
rect 1481 4162 1542 4167
rect 1889 4162 2022 4167
rect 2161 4162 2278 4167
rect 2321 4162 3518 4167
rect 3569 4162 3598 4167
rect 3625 4162 3894 4167
rect 361 4157 366 4162
rect 193 4152 262 4157
rect 337 4152 366 4157
rect 457 4157 462 4162
rect 945 4157 950 4162
rect 457 4152 486 4157
rect 761 4152 870 4157
rect 881 4152 950 4157
rect 1057 4157 1062 4162
rect 1601 4157 1766 4162
rect 2041 4157 2142 4162
rect 3993 4157 4150 4162
rect 1057 4152 1350 4157
rect 1577 4152 1606 4157
rect 1761 4152 1790 4157
rect 1841 4152 2046 4157
rect 2137 4152 3998 4157
rect 4145 4152 4342 4157
rect 233 4142 390 4147
rect 385 4137 390 4142
rect 473 4142 830 4147
rect 473 4137 478 4142
rect 865 4137 870 4152
rect 1841 4147 1846 4152
rect 889 4142 966 4147
rect 1001 4142 1134 4147
rect 1417 4142 1470 4147
rect 1505 4142 1606 4147
rect 1617 4142 1846 4147
rect 1865 4142 1910 4147
rect 1945 4142 1966 4147
rect 2017 4142 2158 4147
rect 2169 4142 2190 4147
rect 2201 4142 2230 4147
rect 2249 4142 2270 4147
rect 2289 4142 2326 4147
rect 2361 4142 2510 4147
rect 2665 4142 2686 4147
rect 2777 4142 2894 4147
rect 2913 4142 3254 4147
rect 3361 4142 3390 4147
rect 3473 4142 3518 4147
rect 3553 4142 3910 4147
rect 4009 4142 4030 4147
rect 4041 4142 4134 4147
rect 1601 4137 1606 4142
rect 2529 4137 2646 4142
rect 2913 4137 2918 4142
rect 0 4132 166 4137
rect 385 4132 478 4137
rect 649 4132 670 4137
rect 865 4132 1110 4137
rect 1153 4132 1350 4137
rect 1401 4132 1478 4137
rect 1489 4132 1534 4137
rect 1601 4132 1830 4137
rect 1841 4132 1886 4137
rect 1993 4132 2310 4137
rect 2321 4132 2534 4137
rect 2641 4132 2694 4137
rect 2785 4132 2918 4137
rect 3017 4132 3062 4137
rect 1153 4127 1158 4132
rect 81 4117 86 4127
rect 145 4122 198 4127
rect 673 4122 742 4127
rect 929 4122 1014 4127
rect 1025 4122 1158 4127
rect 1345 4127 1350 4132
rect 1489 4127 1494 4132
rect 1825 4127 1830 4132
rect 2321 4127 2326 4132
rect 2785 4127 2790 4132
rect 3249 4127 3254 4142
rect 3345 4132 3950 4137
rect 3969 4132 4054 4137
rect 4129 4132 4134 4142
rect 4161 4132 4206 4137
rect 4049 4127 4054 4132
rect 1345 4122 1374 4127
rect 1473 4122 1494 4127
rect 1513 4122 1598 4127
rect 1705 4122 1734 4127
rect 1825 4122 2150 4127
rect 2161 4122 2222 4127
rect 2265 4122 2326 4127
rect 2377 4122 2790 4127
rect 2809 4122 2862 4127
rect 2929 4122 3086 4127
rect 3249 4122 3374 4127
rect 3393 4122 3534 4127
rect 3601 4122 3750 4127
rect 3761 4122 3806 4127
rect 3841 4122 3958 4127
rect 3993 4122 4038 4127
rect 4049 4122 4142 4127
rect 4217 4122 4334 4127
rect 0 4112 134 4117
rect 193 4107 198 4122
rect 1233 4117 1326 4122
rect 1593 4117 1710 4122
rect 2857 4117 2934 4122
rect 3745 4117 3750 4122
rect 641 4112 710 4117
rect 841 4112 910 4117
rect 1057 4112 1238 4117
rect 1321 4112 1382 4117
rect 1425 4112 1462 4117
rect 1489 4112 1526 4117
rect 1769 4112 1830 4117
rect 1865 4112 2038 4117
rect 2049 4112 2086 4117
rect 2097 4112 2166 4117
rect 2225 4112 2558 4117
rect 2649 4112 2710 4117
rect 2753 4112 2838 4117
rect 3201 4112 3422 4117
rect 3449 4112 3734 4117
rect 3745 4112 4054 4117
rect 4081 4112 4174 4117
rect 841 4107 846 4112
rect 193 4102 222 4107
rect 545 4102 662 4107
rect 721 4102 846 4107
rect 905 4107 910 4112
rect 1489 4107 1494 4112
rect 2081 4107 2086 4112
rect 905 4102 1006 4107
rect 1121 4102 1494 4107
rect 1537 4102 1878 4107
rect 1953 4102 2022 4107
rect 2081 4102 2158 4107
rect 2169 4102 2198 4107
rect 2281 4102 2646 4107
rect 2657 4102 2782 4107
rect 2953 4102 2998 4107
rect 3017 4102 3094 4107
rect 3217 4102 3358 4107
rect 3465 4102 3494 4107
rect 3505 4102 3566 4107
rect 3585 4102 3646 4107
rect 3697 4102 3742 4107
rect 3753 4102 3774 4107
rect 3785 4102 3990 4107
rect 4001 4102 4022 4107
rect 4041 4102 4102 4107
rect 4137 4102 4246 4107
rect 1873 4097 1878 4102
rect 2641 4097 2646 4102
rect 3017 4097 3022 4102
rect 0 4092 158 4097
rect 625 4092 654 4097
rect 649 4087 654 4092
rect 777 4092 806 4097
rect 865 4092 950 4097
rect 1097 4092 1126 4097
rect 1329 4092 1470 4097
rect 1481 4092 1566 4097
rect 1713 4092 1862 4097
rect 1873 4092 2134 4097
rect 2145 4092 2262 4097
rect 2273 4092 2310 4097
rect 2473 4092 2550 4097
rect 2641 4092 3022 4097
rect 3089 4097 3094 4102
rect 4443 4097 4448 4127
rect 3089 4092 3854 4097
rect 3921 4092 3974 4097
rect 3985 4092 4102 4097
rect 4121 4092 4214 4097
rect 4377 4092 4448 4097
rect 777 4087 782 4092
rect 1121 4087 1334 4092
rect 1561 4087 1718 4092
rect 2329 4087 2454 4092
rect 4097 4087 4102 4092
rect 121 4082 150 4087
rect 649 4082 782 4087
rect 1353 4082 1390 4087
rect 1481 4082 1542 4087
rect 1537 4077 1542 4082
rect 1737 4082 2334 4087
rect 2449 4082 2502 4087
rect 2529 4082 2598 4087
rect 2641 4082 3078 4087
rect 3233 4082 3270 4087
rect 3297 4082 3350 4087
rect 3433 4082 3614 4087
rect 3657 4082 3926 4087
rect 4025 4082 4054 4087
rect 4097 4082 4158 4087
rect 1737 4077 1742 4082
rect 3097 4077 3174 4082
rect 1105 4072 1502 4077
rect 1537 4072 1742 4077
rect 1777 4072 3102 4077
rect 3169 4072 3222 4077
rect 3305 4072 4086 4077
rect 3217 4067 3310 4072
rect 857 4062 1094 4067
rect 1313 4062 1518 4067
rect 1761 4062 2030 4067
rect 2113 4062 2238 4067
rect 2249 4062 2814 4067
rect 2849 4062 3158 4067
rect 3329 4062 3822 4067
rect 1089 4057 1318 4062
rect 3921 4057 4158 4062
rect 0 4052 22 4057
rect 1489 4052 1542 4057
rect 1577 4052 1638 4057
rect 1649 4052 3606 4057
rect 3737 4052 3926 4057
rect 4153 4052 4286 4057
rect 17 4007 22 4052
rect 1337 4047 1470 4052
rect 3601 4047 3742 4052
rect 321 4042 366 4047
rect 569 4042 638 4047
rect 1113 4042 1190 4047
rect 1113 4037 1118 4042
rect 313 4032 454 4037
rect 553 4032 694 4037
rect 945 4032 1118 4037
rect 1185 4037 1190 4042
rect 1313 4042 1342 4047
rect 1465 4042 1694 4047
rect 1849 4042 2110 4047
rect 2121 4042 2174 4047
rect 2273 4042 2294 4047
rect 2329 4042 2358 4047
rect 2385 4042 2486 4047
rect 2561 4042 2622 4047
rect 2713 4042 2830 4047
rect 3001 4042 3070 4047
rect 3081 4042 3166 4047
rect 3457 4042 3582 4047
rect 3761 4042 3814 4047
rect 1313 4037 1318 4042
rect 1713 4037 1830 4042
rect 2849 4037 2982 4042
rect 3185 4037 3398 4042
rect 3825 4037 3830 4047
rect 3937 4042 4142 4047
rect 1185 4032 1318 4037
rect 1353 4032 1718 4037
rect 1825 4032 2494 4037
rect 2537 4032 2854 4037
rect 2977 4032 3190 4037
rect 3393 4032 3550 4037
rect 3633 4032 3718 4037
rect 3753 4032 3790 4037
rect 3825 4032 4006 4037
rect 4097 4032 4198 4037
rect 337 4022 486 4027
rect 513 4022 702 4027
rect 737 4022 814 4027
rect 977 4022 1110 4027
rect 1161 4022 1230 4027
rect 1257 4022 1326 4027
rect 1385 4022 1766 4027
rect 1777 4022 4030 4027
rect 4265 4022 4318 4027
rect 297 4012 374 4017
rect 481 4012 486 4022
rect 737 4017 742 4022
rect 665 4012 742 4017
rect 809 4017 814 4022
rect 809 4012 902 4017
rect 1137 4012 1366 4017
rect 1497 4012 1830 4017
rect 1913 4012 2894 4017
rect 3041 4012 3126 4017
rect 3313 4012 3454 4017
rect 3569 4012 3774 4017
rect 3801 4012 3918 4017
rect 4113 4012 4158 4017
rect 4353 4012 4448 4017
rect 2937 4007 3046 4012
rect 3145 4007 3294 4012
rect 17 4002 230 4007
rect 225 3997 230 4002
rect 513 4002 646 4007
rect 905 4002 982 4007
rect 1345 4002 1390 4007
rect 513 3997 518 4002
rect 641 3997 750 4002
rect 1385 3997 1390 4002
rect 1521 4002 1894 4007
rect 2009 4002 2078 4007
rect 2137 4002 2334 4007
rect 2345 4002 2398 4007
rect 2489 4002 2942 4007
rect 3073 4002 3150 4007
rect 3289 4002 3462 4007
rect 3521 4002 3598 4007
rect 3609 4002 3686 4007
rect 3745 4002 3766 4007
rect 3777 4002 3870 4007
rect 4017 4002 4118 4007
rect 1521 3997 1526 4002
rect 225 3992 254 3997
rect 385 3992 454 3997
rect 489 3992 518 3997
rect 745 3992 774 3997
rect 793 3992 830 3997
rect 1001 3992 1086 3997
rect 1241 3992 1278 3997
rect 1385 3992 1526 3997
rect 1545 3992 1702 3997
rect 1713 3992 1758 3997
rect 1785 3992 1846 3997
rect 1921 3992 1998 3997
rect 2073 3992 2534 3997
rect 2561 3992 2582 3997
rect 2593 3992 2638 3997
rect 2681 3992 2726 3997
rect 2761 3992 2886 3997
rect 2953 3992 3990 3997
rect 1001 3987 1006 3992
rect 337 3982 630 3987
rect 641 3982 1006 3987
rect 1081 3987 1086 3992
rect 1993 3987 2078 3992
rect 1081 3982 1366 3987
rect 1617 3982 1678 3987
rect 1689 3982 1782 3987
rect 1937 3982 1966 3987
rect 2097 3982 2126 3987
rect 2153 3982 2766 3987
rect 2785 3982 2822 3987
rect 625 3977 630 3982
rect 1801 3977 1918 3982
rect 209 3972 430 3977
rect 625 3972 862 3977
rect 1017 3972 1078 3977
rect 1761 3972 1806 3977
rect 1913 3972 2174 3977
rect 2225 3972 2278 3977
rect 2361 3972 2550 3977
rect 2769 3972 2854 3977
rect 489 3967 606 3972
rect 857 3967 1022 3972
rect 2569 3967 2750 3972
rect 2881 3967 2886 3992
rect 4041 3987 4110 3992
rect 2897 3982 2950 3987
rect 3017 3982 3062 3987
rect 3121 3982 3358 3987
rect 3481 3982 3502 3987
rect 3513 3982 3662 3987
rect 3713 3982 3862 3987
rect 4017 3982 4046 3987
rect 4105 3982 4166 3987
rect 4193 3982 4238 3987
rect 2969 3972 3014 3977
rect 3281 3972 3510 3977
rect 3601 3972 3878 3977
rect 3953 3972 4094 3977
rect 225 3962 494 3967
rect 601 3962 838 3967
rect 1785 3962 1822 3967
rect 1841 3962 1910 3967
rect 2065 3962 2574 3967
rect 2745 3962 2838 3967
rect 2881 3962 3038 3967
rect 3137 3962 3598 3967
rect 3681 3962 3718 3967
rect 3793 3962 3894 3967
rect 4009 3962 4046 3967
rect 4057 3962 4086 3967
rect 505 3952 590 3957
rect 625 3952 686 3957
rect 785 3952 1238 3957
rect 1409 3952 1478 3957
rect 1409 3947 1414 3952
rect 81 3942 270 3947
rect 465 3942 846 3947
rect 1385 3942 1414 3947
rect 1473 3947 1478 3952
rect 1601 3952 1686 3957
rect 1705 3952 1830 3957
rect 1889 3952 1910 3957
rect 1929 3952 2062 3957
rect 2073 3952 2110 3957
rect 2185 3952 2358 3957
rect 2497 3952 2670 3957
rect 2705 3952 2790 3957
rect 2841 3952 2878 3957
rect 2889 3952 2958 3957
rect 2993 3952 3054 3957
rect 1601 3947 1606 3952
rect 1473 3942 1518 3947
rect 1577 3942 1606 3947
rect 1681 3947 1686 3952
rect 3137 3947 3142 3962
rect 3161 3952 3198 3957
rect 3369 3952 3406 3957
rect 3425 3952 3494 3957
rect 3505 3952 3542 3957
rect 3585 3952 3726 3957
rect 3761 3952 3910 3957
rect 4049 3952 4182 3957
rect 4193 3952 4238 3957
rect 3217 3947 3350 3952
rect 1681 3942 1782 3947
rect 1953 3942 2166 3947
rect 2209 3942 2374 3947
rect 2393 3942 2486 3947
rect 2521 3942 2614 3947
rect 2625 3942 2694 3947
rect 2729 3942 2750 3947
rect 2769 3942 2806 3947
rect 2833 3942 3142 3947
rect 3153 3942 3222 3947
rect 3345 3942 3814 3947
rect 3993 3942 4070 3947
rect 4201 3942 4222 3947
rect 1777 3937 1958 3942
rect 297 3932 374 3937
rect 537 3932 566 3937
rect 593 3932 622 3937
rect 617 3927 622 3932
rect 825 3932 878 3937
rect 825 3927 830 3932
rect 617 3922 830 3927
rect 873 3927 878 3932
rect 937 3932 966 3937
rect 1433 3932 1654 3937
rect 1713 3932 1758 3937
rect 1977 3932 2158 3937
rect 2385 3932 2430 3937
rect 2497 3932 2534 3937
rect 2561 3932 2662 3937
rect 2753 3932 2782 3937
rect 2793 3932 2862 3937
rect 2937 3932 2982 3937
rect 3009 3932 3054 3937
rect 3089 3932 3110 3937
rect 3177 3932 3230 3937
rect 3281 3932 3342 3937
rect 3473 3932 3622 3937
rect 3673 3932 3710 3937
rect 4009 3932 4078 3937
rect 4105 3932 4448 3937
rect 937 3927 942 3932
rect 2177 3927 2366 3932
rect 3361 3927 3454 3932
rect 3729 3927 3806 3932
rect 873 3922 942 3927
rect 1337 3922 1374 3927
rect 1609 3922 1638 3927
rect 1657 3922 1694 3927
rect 1857 3922 1926 3927
rect 1937 3922 1966 3927
rect 2025 3922 2182 3927
rect 2361 3922 3366 3927
rect 3449 3922 3734 3927
rect 3801 3922 3958 3927
rect 3985 3922 4174 3927
rect 4257 3922 4286 3927
rect 1369 3917 1374 3922
rect 1473 3917 1614 3922
rect 1369 3912 1478 3917
rect 1641 3912 1766 3917
rect 1841 3912 1886 3917
rect 2009 3912 2046 3917
rect 2089 3912 3190 3917
rect 3233 3912 3270 3917
rect 3313 3912 3470 3917
rect 3481 3912 3518 3917
rect 3697 3912 3790 3917
rect 3953 3912 3958 3922
rect 4169 3917 4262 3922
rect 4089 3912 4150 3917
rect 3537 3907 3662 3912
rect 665 3902 782 3907
rect 1497 3902 1718 3907
rect 1785 3902 1942 3907
rect 1993 3902 2022 3907
rect 2073 3902 2150 3907
rect 2169 3902 3542 3907
rect 3657 3902 3886 3907
rect 3929 3902 4374 3907
rect 1017 3892 1214 3897
rect 1633 3892 2166 3897
rect 2209 3892 2310 3897
rect 2329 3892 2406 3897
rect 2425 3892 3238 3897
rect 3257 3892 3446 3897
rect 3497 3892 3646 3897
rect 3729 3892 3846 3897
rect 4073 3892 4198 3897
rect 1017 3877 1022 3892
rect 113 3872 182 3877
rect 201 3872 262 3877
rect 537 3872 670 3877
rect 993 3872 1022 3877
rect 1209 3877 1214 3892
rect 2161 3887 2166 3892
rect 2305 3887 2310 3892
rect 1561 3882 1678 3887
rect 2017 3882 2078 3887
rect 2161 3882 2246 3887
rect 2305 3882 2350 3887
rect 2369 3882 2854 3887
rect 2897 3882 2942 3887
rect 3177 3882 3822 3887
rect 3865 3882 3934 3887
rect 4025 3882 4278 3887
rect 1809 3877 1894 3882
rect 1929 3877 1998 3882
rect 2961 3877 3086 3882
rect 3865 3877 3870 3882
rect 1209 3872 1358 3877
rect 1649 3872 1814 3877
rect 1889 3872 1934 3877
rect 1993 3872 2966 3877
rect 3081 3872 3110 3877
rect 3193 3872 3254 3877
rect 3265 3872 3294 3877
rect 3393 3872 3494 3877
rect 3521 3872 3870 3877
rect 3929 3877 3934 3882
rect 3929 3872 4118 3877
rect 4137 3872 4270 3877
rect 537 3867 542 3872
rect 473 3862 542 3867
rect 665 3867 670 3872
rect 3289 3867 3398 3872
rect 665 3862 1198 3867
rect 1825 3862 1878 3867
rect 1945 3862 2046 3867
rect 2161 3862 2278 3867
rect 2361 3862 2430 3867
rect 2457 3862 2510 3867
rect 2521 3862 2662 3867
rect 2689 3862 2710 3867
rect 2737 3862 3006 3867
rect 3025 3862 3142 3867
rect 3217 3862 3254 3867
rect 3417 3862 3486 3867
rect 3673 3862 3918 3867
rect 4057 3862 4166 3867
rect 4225 3862 4310 3867
rect 3505 3857 3654 3862
rect 4161 3857 4166 3862
rect 281 3852 438 3857
rect 1609 3852 1686 3857
rect 1705 3852 3510 3857
rect 3649 3852 3678 3857
rect 3785 3852 3998 3857
rect 4017 3852 4086 3857
rect 4161 3852 4382 3857
rect 281 3847 286 3852
rect 65 3842 286 3847
rect 433 3847 438 3852
rect 3673 3847 3790 3852
rect 4017 3847 4022 3852
rect 433 3842 462 3847
rect 553 3842 654 3847
rect 1657 3842 1774 3847
rect 1793 3842 1830 3847
rect 1841 3842 2118 3847
rect 2129 3842 2310 3847
rect 2321 3842 2382 3847
rect 2529 3842 2558 3847
rect 2665 3842 2734 3847
rect 2761 3842 3006 3847
rect 3017 3842 3150 3847
rect 3417 3842 3654 3847
rect 3809 3842 3838 3847
rect 1793 3837 1798 3842
rect 465 3832 550 3837
rect 665 3832 1254 3837
rect 1521 3832 1622 3837
rect 1769 3832 1798 3837
rect 1809 3832 1862 3837
rect 2033 3832 2086 3837
rect 545 3827 670 3832
rect 1249 3827 1254 3832
rect 1881 3827 2014 3832
rect 0 3822 526 3827
rect 1249 3822 1286 3827
rect 1425 3822 1550 3827
rect 1689 3822 1718 3827
rect 1737 3822 1886 3827
rect 2009 3822 2054 3827
rect 2113 3817 2118 3842
rect 2321 3837 2326 3842
rect 2401 3837 2510 3842
rect 3169 3837 3270 3842
rect 3833 3837 3838 3842
rect 3953 3842 4022 3847
rect 4065 3842 4102 3847
rect 4113 3842 4448 3847
rect 3953 3837 3958 3842
rect 4113 3837 4118 3842
rect 2169 3832 2230 3837
rect 2257 3832 2326 3837
rect 2337 3832 2406 3837
rect 2505 3832 3174 3837
rect 3265 3832 3462 3837
rect 3489 3832 3558 3837
rect 3681 3832 3790 3837
rect 3833 3832 3958 3837
rect 4017 3832 4118 3837
rect 4145 3832 4206 3837
rect 4225 3827 4334 3832
rect 2137 3822 2270 3827
rect 2281 3822 2318 3827
rect 2353 3822 2726 3827
rect 2809 3822 2870 3827
rect 2881 3822 2998 3827
rect 3065 3822 3134 3827
rect 3169 3822 3230 3827
rect 3369 3822 3526 3827
rect 3601 3822 3758 3827
rect 3993 3822 4102 3827
rect 4121 3822 4230 3827
rect 4329 3822 4358 3827
rect 3249 3817 3374 3822
rect 4353 3817 4358 3822
rect 257 3812 286 3817
rect 497 3812 702 3817
rect 1345 3812 1486 3817
rect 1601 3812 1750 3817
rect 1881 3812 1982 3817
rect 1993 3812 2054 3817
rect 2113 3812 2494 3817
rect 2561 3812 2694 3817
rect 2713 3812 2766 3817
rect 281 3807 286 3812
rect 409 3807 502 3812
rect 1481 3807 1590 3812
rect 1769 3807 1854 3812
rect 2785 3807 2790 3817
rect 2817 3812 3182 3817
rect 3233 3812 3254 3817
rect 3393 3812 3518 3817
rect 3561 3812 3686 3817
rect 3809 3812 3886 3817
rect 4129 3812 4334 3817
rect 4353 3812 4448 3817
rect 3249 3807 3254 3812
rect 3705 3807 3814 3812
rect 3881 3807 3886 3812
rect 97 3802 134 3807
rect 281 3802 414 3807
rect 561 3802 638 3807
rect 1065 3802 1134 3807
rect 1585 3802 1774 3807
rect 1849 3802 2790 3807
rect 2865 3802 2942 3807
rect 3041 3802 3254 3807
rect 3297 3802 3358 3807
rect 3449 3802 3710 3807
rect 3881 3802 3918 3807
rect 3977 3802 4086 3807
rect 4097 3802 4262 3807
rect 1065 3797 1070 3802
rect 201 3792 246 3797
rect 241 3787 246 3792
rect 433 3792 470 3797
rect 601 3792 790 3797
rect 881 3792 1014 3797
rect 1041 3792 1070 3797
rect 1129 3797 1134 3802
rect 2785 3797 2790 3802
rect 4081 3797 4086 3802
rect 4281 3797 4374 3802
rect 1129 3792 1158 3797
rect 1193 3792 1302 3797
rect 1505 3792 1574 3797
rect 1593 3792 1630 3797
rect 1665 3792 1702 3797
rect 1737 3792 1838 3797
rect 1945 3792 1998 3797
rect 2017 3792 2070 3797
rect 2097 3792 2166 3797
rect 2209 3792 2382 3797
rect 2409 3792 2446 3797
rect 2457 3792 2518 3797
rect 2529 3792 2598 3797
rect 2609 3792 2750 3797
rect 2785 3792 3022 3797
rect 3105 3792 3318 3797
rect 3329 3792 3422 3797
rect 3489 3792 3582 3797
rect 3641 3792 3870 3797
rect 3961 3792 4046 3797
rect 4081 3792 4286 3797
rect 4369 3792 4448 3797
rect 433 3787 438 3792
rect 881 3787 886 3792
rect 241 3782 438 3787
rect 457 3782 590 3787
rect 801 3782 886 3787
rect 1009 3787 1014 3792
rect 2593 3787 2598 3792
rect 3313 3787 3318 3792
rect 1009 3782 1030 3787
rect 585 3777 590 3782
rect 665 3777 806 3782
rect 1025 3777 1030 3782
rect 1113 3782 1238 3787
rect 1417 3782 1486 3787
rect 1697 3782 1774 3787
rect 1793 3782 2574 3787
rect 2593 3782 2622 3787
rect 2657 3782 2878 3787
rect 2913 3782 3046 3787
rect 3145 3782 3206 3787
rect 3217 3782 3294 3787
rect 3313 3782 3334 3787
rect 3345 3782 3430 3787
rect 3505 3782 3654 3787
rect 3689 3782 3806 3787
rect 3937 3782 3990 3787
rect 4073 3782 4358 3787
rect 1113 3777 1118 3782
rect 1417 3777 1422 3782
rect 1481 3777 1582 3782
rect 4353 3777 4358 3782
rect 585 3772 670 3777
rect 1025 3772 1118 3777
rect 1225 3772 1366 3777
rect 1393 3772 1422 3777
rect 1577 3772 1606 3777
rect 1657 3772 1734 3777
rect 1753 3772 1814 3777
rect 1825 3772 1886 3777
rect 1985 3772 2022 3777
rect 2049 3772 2534 3777
rect 2609 3772 2654 3777
rect 2665 3772 2838 3777
rect 2849 3772 3070 3777
rect 3193 3772 3358 3777
rect 3513 3772 3598 3777
rect 3609 3772 3686 3777
rect 3985 3772 4022 3777
rect 4033 3772 4110 3777
rect 4209 3772 4302 3777
rect 4353 3772 4448 3777
rect 2833 3767 2838 3772
rect 689 3762 846 3767
rect 689 3757 694 3762
rect 377 3752 694 3757
rect 841 3757 846 3762
rect 897 3762 998 3767
rect 1137 3762 1382 3767
rect 1537 3762 2214 3767
rect 2225 3762 2262 3767
rect 2289 3762 2574 3767
rect 2617 3762 2662 3767
rect 2737 3762 2766 3767
rect 2777 3762 2822 3767
rect 2833 3762 2918 3767
rect 2945 3762 3742 3767
rect 3889 3762 4198 3767
rect 4233 3762 4278 3767
rect 4329 3762 4366 3767
rect 897 3757 902 3762
rect 1377 3757 1542 3762
rect 841 3752 902 3757
rect 913 3752 998 3757
rect 1257 3752 1358 3757
rect 1561 3752 1598 3757
rect 1681 3752 1710 3757
rect 1777 3752 1926 3757
rect 2001 3752 2046 3757
rect 2057 3752 2614 3757
rect 2625 3752 2902 3757
rect 2953 3752 2982 3757
rect 3105 3752 3158 3757
rect 3169 3752 3190 3757
rect 3281 3752 3374 3757
rect 3537 3752 3566 3757
rect 3585 3752 4214 3757
rect 4353 3752 4448 3757
rect 89 3742 406 3747
rect 705 3742 1198 3747
rect 1289 3742 1614 3747
rect 1841 3742 1886 3747
rect 1897 3742 2118 3747
rect 2137 3742 2366 3747
rect 2465 3742 2934 3747
rect 2977 3742 2982 3752
rect 2993 3742 3062 3747
rect 3129 3742 3414 3747
rect 3465 3742 3582 3747
rect 3593 3742 3630 3747
rect 3641 3742 3710 3747
rect 3873 3742 3990 3747
rect 4113 3742 4206 3747
rect 4217 3742 4246 3747
rect 4289 3742 4334 3747
rect 4353 3737 4358 3752
rect 1513 3732 1742 3737
rect 1793 3732 2238 3737
rect 2377 3732 3286 3737
rect 3297 3732 3726 3737
rect 3809 3732 3846 3737
rect 4065 3732 4358 3737
rect 873 3727 942 3732
rect 2233 3727 2382 3732
rect 3297 3727 3302 3732
rect 737 3722 766 3727
rect 761 3717 766 3722
rect 825 3722 878 3727
rect 937 3722 1062 3727
rect 825 3717 830 3722
rect 1057 3717 1062 3722
rect 1137 3722 1166 3727
rect 1353 3722 1558 3727
rect 1625 3722 1758 3727
rect 1809 3722 2142 3727
rect 2177 3722 2214 3727
rect 2417 3722 2478 3727
rect 2497 3722 2614 3727
rect 2633 3722 2758 3727
rect 2777 3722 2798 3727
rect 2833 3722 2854 3727
rect 2865 3722 2902 3727
rect 2937 3722 3302 3727
rect 3329 3722 3494 3727
rect 3513 3722 3534 3727
rect 3545 3722 3590 3727
rect 3681 3722 3758 3727
rect 3873 3722 4270 3727
rect 4369 3722 4448 3727
rect 1137 3717 1142 3722
rect 761 3712 830 3717
rect 897 3712 926 3717
rect 921 3707 926 3712
rect 1009 3712 1038 3717
rect 1057 3712 1142 3717
rect 1209 3712 1286 3717
rect 1361 3712 1430 3717
rect 1009 3707 1014 3712
rect 449 3702 542 3707
rect 921 3702 1014 3707
rect 1553 3707 1558 3722
rect 2753 3717 2758 3722
rect 2849 3717 2854 3722
rect 3489 3717 3494 3722
rect 4289 3717 4374 3722
rect 1577 3712 1726 3717
rect 1785 3712 1838 3717
rect 1865 3712 2470 3717
rect 2489 3712 2710 3717
rect 2753 3712 2830 3717
rect 2849 3712 2870 3717
rect 2881 3712 2942 3717
rect 3225 3712 3310 3717
rect 3409 3712 3438 3717
rect 3489 3712 3542 3717
rect 3553 3712 3646 3717
rect 3833 3712 3934 3717
rect 4049 3712 4086 3717
rect 4097 3712 4294 3717
rect 2705 3707 2710 3712
rect 2881 3707 2886 3712
rect 3033 3707 3126 3712
rect 3553 3707 3558 3712
rect 1553 3702 1582 3707
rect 1649 3702 1910 3707
rect 1969 3702 2030 3707
rect 2065 3702 2118 3707
rect 2241 3702 2582 3707
rect 2593 3702 2686 3707
rect 2705 3702 2886 3707
rect 2897 3702 3038 3707
rect 3121 3702 3254 3707
rect 3268 3702 3342 3707
rect 3353 3702 3558 3707
rect 3577 3702 3838 3707
rect 2577 3697 2582 3702
rect 3268 3697 3273 3702
rect 3833 3697 3838 3702
rect 3921 3702 3998 3707
rect 4041 3702 4166 3707
rect 4177 3702 4448 3707
rect 3921 3697 3926 3702
rect 4177 3697 4182 3702
rect 1697 3692 1990 3697
rect 2033 3692 2078 3697
rect 2185 3692 2270 3697
rect 2353 3692 2414 3697
rect 2441 3692 2542 3697
rect 2577 3692 2766 3697
rect 2801 3692 3238 3697
rect 3257 3692 3273 3697
rect 3281 3692 3630 3697
rect 3785 3692 3814 3697
rect 3833 3692 3926 3697
rect 3969 3692 4182 3697
rect 4225 3692 4246 3697
rect 2801 3687 2806 3692
rect 3625 3687 3790 3692
rect 1345 3682 1502 3687
rect 1521 3682 1590 3687
rect 1521 3677 1526 3682
rect 1441 3672 1526 3677
rect 1585 3677 1590 3682
rect 1697 3682 1822 3687
rect 1889 3682 1926 3687
rect 2041 3682 2062 3687
rect 2113 3682 2806 3687
rect 2817 3682 3606 3687
rect 3945 3682 4126 3687
rect 4185 3682 4448 3687
rect 1697 3677 1702 3682
rect 1585 3672 1702 3677
rect 1777 3672 2654 3677
rect 2729 3672 3526 3677
rect 3553 3672 3662 3677
rect 3697 3672 3750 3677
rect 4033 3672 4374 3677
rect 1305 3667 1406 3672
rect 4369 3667 4374 3672
rect 1281 3662 1310 3667
rect 1401 3662 1678 3667
rect 1713 3662 2086 3667
rect 2105 3662 2358 3667
rect 2409 3662 2462 3667
rect 2497 3662 2630 3667
rect 2665 3662 2694 3667
rect 2705 3662 2734 3667
rect 2793 3662 2902 3667
rect 2913 3662 2990 3667
rect 3065 3662 3670 3667
rect 3937 3662 3966 3667
rect 4169 3662 4254 3667
rect 4305 3657 4310 3667
rect 4369 3662 4448 3667
rect 1297 3652 1526 3657
rect 1601 3652 1766 3657
rect 1857 3652 2094 3657
rect 2233 3652 2262 3657
rect 2273 3652 2478 3657
rect 2489 3652 2638 3657
rect 2689 3652 3622 3657
rect 3657 3652 3774 3657
rect 3865 3652 4310 3657
rect 1761 3647 1862 3652
rect 2145 3647 2214 3652
rect 209 3642 246 3647
rect 241 3637 246 3642
rect 1201 3642 1246 3647
rect 1273 3642 1622 3647
rect 1713 3642 1742 3647
rect 1881 3642 2150 3647
rect 2209 3642 3190 3647
rect 3233 3642 3270 3647
rect 3289 3642 3326 3647
rect 3337 3642 3390 3647
rect 3409 3642 3702 3647
rect 4105 3642 4182 3647
rect 4377 3642 4448 3647
rect 0 3632 166 3637
rect 241 3632 278 3637
rect 961 3632 1022 3637
rect 161 3627 166 3632
rect 1201 3627 1206 3642
rect 1337 3632 1446 3637
rect 1561 3632 1638 3637
rect 1657 3632 1734 3637
rect 1753 3632 2078 3637
rect 2161 3632 2422 3637
rect 2497 3632 2590 3637
rect 2721 3632 2838 3637
rect 2857 3632 2918 3637
rect 2929 3632 2950 3637
rect 2977 3632 3118 3637
rect 3129 3632 3166 3637
rect 2073 3627 2166 3632
rect 3185 3627 3190 3642
rect 3409 3637 3414 3642
rect 3201 3632 3414 3637
rect 3505 3632 3534 3637
rect 3569 3632 3686 3637
rect 3201 3627 3206 3632
rect 3697 3627 3702 3642
rect 3753 3632 3830 3637
rect 3881 3632 3998 3637
rect 4161 3632 4230 3637
rect 4257 3632 4342 3637
rect 4337 3627 4342 3632
rect 161 3622 278 3627
rect 289 3622 358 3627
rect 417 3622 662 3627
rect 833 3622 1078 3627
rect 1121 3622 1206 3627
rect 1217 3622 1422 3627
rect 1481 3622 1598 3627
rect 273 3617 278 3622
rect 417 3617 422 3622
rect 273 3612 422 3617
rect 985 3612 1062 3617
rect 1393 3612 1694 3617
rect 1713 3607 1718 3627
rect 1745 3622 1806 3627
rect 1937 3622 2054 3627
rect 2185 3622 2214 3627
rect 2281 3622 2310 3627
rect 2337 3622 2358 3627
rect 2385 3622 2694 3627
rect 2705 3622 2750 3627
rect 2769 3622 2790 3627
rect 2801 3622 2886 3627
rect 2905 3622 3174 3627
rect 3185 3622 3206 3627
rect 3249 3622 3358 3627
rect 3489 3622 3662 3627
rect 3697 3622 3806 3627
rect 3905 3622 4038 3627
rect 4057 3622 4142 3627
rect 4201 3622 4230 3627
rect 4241 3622 4318 3627
rect 4337 3622 4448 3627
rect 2385 3617 2390 3622
rect 2881 3617 2886 3622
rect 3169 3617 3174 3622
rect 1849 3612 2118 3617
rect 2177 3612 2390 3617
rect 2409 3612 2502 3617
rect 2577 3612 2870 3617
rect 2881 3612 2902 3617
rect 2993 3612 3094 3617
rect 3113 3612 3142 3617
rect 3169 3612 3190 3617
rect 3201 3612 3226 3617
rect 2865 3607 2870 3612
rect 2897 3607 2902 3612
rect 3249 3607 3254 3622
rect 3409 3617 3494 3622
rect 3289 3612 3414 3617
rect 3505 3612 3598 3617
rect 3793 3612 3886 3617
rect 3905 3612 4006 3617
rect 4033 3607 4038 3622
rect 193 3602 270 3607
rect 441 3602 582 3607
rect 809 3602 878 3607
rect 945 3602 1014 3607
rect 1401 3602 1510 3607
rect 1521 3602 1718 3607
rect 1737 3602 1830 3607
rect 1841 3602 2038 3607
rect 2145 3602 2238 3607
rect 2345 3602 2782 3607
rect 2865 3602 2886 3607
rect 2897 3602 3014 3607
rect 3105 3602 3254 3607
rect 3265 3602 3318 3607
rect 3353 3602 3550 3607
rect 3609 3602 3758 3607
rect 4033 3602 4070 3607
rect 4361 3602 4448 3607
rect 289 3597 446 3602
rect 577 3597 582 3602
rect 3105 3597 3110 3602
rect 3545 3597 3614 3602
rect 0 3592 294 3597
rect 577 3592 606 3597
rect 937 3592 966 3597
rect 1025 3592 1158 3597
rect 1225 3592 1374 3597
rect 1409 3592 1470 3597
rect 1625 3592 1782 3597
rect 1801 3592 1830 3597
rect 1873 3592 3110 3597
rect 3129 3592 3494 3597
rect 3713 3592 3750 3597
rect 3953 3592 4046 3597
rect 4265 3592 4374 3597
rect 177 3582 182 3592
rect 961 3587 1030 3592
rect 1225 3587 1230 3592
rect 233 3582 318 3587
rect 345 3582 430 3587
rect 449 3582 702 3587
rect 1089 3582 1150 3587
rect 1201 3582 1230 3587
rect 1369 3587 1374 3592
rect 1489 3587 1582 3592
rect 1369 3582 1406 3587
rect 1417 3582 1494 3587
rect 1577 3582 1638 3587
rect 1657 3582 1718 3587
rect 1729 3582 2390 3587
rect 2401 3582 2910 3587
rect 2921 3582 3054 3587
rect 3113 3582 3174 3587
rect 3185 3582 3268 3587
rect 3273 3582 3582 3587
rect 3593 3582 3870 3587
rect 3913 3582 3982 3587
rect 4041 3582 4078 3587
rect 4417 3582 4448 3587
rect 2385 3577 2390 3582
rect 3263 3577 3268 3582
rect 1025 3572 1358 3577
rect 1369 3572 1686 3577
rect 1777 3572 1838 3577
rect 1857 3572 1902 3577
rect 1913 3572 1950 3577
rect 1961 3572 2022 3577
rect 2033 3572 2086 3577
rect 2121 3572 2158 3577
rect 2225 3572 2278 3577
rect 2385 3572 2974 3577
rect 2993 3572 3078 3577
rect 3161 3572 3198 3577
rect 3209 3572 3254 3577
rect 3263 3572 3294 3577
rect 3305 3572 3334 3577
rect 3353 3572 3446 3577
rect 3457 3572 3630 3577
rect 3721 3572 3790 3577
rect 3929 3572 4286 3577
rect 201 3567 302 3572
rect 1777 3567 1782 3572
rect 3441 3567 3446 3572
rect 0 3562 206 3567
rect 297 3562 486 3567
rect 817 3562 902 3567
rect 1153 3562 1614 3567
rect 1689 3562 1782 3567
rect 1865 3562 1910 3567
rect 2001 3562 2054 3567
rect 2097 3562 2382 3567
rect 2481 3562 2582 3567
rect 2593 3562 2638 3567
rect 2665 3562 2718 3567
rect 2745 3562 2774 3567
rect 2825 3562 3286 3567
rect 3297 3562 3414 3567
rect 3441 3562 3574 3567
rect 3657 3562 3718 3567
rect 3737 3562 3862 3567
rect 3913 3562 3966 3567
rect 4105 3562 4246 3567
rect 817 3557 822 3562
rect 2577 3557 2582 3562
rect 4417 3557 4422 3582
rect 217 3552 414 3557
rect 409 3547 414 3552
rect 473 3552 502 3557
rect 689 3552 822 3557
rect 841 3552 1070 3557
rect 1137 3552 1166 3557
rect 1273 3552 1558 3557
rect 1569 3552 2070 3557
rect 2081 3552 2222 3557
rect 2233 3552 2278 3557
rect 2321 3552 2566 3557
rect 2577 3552 2630 3557
rect 2641 3552 2830 3557
rect 2841 3552 2942 3557
rect 2953 3552 3446 3557
rect 3481 3552 3526 3557
rect 3753 3552 3878 3557
rect 3897 3552 4206 3557
rect 4305 3552 4422 3557
rect 473 3547 478 3552
rect 2977 3547 2982 3552
rect 4305 3547 4310 3552
rect 265 3542 374 3547
rect 409 3542 478 3547
rect 713 3542 934 3547
rect 1097 3542 1262 3547
rect 1329 3542 2118 3547
rect 2129 3542 2166 3547
rect 2281 3542 2318 3547
rect 2425 3542 2494 3547
rect 2505 3542 2534 3547
rect 2545 3542 2982 3547
rect 3001 3542 3030 3547
rect 3145 3542 3214 3547
rect 3233 3542 3262 3547
rect 3273 3542 3334 3547
rect 3361 3542 3550 3547
rect 3625 3542 3670 3547
rect 3729 3542 3774 3547
rect 3849 3542 3966 3547
rect 4057 3542 4102 3547
rect 4113 3542 4310 3547
rect 369 3527 374 3542
rect 1257 3537 1334 3542
rect 2129 3537 2134 3542
rect 3025 3537 3126 3542
rect 3233 3537 3238 3542
rect 3665 3537 3670 3542
rect 737 3532 830 3537
rect 857 3532 950 3537
rect 969 3532 1078 3537
rect 1113 3532 1142 3537
rect 969 3527 974 3532
rect 161 3522 286 3527
rect 369 3522 390 3527
rect 529 3522 974 3527
rect 1073 3527 1078 3532
rect 1193 3527 1198 3537
rect 1353 3532 1382 3537
rect 1417 3532 1462 3537
rect 1473 3532 1646 3537
rect 1665 3532 2134 3537
rect 2193 3532 2230 3537
rect 2241 3532 2374 3537
rect 2401 3532 2422 3537
rect 2433 3532 2886 3537
rect 3121 3532 3238 3537
rect 3273 3532 3350 3537
rect 3441 3532 3566 3537
rect 3665 3532 3710 3537
rect 1473 3527 1478 3532
rect 1665 3527 1670 3532
rect 1073 3522 1150 3527
rect 1177 3522 1222 3527
rect 1257 3522 1478 3527
rect 1489 3522 1670 3527
rect 1713 3522 1830 3527
rect 1841 3522 2174 3527
rect 2225 3522 2230 3532
rect 2417 3527 2422 3532
rect 2881 3527 2886 3532
rect 3825 3527 3830 3537
rect 4361 3532 4382 3537
rect 2273 3522 2398 3527
rect 2417 3522 2534 3527
rect 2697 3522 2862 3527
rect 2881 3522 2926 3527
rect 2969 3522 3046 3527
rect 3105 3522 3190 3527
rect 3201 3522 3230 3527
rect 3241 3522 3270 3527
rect 3281 3522 3326 3527
rect 3337 3522 3558 3527
rect 3569 3522 3702 3527
rect 3769 3522 3886 3527
rect 3945 3522 4046 3527
rect 4193 3522 4350 3527
rect 4417 3522 4448 3527
rect 1217 3517 1222 3522
rect 1825 3517 1830 3522
rect 2553 3517 2678 3522
rect 4345 3517 4422 3522
rect 673 3512 702 3517
rect 697 3507 702 3512
rect 793 3512 1102 3517
rect 1113 3512 1198 3517
rect 1217 3512 1278 3517
rect 1321 3512 1430 3517
rect 1473 3512 1494 3517
rect 1505 3512 1558 3517
rect 1673 3512 1750 3517
rect 793 3507 798 3512
rect 1761 3507 1766 3517
rect 1825 3512 1846 3517
rect 1905 3512 1926 3517
rect 1945 3512 1974 3517
rect 1993 3512 2150 3517
rect 2177 3512 2294 3517
rect 2313 3512 2558 3517
rect 2673 3512 3430 3517
rect 3473 3512 3654 3517
rect 3777 3512 3854 3517
rect 3889 3512 4022 3517
rect 4081 3512 4190 3517
rect 1921 3507 1926 3512
rect 4017 3507 4022 3512
rect 0 3502 342 3507
rect 353 3502 414 3507
rect 697 3502 798 3507
rect 841 3502 950 3507
rect 1041 3502 1222 3507
rect 1377 3502 1502 3507
rect 1569 3502 1734 3507
rect 1745 3502 1766 3507
rect 1809 3502 1886 3507
rect 1921 3502 1958 3507
rect 1969 3502 2510 3507
rect 2521 3502 2566 3507
rect 2577 3502 2638 3507
rect 2649 3502 2774 3507
rect 2801 3502 2854 3507
rect 2905 3502 3206 3507
rect 3217 3502 3310 3507
rect 3345 3502 3446 3507
rect 3513 3502 3622 3507
rect 3649 3502 3806 3507
rect 3881 3502 3926 3507
rect 4017 3502 4078 3507
rect 1497 3497 1574 3502
rect 1953 3497 1958 3502
rect 2769 3497 2774 3502
rect 2849 3497 2854 3502
rect 3201 3497 3206 3502
rect 401 3492 486 3497
rect 1065 3492 1126 3497
rect 1393 3492 1438 3497
rect 1457 3492 1478 3497
rect 1689 3492 1710 3497
rect 1721 3492 1878 3497
rect 1889 3492 1942 3497
rect 1953 3492 1982 3497
rect 2041 3492 2342 3497
rect 2369 3492 2454 3497
rect 2465 3492 2638 3497
rect 2689 3492 2710 3497
rect 2769 3492 2838 3497
rect 2849 3492 2990 3497
rect 3089 3492 3126 3497
rect 3201 3492 3414 3497
rect 3425 3492 3518 3497
rect 3537 3492 3590 3497
rect 3641 3492 3670 3497
rect 1457 3487 1462 3492
rect 2985 3487 3094 3492
rect 3665 3487 3670 3492
rect 3737 3492 3766 3497
rect 3921 3492 4022 3497
rect 4209 3492 4448 3497
rect 3737 3487 3742 3492
rect 817 3482 846 3487
rect 841 3477 846 3482
rect 905 3482 990 3487
rect 1089 3482 1222 3487
rect 1241 3482 1358 3487
rect 1401 3482 1462 3487
rect 1481 3482 1590 3487
rect 1633 3482 1822 3487
rect 1881 3482 2006 3487
rect 2081 3482 2126 3487
rect 2153 3482 2462 3487
rect 2481 3482 2534 3487
rect 2593 3482 2758 3487
rect 2913 3482 2966 3487
rect 3113 3482 3150 3487
rect 3169 3482 3582 3487
rect 3665 3482 3742 3487
rect 4289 3482 4334 3487
rect 905 3477 910 3482
rect 1241 3477 1246 3482
rect 841 3472 910 3477
rect 929 3472 1078 3477
rect 1161 3472 1246 3477
rect 1353 3477 1358 3482
rect 2081 3477 2086 3482
rect 2793 3477 2894 3482
rect 3169 3477 3174 3482
rect 1353 3472 2086 3477
rect 2145 3472 2182 3477
rect 2193 3472 2230 3477
rect 2281 3472 2318 3477
rect 2361 3472 2422 3477
rect 2449 3472 2550 3477
rect 2569 3472 2614 3477
rect 2641 3472 2798 3477
rect 2889 3472 3174 3477
rect 3193 3472 3238 3477
rect 3249 3472 3334 3477
rect 3345 3472 3582 3477
rect 4001 3472 4022 3477
rect 1073 3467 1166 3472
rect 129 3462 190 3467
rect 361 3462 630 3467
rect 1185 3462 1214 3467
rect 1361 3462 1518 3467
rect 1537 3462 1582 3467
rect 1665 3462 1878 3467
rect 1977 3462 2110 3467
rect 2169 3462 2582 3467
rect 2625 3462 2670 3467
rect 2713 3462 2742 3467
rect 2809 3462 2902 3467
rect 2921 3462 3374 3467
rect 3409 3462 3454 3467
rect 3481 3462 3510 3467
rect 3553 3462 3590 3467
rect 3609 3462 3742 3467
rect 361 3447 366 3462
rect 625 3447 630 3462
rect 1233 3457 1342 3462
rect 3609 3457 3614 3462
rect 1001 3452 1070 3457
rect 1145 3452 1238 3457
rect 1337 3452 2062 3457
rect 2081 3452 2134 3457
rect 2313 3452 2366 3457
rect 2377 3452 2606 3457
rect 2625 3452 3614 3457
rect 3737 3457 3742 3462
rect 3737 3452 3870 3457
rect 4049 3452 4094 3457
rect 4145 3452 4310 3457
rect 2153 3447 2294 3452
rect 337 3442 366 3447
rect 433 3442 542 3447
rect 625 3442 654 3447
rect 825 3442 934 3447
rect 953 3442 1054 3447
rect 1073 3442 1134 3447
rect 1241 3442 1390 3447
rect 1417 3442 1566 3447
rect 1641 3442 2158 3447
rect 2289 3442 3350 3447
rect 3457 3442 3550 3447
rect 3569 3442 3726 3447
rect 3769 3442 3806 3447
rect 3897 3442 3942 3447
rect 433 3437 438 3442
rect 209 3432 278 3437
rect 289 3432 318 3437
rect 377 3432 438 3437
rect 537 3437 542 3442
rect 825 3437 830 3442
rect 537 3432 830 3437
rect 929 3437 934 3442
rect 929 3432 2134 3437
rect 2177 3432 2302 3437
rect 2329 3432 2806 3437
rect 2817 3432 2838 3437
rect 2905 3432 2958 3437
rect 3001 3432 3822 3437
rect 209 3427 214 3432
rect 313 3427 382 3432
rect 113 3422 238 3427
rect 449 3422 526 3427
rect 841 3422 1102 3427
rect 1225 3422 1478 3427
rect 1537 3422 1590 3427
rect 1665 3422 1710 3427
rect 1737 3422 1814 3427
rect 1897 3422 1974 3427
rect 2017 3422 2046 3427
rect 2081 3422 2238 3427
rect 2353 3422 2454 3427
rect 2481 3422 2502 3427
rect 2529 3422 3430 3427
rect 3449 3422 3478 3427
rect 3489 3422 3614 3427
rect 3697 3422 3846 3427
rect 3977 3422 4078 3427
rect 449 3417 454 3422
rect 3473 3417 3478 3422
rect 0 3412 246 3417
rect 241 3407 246 3412
rect 353 3412 454 3417
rect 745 3412 822 3417
rect 961 3412 1086 3417
rect 1153 3412 1254 3417
rect 1265 3412 1614 3417
rect 1689 3412 1998 3417
rect 2033 3412 2990 3417
rect 3057 3412 3102 3417
rect 3137 3412 3222 3417
rect 3241 3412 3286 3417
rect 3297 3412 3342 3417
rect 3377 3412 3422 3417
rect 3433 3412 3462 3417
rect 3473 3412 3574 3417
rect 3617 3412 3702 3417
rect 3857 3412 3886 3417
rect 3969 3412 4134 3417
rect 4257 3412 4358 3417
rect 353 3407 358 3412
rect 745 3407 750 3412
rect 817 3407 902 3412
rect 3457 3407 3462 3412
rect 137 3402 206 3407
rect 241 3402 358 3407
rect 585 3402 750 3407
rect 897 3402 926 3407
rect 1057 3402 1262 3407
rect 1337 3402 1406 3407
rect 1441 3402 1462 3407
rect 1497 3402 1566 3407
rect 1657 3402 1742 3407
rect 1753 3402 1862 3407
rect 1953 3402 2454 3407
rect 2481 3402 2534 3407
rect 2577 3402 2766 3407
rect 2801 3402 2854 3407
rect 2865 3402 3030 3407
rect 3209 3402 3254 3407
rect 3297 3402 3326 3407
rect 3369 3402 3446 3407
rect 3457 3402 3494 3407
rect 3513 3402 3558 3407
rect 3569 3402 3574 3412
rect 3697 3407 3862 3412
rect 3601 3402 3678 3407
rect 4009 3402 4126 3407
rect 4233 3402 4318 3407
rect 377 3392 606 3397
rect 761 3392 862 3397
rect 969 3392 1798 3397
rect 1873 3392 2070 3397
rect 2113 3392 2318 3397
rect 2353 3392 3262 3397
rect 3273 3392 3318 3397
rect 3353 3392 3478 3397
rect 3529 3392 3694 3397
rect 3761 3392 3798 3397
rect 3833 3392 3918 3397
rect 3929 3392 4174 3397
rect 4201 3392 4254 3397
rect 1793 3387 1878 3392
rect 4369 3387 4374 3427
rect 593 3382 870 3387
rect 881 3382 982 3387
rect 1169 3382 1214 3387
rect 1257 3382 1670 3387
rect 1729 3382 1774 3387
rect 1921 3382 2654 3387
rect 2665 3382 3142 3387
rect 3153 3382 3238 3387
rect 3249 3382 3494 3387
rect 3505 3382 3542 3387
rect 3569 3382 3662 3387
rect 3737 3382 3782 3387
rect 3801 3382 3942 3387
rect 4009 3382 4038 3387
rect 4353 3382 4374 3387
rect 1001 3377 1134 3382
rect 3505 3377 3510 3382
rect 4033 3377 4214 3382
rect 4353 3377 4358 3382
rect 73 3372 206 3377
rect 641 3372 670 3377
rect 73 3357 78 3372
rect 0 3352 78 3357
rect 201 3357 206 3372
rect 665 3367 670 3372
rect 809 3372 1006 3377
rect 1129 3372 1158 3377
rect 809 3367 814 3372
rect 1153 3367 1158 3372
rect 1257 3372 1286 3377
rect 1297 3372 1374 3377
rect 1473 3372 1510 3377
rect 1577 3372 1614 3377
rect 1625 3372 1846 3377
rect 1929 3372 2414 3377
rect 2425 3372 2646 3377
rect 2665 3372 2742 3377
rect 2753 3372 3462 3377
rect 3473 3372 3510 3377
rect 3521 3372 3622 3377
rect 3689 3372 3878 3377
rect 4209 3372 4358 3377
rect 1257 3367 1262 3372
rect 241 3362 526 3367
rect 665 3362 814 3367
rect 833 3362 862 3367
rect 945 3362 1110 3367
rect 1153 3362 1262 3367
rect 1313 3362 1382 3367
rect 1521 3362 1670 3367
rect 1809 3362 1830 3367
rect 1897 3362 1958 3367
rect 1977 3362 2006 3367
rect 2041 3362 2110 3367
rect 2137 3362 2262 3367
rect 2289 3362 2342 3367
rect 2353 3362 2398 3367
rect 2425 3362 2582 3367
rect 2593 3362 3206 3367
rect 3233 3362 3438 3367
rect 3449 3362 3502 3367
rect 3513 3362 3566 3367
rect 3609 3362 3774 3367
rect 3873 3362 4190 3367
rect 241 3357 246 3362
rect 857 3357 950 3362
rect 2289 3357 2294 3362
rect 201 3352 246 3357
rect 969 3352 1022 3357
rect 1353 3352 1398 3357
rect 1425 3352 1510 3357
rect 1569 3352 1654 3357
rect 1689 3352 2038 3357
rect 2073 3352 2110 3357
rect 2121 3352 2182 3357
rect 2201 3352 2294 3357
rect 2321 3352 3638 3357
rect 3649 3352 3734 3357
rect 3753 3347 3902 3352
rect 89 3342 150 3347
rect 193 3342 270 3347
rect 721 3342 814 3347
rect 913 3342 1158 3347
rect 1249 3342 1686 3347
rect 1777 3342 1830 3347
rect 1953 3342 2486 3347
rect 2545 3342 2590 3347
rect 2609 3342 2662 3347
rect 2689 3342 2774 3347
rect 2817 3342 2878 3347
rect 2929 3342 3078 3347
rect 3129 3342 3182 3347
rect 3265 3342 3310 3347
rect 3353 3342 3470 3347
rect 3529 3342 3558 3347
rect 3569 3342 3758 3347
rect 3897 3342 3926 3347
rect 4033 3342 4078 3347
rect 4089 3342 4198 3347
rect 4209 3342 4254 3347
rect 4265 3342 4374 3347
rect 721 3337 726 3342
rect 289 3332 382 3337
rect 697 3332 726 3337
rect 809 3337 814 3342
rect 809 3332 990 3337
rect 1113 3332 1238 3337
rect 1337 3332 1718 3337
rect 1745 3332 1894 3337
rect 2017 3332 2462 3337
rect 289 3327 294 3332
rect 113 3322 294 3327
rect 377 3327 382 3332
rect 1233 3327 1342 3332
rect 377 3322 806 3327
rect 977 3322 1062 3327
rect 1361 3322 1542 3327
rect 1561 3322 1622 3327
rect 1633 3322 1894 3327
rect 2009 3322 2142 3327
rect 2153 3322 2310 3327
rect 2353 3322 2462 3327
rect 113 3317 118 3322
rect 1633 3317 1638 3322
rect 2481 3317 2486 3342
rect 2769 3337 2774 3342
rect 2929 3337 2934 3342
rect 2497 3332 2758 3337
rect 2769 3332 2814 3337
rect 2825 3332 2934 3337
rect 2945 3332 3046 3337
rect 3057 3332 3126 3337
rect 3177 3332 3606 3337
rect 3633 3332 3870 3337
rect 4049 3332 4142 3337
rect 2505 3322 2542 3327
rect 2585 3322 3502 3327
rect 3513 3322 3678 3327
rect 3737 3322 3822 3327
rect 3897 3322 4110 3327
rect 4105 3317 4110 3322
rect 4177 3322 4206 3327
rect 4177 3317 4182 3322
rect 0 3312 118 3317
rect 729 3312 758 3317
rect 753 3307 758 3312
rect 897 3312 1030 3317
rect 1249 3312 1310 3317
rect 1377 3312 1542 3317
rect 1601 3312 1638 3317
rect 1665 3312 1782 3317
rect 1865 3312 2470 3317
rect 2481 3312 2846 3317
rect 2865 3312 3006 3317
rect 3049 3312 3142 3317
rect 3185 3312 3326 3317
rect 3409 3312 3558 3317
rect 3593 3312 3670 3317
rect 3801 3312 3894 3317
rect 4049 3312 4086 3317
rect 4105 3312 4182 3317
rect 4233 3312 4318 3317
rect 897 3307 902 3312
rect 145 3302 174 3307
rect 169 3297 174 3302
rect 241 3302 382 3307
rect 241 3297 246 3302
rect 169 3292 246 3297
rect 377 3297 382 3302
rect 585 3302 614 3307
rect 753 3302 902 3307
rect 1217 3302 1334 3307
rect 1369 3302 1406 3307
rect 1417 3302 1486 3307
rect 1537 3302 1542 3312
rect 1593 3302 1702 3307
rect 1737 3302 1830 3307
rect 1857 3302 1910 3307
rect 1929 3302 2102 3307
rect 2113 3302 2366 3307
rect 2377 3302 2654 3307
rect 2713 3302 2742 3307
rect 2753 3302 3494 3307
rect 3513 3302 3542 3307
rect 3585 3302 3630 3307
rect 3705 3302 3814 3307
rect 585 3297 590 3302
rect 377 3292 590 3297
rect 921 3292 1110 3297
rect 1289 3292 1686 3297
rect 1697 3292 1702 3302
rect 1905 3297 1910 3302
rect 2097 3297 2102 3302
rect 1801 3292 1854 3297
rect 1905 3292 2086 3297
rect 2097 3292 2846 3297
rect 2945 3292 2990 3297
rect 3089 3292 3222 3297
rect 3233 3292 3294 3297
rect 3345 3292 3374 3297
rect 3457 3292 3646 3297
rect 3761 3292 3886 3297
rect 1305 3282 1382 3287
rect 1489 3282 1582 3287
rect 1617 3282 1670 3287
rect 1689 3282 1742 3287
rect 1753 3282 2630 3287
rect 2649 3282 2742 3287
rect 2833 3282 3022 3287
rect 3105 3282 3126 3287
rect 3217 3277 3222 3292
rect 3273 3282 3534 3287
rect 993 3272 2934 3277
rect 2945 3272 3102 3277
rect 3129 3272 3158 3277
rect 3217 3272 3350 3277
rect 3361 3272 3606 3277
rect 3633 3272 4030 3277
rect 1265 3262 1350 3267
rect 1537 3262 1598 3267
rect 1633 3262 1766 3267
rect 1777 3262 1862 3267
rect 1953 3262 2086 3267
rect 2137 3262 2286 3267
rect 2361 3262 2958 3267
rect 3113 3262 3190 3267
rect 3281 3262 3334 3267
rect 1953 3257 1958 3262
rect 3185 3257 3190 3262
rect 3345 3257 3350 3272
rect 3385 3262 3422 3267
rect 3441 3262 3606 3267
rect 3753 3257 3822 3262
rect 449 3252 518 3257
rect 1089 3252 1206 3257
rect 1489 3252 1558 3257
rect 1569 3252 1774 3257
rect 1841 3252 1958 3257
rect 1969 3252 2174 3257
rect 2225 3252 2278 3257
rect 2289 3252 2566 3257
rect 2577 3252 2846 3257
rect 2857 3252 2894 3257
rect 3001 3252 3134 3257
rect 3185 3252 3270 3257
rect 3345 3252 3582 3257
rect 3609 3252 3758 3257
rect 3817 3252 3846 3257
rect 449 3247 454 3252
rect 129 3242 454 3247
rect 513 3247 518 3252
rect 1969 3247 1974 3252
rect 2577 3247 2582 3252
rect 513 3242 646 3247
rect 1097 3242 1126 3247
rect 1209 3242 1238 3247
rect 1257 3242 1470 3247
rect 1513 3242 1710 3247
rect 1753 3242 1974 3247
rect 1993 3242 2070 3247
rect 2089 3242 2142 3247
rect 2161 3242 2334 3247
rect 2401 3242 2582 3247
rect 2633 3242 2710 3247
rect 2737 3242 3422 3247
rect 3433 3242 3678 3247
rect 3769 3242 3854 3247
rect 3921 3242 4102 3247
rect 1257 3237 1262 3242
rect 625 3227 630 3237
rect 137 3222 190 3227
rect 465 3222 630 3227
rect 753 3232 846 3237
rect 873 3232 1262 3237
rect 1465 3237 1470 3242
rect 1465 3232 1590 3237
rect 1721 3232 2974 3237
rect 3081 3232 3190 3237
rect 3273 3232 3478 3237
rect 3601 3232 3790 3237
rect 753 3217 758 3232
rect 841 3227 846 3232
rect 1585 3227 1726 3232
rect 3473 3227 3606 3232
rect 841 3222 918 3227
rect 1145 3222 1470 3227
rect 1497 3222 1566 3227
rect 1745 3222 1766 3227
rect 1809 3222 1950 3227
rect 1977 3222 2262 3227
rect 2297 3222 2374 3227
rect 2417 3222 2438 3227
rect 913 3217 918 3222
rect 241 3212 518 3217
rect 665 3212 758 3217
rect 793 3212 878 3217
rect 913 3212 942 3217
rect 1081 3212 1270 3217
rect 1281 3212 1638 3217
rect 1761 3207 1766 3222
rect 2449 3217 2454 3227
rect 2473 3222 2526 3227
rect 2537 3222 2670 3227
rect 2705 3222 2782 3227
rect 2801 3217 2806 3227
rect 2825 3222 3358 3227
rect 3363 3222 3454 3227
rect 3625 3222 3830 3227
rect 3945 3222 3982 3227
rect 4001 3222 4038 3227
rect 4073 3222 4182 3227
rect 4001 3217 4006 3222
rect 1833 3212 1870 3217
rect 2065 3212 2454 3217
rect 2465 3212 3502 3217
rect 3681 3212 3774 3217
rect 3817 3212 3886 3217
rect 3921 3212 4006 3217
rect 1865 3207 2070 3212
rect 169 3202 270 3207
rect 393 3202 526 3207
rect 809 3202 998 3207
rect 1193 3202 1270 3207
rect 1393 3202 1430 3207
rect 1529 3202 1726 3207
rect 1737 3202 1766 3207
rect 1793 3202 1846 3207
rect 2089 3202 2382 3207
rect 2425 3202 2470 3207
rect 2529 3202 2558 3207
rect 2569 3202 2574 3212
rect 2649 3202 2726 3207
rect 2737 3202 2830 3207
rect 1017 3197 1126 3202
rect 1393 3197 1398 3202
rect 1841 3197 1846 3202
rect 2849 3197 2854 3212
rect 3561 3207 3662 3212
rect 2873 3202 3206 3207
rect 3305 3202 3430 3207
rect 3537 3202 3566 3207
rect 3657 3202 3718 3207
rect 3937 3202 4038 3207
rect 4049 3202 4126 3207
rect 4233 3202 4310 3207
rect 3537 3197 3542 3202
rect 4033 3197 4038 3202
rect 281 3192 382 3197
rect 849 3192 878 3197
rect 961 3192 1022 3197
rect 1121 3192 1150 3197
rect 1313 3192 1366 3197
rect 1377 3192 1398 3197
rect 1585 3192 1702 3197
rect 1841 3192 2110 3197
rect 2121 3192 2158 3197
rect 2177 3192 2230 3197
rect 2273 3192 2662 3197
rect 2769 3192 2838 3197
rect 2849 3192 2878 3197
rect 2969 3192 3046 3197
rect 3105 3192 3190 3197
rect 3209 3192 3486 3197
rect 3505 3192 3542 3197
rect 3553 3192 3670 3197
rect 3681 3192 3758 3197
rect 3849 3192 3918 3197
rect 4033 3192 4214 3197
rect 4257 3192 4366 3197
rect 873 3187 966 3192
rect 1585 3187 1590 3192
rect 3505 3187 3510 3192
rect 3681 3187 3686 3192
rect 257 3182 286 3187
rect 281 3177 286 3182
rect 345 3182 470 3187
rect 713 3182 790 3187
rect 985 3182 1134 3187
rect 1353 3182 1518 3187
rect 1537 3182 1590 3187
rect 1609 3182 1846 3187
rect 1865 3182 2510 3187
rect 2537 3182 3414 3187
rect 3449 3182 3510 3187
rect 3649 3182 3686 3187
rect 3737 3182 4022 3187
rect 345 3177 350 3182
rect 713 3177 718 3182
rect 281 3172 350 3177
rect 513 3172 598 3177
rect 617 3172 718 3177
rect 785 3177 790 3182
rect 1841 3177 1846 3182
rect 4017 3177 4022 3182
rect 4161 3182 4190 3187
rect 4201 3182 4254 3187
rect 4161 3177 4166 3182
rect 785 3172 966 3177
rect 1065 3172 1126 3177
rect 1201 3172 1358 3177
rect 1369 3172 1566 3177
rect 1601 3172 1734 3177
rect 1841 3172 1958 3177
rect 2017 3172 2686 3177
rect 2713 3172 2750 3177
rect 2849 3172 2934 3177
rect 2945 3172 3030 3177
rect 3113 3172 3134 3177
rect 3161 3172 3478 3177
rect 3577 3172 3894 3177
rect 4017 3172 4166 3177
rect 513 3167 518 3172
rect 489 3162 518 3167
rect 593 3167 598 3172
rect 593 3162 806 3167
rect 1097 3162 1270 3167
rect 1337 3162 1398 3167
rect 1417 3162 1534 3167
rect 1633 3162 1910 3167
rect 1945 3162 2006 3167
rect 2089 3162 2942 3167
rect 3041 3162 3686 3167
rect 3705 3162 3934 3167
rect 801 3157 806 3162
rect 2937 3157 3046 3162
rect 4121 3157 4190 3162
rect 137 3152 230 3157
rect 481 3152 662 3157
rect 801 3152 878 3157
rect 961 3152 1182 3157
rect 1225 3152 1326 3157
rect 1337 3152 1638 3157
rect 1681 3152 1798 3157
rect 1809 3152 2318 3157
rect 2329 3152 2918 3157
rect 3121 3152 3382 3157
rect 3393 3152 3566 3157
rect 3633 3152 3862 3157
rect 4017 3152 4126 3157
rect 4185 3152 4286 3157
rect 601 3142 830 3147
rect 1161 3142 1670 3147
rect 1721 3142 1862 3147
rect 1937 3142 2022 3147
rect 2033 3142 2902 3147
rect 3025 3142 3174 3147
rect 3201 3142 3254 3147
rect 3289 3142 3334 3147
rect 3369 3142 3622 3147
rect 3705 3142 3734 3147
rect 3801 3142 3846 3147
rect 1857 3137 1862 3142
rect 3617 3137 3710 3142
rect 3841 3137 3846 3142
rect 3945 3142 4006 3147
rect 3945 3137 3950 3142
rect 209 3132 590 3137
rect 585 3117 590 3132
rect 841 3132 1846 3137
rect 1857 3132 1910 3137
rect 1929 3132 2046 3137
rect 2065 3132 2094 3137
rect 2105 3132 2206 3137
rect 2233 3132 2294 3137
rect 2417 3132 2798 3137
rect 2809 3132 3566 3137
rect 3841 3132 3950 3137
rect 4001 3137 4006 3142
rect 4145 3142 4174 3147
rect 4241 3142 4366 3147
rect 4145 3137 4150 3142
rect 4001 3132 4150 3137
rect 4225 3132 4310 3137
rect 841 3117 846 3132
rect 1105 3122 1206 3127
rect 1489 3122 2270 3127
rect 2425 3122 3510 3127
rect 3649 3122 3822 3127
rect 953 3117 1022 3122
rect 1201 3117 1494 3122
rect 2289 3117 2406 3122
rect 145 3112 190 3117
rect 217 3112 254 3117
rect 585 3112 846 3117
rect 897 3112 958 3117
rect 1017 3112 1094 3117
rect 1153 3112 1182 3117
rect 1513 3112 1582 3117
rect 1593 3112 1638 3117
rect 1713 3112 1998 3117
rect 2017 3112 2294 3117
rect 2401 3112 3638 3117
rect 1089 3107 1158 3112
rect 3633 3107 3638 3112
rect 3769 3112 3798 3117
rect 3769 3107 3774 3112
rect 177 3102 310 3107
rect 401 3102 510 3107
rect 969 3102 1006 3107
rect 1265 3102 1534 3107
rect 1561 3102 1606 3107
rect 1705 3102 3126 3107
rect 3137 3102 3454 3107
rect 3497 3102 3614 3107
rect 3633 3102 3774 3107
rect 4081 3102 4254 3107
rect 1105 3092 1246 3097
rect 1625 3092 1942 3097
rect 2009 3092 2374 3097
rect 2433 3092 2814 3097
rect 2841 3092 2886 3097
rect 2897 3092 2934 3097
rect 3009 3092 3078 3097
rect 3145 3092 3398 3097
rect 3409 3092 3470 3097
rect 3481 3092 3598 3097
rect 1105 3087 1110 3092
rect 297 3082 422 3087
rect 1081 3082 1110 3087
rect 1241 3087 1246 3092
rect 1361 3087 1550 3092
rect 2897 3087 2902 3092
rect 3009 3087 3014 3092
rect 1241 3082 1310 3087
rect 1337 3082 1366 3087
rect 1545 3082 1574 3087
rect 1617 3082 1686 3087
rect 1705 3082 1782 3087
rect 1825 3082 1878 3087
rect 1905 3082 1966 3087
rect 1985 3082 2262 3087
rect 2273 3082 2318 3087
rect 2361 3082 2526 3087
rect 2585 3082 2630 3087
rect 2641 3082 2678 3087
rect 2721 3082 2758 3087
rect 2801 3082 2902 3087
rect 2913 3082 3014 3087
rect 3025 3082 3174 3087
rect 3209 3082 3270 3087
rect 3281 3082 3350 3087
rect 3441 3082 3566 3087
rect 1617 3077 1622 3082
rect 1065 3072 1238 3077
rect 1297 3072 1622 3077
rect 1633 3072 1742 3077
rect 1793 3072 1814 3077
rect 1985 3072 1990 3082
rect 2057 3072 2118 3077
rect 2305 3072 3038 3077
rect 3121 3072 3150 3077
rect 3177 3072 3206 3077
rect 3361 3072 3630 3077
rect 3817 3072 3902 3077
rect 1833 3067 1990 3072
rect 2113 3067 2310 3072
rect 3033 3067 3126 3072
rect 3201 3067 3366 3072
rect 1041 3062 1070 3067
rect 1193 3062 1838 3067
rect 2017 3062 2094 3067
rect 2329 3062 2446 3067
rect 2465 3062 2534 3067
rect 2617 3062 2830 3067
rect 2849 3062 2894 3067
rect 2921 3062 3014 3067
rect 3401 3062 3518 3067
rect 1065 3057 1198 3062
rect 505 3052 766 3057
rect 505 3037 510 3052
rect 409 3032 510 3037
rect 761 3037 766 3052
rect 881 3052 1022 3057
rect 1217 3052 1590 3057
rect 1625 3052 2302 3057
rect 2377 3052 3046 3057
rect 3065 3052 3158 3057
rect 3177 3052 3342 3057
rect 3361 3052 3622 3057
rect 881 3037 886 3052
rect 761 3032 790 3037
rect 857 3032 886 3037
rect 1017 3037 1022 3052
rect 3041 3047 3046 3052
rect 3177 3047 3182 3052
rect 1073 3042 1118 3047
rect 1185 3042 1358 3047
rect 1401 3042 1478 3047
rect 1489 3042 1558 3047
rect 1577 3042 1622 3047
rect 1665 3042 2006 3047
rect 2073 3042 2246 3047
rect 2257 3042 2286 3047
rect 2457 3042 2486 3047
rect 2585 3042 2622 3047
rect 2673 3042 2766 3047
rect 2785 3042 2862 3047
rect 2873 3042 2966 3047
rect 3041 3042 3182 3047
rect 3337 3047 3342 3052
rect 3337 3042 3574 3047
rect 2481 3037 2590 3042
rect 3201 3037 3318 3042
rect 1017 3032 1262 3037
rect 1273 3032 1662 3037
rect 1721 3032 1822 3037
rect 1913 3032 1958 3037
rect 2065 3032 2214 3037
rect 2353 3032 2438 3037
rect 2609 3032 2694 3037
rect 2729 3032 3062 3037
rect 3113 3032 3206 3037
rect 3313 3032 3542 3037
rect 3641 3032 3814 3037
rect 3833 3032 3870 3037
rect 2249 3027 2358 3032
rect 3641 3027 3646 3032
rect 161 3022 318 3027
rect 521 3022 622 3027
rect 633 3022 966 3027
rect 1017 3022 1070 3027
rect 1153 3022 2254 3027
rect 2369 3022 2542 3027
rect 2553 3022 2710 3027
rect 2761 3022 2822 3027
rect 961 3017 966 3022
rect 2705 3017 2710 3022
rect 81 3012 190 3017
rect 961 3012 990 3017
rect 1081 3012 1142 3017
rect 985 3007 1086 3012
rect 1137 3007 1142 3012
rect 1217 3012 2190 3017
rect 2265 3012 2310 3017
rect 2361 3012 2614 3017
rect 2625 3012 2686 3017
rect 2705 3012 2758 3017
rect 1217 3007 1222 3012
rect 2865 3007 2870 3027
rect 2961 3022 3046 3027
rect 3121 3022 3646 3027
rect 3809 3027 3814 3032
rect 3809 3022 3910 3027
rect 3921 3022 4022 3027
rect 4177 3022 4278 3027
rect 3905 3017 3910 3022
rect 2897 3012 2958 3017
rect 2977 3012 3086 3017
rect 3153 3012 3214 3017
rect 3249 3012 3366 3017
rect 3681 3012 3774 3017
rect 3905 3012 4142 3017
rect 3385 3007 3662 3012
rect 337 3002 446 3007
rect 1137 3002 1222 3007
rect 1265 3002 2534 3007
rect 2665 3002 2870 3007
rect 3129 3002 3206 3007
rect 3233 3002 3390 3007
rect 3657 3002 3918 3007
rect 3961 3002 4078 3007
rect 2553 2997 2646 3002
rect 145 2992 230 2997
rect 313 2992 414 2997
rect 449 2992 558 2997
rect 577 2992 846 2997
rect 865 2992 1054 2997
rect 1241 2992 1390 2997
rect 1433 2992 1494 2997
rect 1529 2992 2254 2997
rect 2265 2992 2558 2997
rect 2641 2992 2782 2997
rect 3217 2992 3446 2997
rect 3465 2992 3678 2997
rect 3689 2992 3734 2997
rect 3761 2992 3846 2997
rect 3857 2992 4118 2997
rect 577 2987 582 2992
rect 417 2982 518 2987
rect 529 2982 582 2987
rect 841 2987 846 2992
rect 3441 2987 3446 2992
rect 841 2982 982 2987
rect 1065 2982 2126 2987
rect 2169 2982 2462 2987
rect 2529 2982 2870 2987
rect 3033 2982 3166 2987
rect 3297 2982 3390 2987
rect 3441 2982 3606 2987
rect 3617 2982 3710 2987
rect 3833 2982 4086 2987
rect 4201 2982 4334 2987
rect 601 2977 822 2982
rect 977 2977 1070 2982
rect 3601 2977 3606 2982
rect 529 2972 606 2977
rect 817 2972 958 2977
rect 1249 2972 1326 2977
rect 1465 2972 2214 2977
rect 2385 2972 2742 2977
rect 2753 2972 2798 2977
rect 2977 2972 3414 2977
rect 3601 2972 4246 2977
rect 1345 2967 1446 2972
rect 2209 2967 2390 2972
rect 3409 2967 3502 2972
rect 441 2962 1014 2967
rect 1081 2962 1190 2967
rect 1209 2962 1350 2967
rect 1441 2962 1726 2967
rect 1793 2962 1878 2967
rect 1889 2962 1998 2967
rect 2081 2962 2190 2967
rect 2409 2962 2606 2967
rect 2697 2962 2726 2967
rect 2881 2962 3182 2967
rect 3497 2962 4198 2967
rect 1081 2957 1086 2962
rect 369 2952 566 2957
rect 705 2952 878 2957
rect 1025 2952 1086 2957
rect 1185 2957 1190 2962
rect 2601 2957 2702 2962
rect 2881 2957 2886 2962
rect 3305 2957 3390 2962
rect 1185 2952 2198 2957
rect 2217 2952 2390 2957
rect 369 2947 374 2952
rect 585 2947 686 2952
rect 873 2947 1030 2952
rect 2217 2947 2222 2952
rect 185 2942 374 2947
rect 401 2942 590 2947
rect 681 2942 854 2947
rect 1097 2942 1246 2947
rect 1257 2942 1910 2947
rect 1993 2942 2022 2947
rect 2033 2942 2102 2947
rect 2113 2942 2142 2947
rect 2161 2942 2222 2947
rect 2385 2947 2390 2952
rect 2753 2952 2886 2957
rect 2913 2952 3310 2957
rect 3385 2952 3846 2957
rect 3937 2952 4254 2957
rect 2753 2947 2758 2952
rect 3841 2947 3942 2952
rect 2385 2942 2758 2947
rect 2993 2942 3214 2947
rect 3321 2942 3446 2947
rect 3537 2942 3630 2947
rect 3649 2942 3702 2947
rect 3737 2942 3822 2947
rect 3961 2942 4142 2947
rect 1905 2937 1998 2942
rect 2241 2937 2358 2942
rect 3649 2937 3654 2942
rect 4137 2937 4142 2942
rect 4265 2942 4294 2947
rect 4265 2937 4270 2942
rect 417 2932 806 2937
rect 921 2932 974 2937
rect 1185 2932 1214 2937
rect 1361 2932 1470 2937
rect 1569 2932 1646 2937
rect 1729 2932 1886 2937
rect 2057 2932 2246 2937
rect 2353 2932 2382 2937
rect 2929 2932 3006 2937
rect 3105 2932 3182 2937
rect 3193 2932 3222 2937
rect 3465 2932 3654 2937
rect 1233 2927 1342 2932
rect 2681 2927 2822 2932
rect 3681 2927 3686 2937
rect 3729 2932 3846 2937
rect 3937 2932 4046 2937
rect 4137 2932 4270 2937
rect 657 2922 766 2927
rect 785 2922 1238 2927
rect 1337 2922 1798 2927
rect 1849 2922 1894 2927
rect 2017 2922 2630 2927
rect 2657 2922 2686 2927
rect 2817 2922 2846 2927
rect 3009 2922 3230 2927
rect 3265 2922 3334 2927
rect 3353 2922 3446 2927
rect 3681 2922 3726 2927
rect 545 2917 638 2922
rect 657 2917 662 2922
rect 441 2912 550 2917
rect 633 2912 662 2917
rect 737 2917 742 2922
rect 737 2912 886 2917
rect 913 2912 1038 2917
rect 1121 2912 1446 2917
rect 1457 2912 2006 2917
rect 2017 2912 2022 2922
rect 2625 2917 2630 2922
rect 3353 2917 3358 2922
rect 2105 2912 2166 2917
rect 2241 2912 2310 2917
rect 2625 2912 2646 2917
rect 2657 2912 2742 2917
rect 2769 2912 2910 2917
rect 3017 2912 3358 2917
rect 3441 2917 3446 2922
rect 3553 2917 3662 2922
rect 3441 2912 3558 2917
rect 3657 2912 3894 2917
rect 3905 2912 3990 2917
rect 4065 2912 4142 2917
rect 4233 2912 4318 2917
rect 1441 2907 1446 2912
rect 2641 2907 2646 2912
rect 3889 2907 3894 2912
rect 233 2902 302 2907
rect 561 2902 1342 2907
rect 1377 2902 1422 2907
rect 1441 2902 2094 2907
rect 2177 2902 2422 2907
rect 449 2897 542 2902
rect 2089 2897 2182 2902
rect 2417 2897 2422 2902
rect 2481 2902 2542 2907
rect 2553 2902 2622 2907
rect 2641 2902 2854 2907
rect 2881 2902 3150 2907
rect 3161 2902 3486 2907
rect 3593 2902 3686 2907
rect 3889 2902 3918 2907
rect 4081 2902 4278 2907
rect 2481 2897 2486 2902
rect 3481 2897 3574 2902
rect 3713 2897 3814 2902
rect 4081 2897 4086 2902
rect 345 2892 454 2897
rect 537 2892 910 2897
rect 1009 2892 1782 2897
rect 1793 2892 2070 2897
rect 2225 2892 2326 2897
rect 2417 2892 2486 2897
rect 2817 2892 3422 2897
rect 3569 2892 3718 2897
rect 3809 2892 3838 2897
rect 3897 2892 4086 2897
rect 4097 2892 4206 2897
rect 185 2882 334 2887
rect 329 2877 334 2882
rect 465 2882 750 2887
rect 857 2882 886 2887
rect 897 2882 942 2887
rect 961 2882 1150 2887
rect 1161 2882 1246 2887
rect 1281 2882 1366 2887
rect 1441 2882 1526 2887
rect 1641 2882 1670 2887
rect 1721 2882 2062 2887
rect 2169 2882 2254 2887
rect 2625 2882 2798 2887
rect 2873 2882 2966 2887
rect 3217 2882 3558 2887
rect 3673 2882 3862 2887
rect 4073 2882 4374 2887
rect 465 2877 470 2882
rect 745 2877 862 2882
rect 1281 2877 1286 2882
rect 1521 2877 1606 2882
rect 2273 2877 2374 2882
rect 2625 2877 2630 2882
rect 329 2872 470 2877
rect 489 2872 726 2877
rect 905 2872 1094 2877
rect 1153 2872 1286 2877
rect 1297 2872 1502 2877
rect 1601 2872 2278 2877
rect 2369 2872 2398 2877
rect 2497 2872 2630 2877
rect 2793 2877 2798 2882
rect 2985 2877 3102 2882
rect 3553 2877 3678 2882
rect 2793 2872 2926 2877
rect 2937 2872 2990 2877
rect 3097 2872 3126 2877
rect 2665 2867 2774 2872
rect 3321 2867 3510 2872
rect 4017 2867 4182 2872
rect 113 2862 214 2867
rect 505 2862 702 2867
rect 849 2862 1014 2867
rect 1113 2862 1454 2867
rect 1489 2862 1862 2867
rect 2105 2862 2286 2867
rect 2297 2862 2366 2867
rect 2641 2862 2670 2867
rect 2769 2862 3326 2867
rect 3505 2862 3534 2867
rect 3553 2862 3622 2867
rect 3729 2862 3878 2867
rect 3993 2862 4022 2867
rect 4177 2862 4238 2867
rect 721 2857 830 2862
rect 3553 2857 3558 2862
rect 233 2852 342 2857
rect 361 2852 414 2857
rect 569 2852 726 2857
rect 825 2852 3110 2857
rect 3265 2852 3558 2857
rect 3617 2857 3622 2862
rect 3617 2852 4166 2857
rect 233 2847 238 2852
rect 201 2842 238 2847
rect 337 2847 342 2852
rect 3129 2847 3246 2852
rect 337 2842 718 2847
rect 761 2842 790 2847
rect 841 2842 958 2847
rect 1177 2842 1278 2847
rect 1289 2842 1494 2847
rect 1537 2842 1766 2847
rect 1777 2842 1814 2847
rect 1825 2842 1902 2847
rect 2097 2842 2150 2847
rect 2177 2842 2334 2847
rect 2441 2842 2510 2847
rect 2609 2842 2758 2847
rect 2873 2842 2918 2847
rect 2945 2842 3134 2847
rect 3241 2842 3294 2847
rect 3369 2842 3454 2847
rect 3497 2842 3630 2847
rect 3793 2842 3910 2847
rect 1537 2837 1542 2842
rect 3649 2837 3742 2842
rect 601 2832 758 2837
rect 793 2832 822 2837
rect 833 2832 862 2837
rect 1033 2832 1206 2837
rect 1273 2832 1542 2837
rect 1561 2832 1638 2837
rect 1697 2832 1774 2837
rect 1793 2832 1934 2837
rect 1961 2832 2086 2837
rect 2201 2832 2246 2837
rect 2289 2832 2366 2837
rect 2385 2832 2470 2837
rect 2513 2832 2742 2837
rect 2777 2832 2814 2837
rect 2865 2832 3654 2837
rect 3737 2832 3766 2837
rect 4065 2832 4150 2837
rect 329 2827 438 2832
rect 2081 2827 2206 2832
rect 137 2822 230 2827
rect 257 2822 334 2827
rect 433 2822 462 2827
rect 505 2822 550 2827
rect 561 2822 654 2827
rect 721 2822 854 2827
rect 953 2822 1094 2827
rect 1161 2822 1206 2827
rect 1233 2822 1294 2827
rect 1305 2822 1374 2827
rect 1441 2822 1550 2827
rect 1577 2822 1622 2827
rect 1641 2822 1662 2827
rect 1761 2822 1830 2827
rect 1889 2822 1966 2827
rect 1977 2822 2022 2827
rect 2225 2817 2230 2827
rect 313 2812 606 2817
rect 625 2812 1150 2817
rect 1249 2812 1702 2817
rect 1713 2812 1790 2817
rect 2009 2812 2134 2817
rect 2169 2812 2230 2817
rect 2241 2817 2246 2832
rect 2385 2827 2390 2832
rect 2737 2827 2742 2832
rect 2257 2822 2294 2827
rect 2321 2822 2390 2827
rect 2321 2817 2326 2822
rect 2401 2817 2406 2827
rect 2601 2822 2638 2827
rect 2689 2822 2718 2827
rect 2737 2822 2814 2827
rect 2889 2822 3206 2827
rect 3233 2822 3286 2827
rect 3313 2822 3438 2827
rect 3505 2822 3526 2827
rect 3633 2822 3710 2827
rect 3865 2822 3934 2827
rect 4081 2822 4126 2827
rect 3505 2817 3510 2822
rect 2241 2812 2326 2817
rect 2337 2812 2406 2817
rect 2545 2812 3510 2817
rect 3529 2812 4038 2817
rect 4185 2812 4294 2817
rect 625 2807 630 2812
rect 1145 2807 1254 2812
rect 1809 2807 1990 2812
rect 2545 2807 2550 2812
rect 4185 2807 4190 2812
rect 201 2802 238 2807
rect 289 2802 534 2807
rect 609 2802 630 2807
rect 639 2802 678 2807
rect 721 2802 806 2807
rect 865 2802 902 2807
rect 985 2802 1030 2807
rect 1273 2802 1318 2807
rect 1353 2802 1398 2807
rect 1417 2802 1438 2807
rect 1497 2802 1814 2807
rect 1985 2802 2550 2807
rect 2561 2802 2654 2807
rect 2705 2802 2758 2807
rect 2769 2802 2942 2807
rect 3001 2802 3150 2807
rect 3177 2802 3270 2807
rect 3289 2802 3318 2807
rect 639 2797 644 2802
rect 721 2797 726 2802
rect 2753 2797 2758 2802
rect 3393 2797 3398 2807
rect 3489 2802 3542 2807
rect 3609 2802 3646 2807
rect 4033 2802 4150 2807
rect 4161 2802 4190 2807
rect 4289 2807 4294 2812
rect 4289 2802 4318 2807
rect 3841 2797 3966 2802
rect 4033 2797 4038 2802
rect 209 2792 342 2797
rect 369 2792 644 2797
rect 649 2792 726 2797
rect 737 2792 982 2797
rect 1001 2792 1038 2797
rect 1049 2792 1086 2797
rect 1105 2792 1182 2797
rect 1201 2792 1270 2797
rect 1305 2792 1326 2797
rect 1337 2792 1390 2797
rect 1425 2792 2598 2797
rect 2617 2792 2734 2797
rect 2753 2792 2838 2797
rect 2857 2792 2918 2797
rect 3113 2792 3262 2797
rect 3393 2792 3526 2797
rect 3577 2792 3774 2797
rect 3785 2792 3846 2797
rect 3961 2792 3990 2797
rect 4001 2792 4062 2797
rect 4089 2792 4214 2797
rect 337 2787 342 2792
rect 1105 2787 1110 2792
rect 2833 2787 2838 2792
rect 3393 2787 3398 2792
rect 3521 2787 3526 2792
rect 4001 2787 4006 2792
rect 337 2782 430 2787
rect 465 2782 886 2787
rect 993 2782 1030 2787
rect 1041 2782 1110 2787
rect 1121 2782 1446 2787
rect 1465 2782 1494 2787
rect 1513 2782 1534 2787
rect 1577 2782 1638 2787
rect 1697 2782 2510 2787
rect 2689 2782 2822 2787
rect 2833 2782 3006 2787
rect 3017 2782 3126 2787
rect 3145 2782 3398 2787
rect 3417 2782 3510 2787
rect 3521 2782 4006 2787
rect 4025 2782 4374 2787
rect 1041 2777 1046 2782
rect 281 2772 446 2777
rect 537 2772 678 2777
rect 689 2772 726 2777
rect 745 2772 1046 2777
rect 1057 2772 1766 2777
rect 1825 2772 1878 2777
rect 1921 2772 1982 2777
rect 1993 2772 2014 2777
rect 2025 2772 2078 2777
rect 2097 2772 2198 2777
rect 2225 2772 2278 2777
rect 2329 2772 2446 2777
rect 2481 2772 2830 2777
rect 2849 2772 3094 2777
rect 3121 2772 3126 2782
rect 3505 2777 3510 2782
rect 3161 2772 3238 2777
rect 3449 2772 3486 2777
rect 3505 2772 3542 2777
rect 3585 2772 3702 2777
rect 3745 2772 3918 2777
rect 1057 2767 1062 2772
rect 1761 2767 1766 2772
rect 3257 2767 3430 2772
rect 185 2762 246 2767
rect 257 2762 422 2767
rect 513 2762 566 2767
rect 593 2762 678 2767
rect 697 2762 814 2767
rect 841 2762 862 2767
rect 881 2762 990 2767
rect 1025 2762 1062 2767
rect 1137 2762 1238 2767
rect 1257 2762 1286 2767
rect 1361 2762 1454 2767
rect 1465 2762 1606 2767
rect 1681 2762 1742 2767
rect 1761 2762 3262 2767
rect 3425 2762 3670 2767
rect 3745 2757 3750 2772
rect 3913 2767 3918 2772
rect 4025 2772 4054 2777
rect 4081 2772 4270 2777
rect 4025 2767 4030 2772
rect 3817 2762 3886 2767
rect 3913 2762 4030 2767
rect 4073 2762 4326 2767
rect 217 2752 926 2757
rect 945 2752 1006 2757
rect 1217 2752 1670 2757
rect 1689 2752 1750 2757
rect 1769 2752 1878 2757
rect 1905 2752 1950 2757
rect 2009 2752 2070 2757
rect 2113 2752 2166 2757
rect 2233 2752 2374 2757
rect 2417 2752 2486 2757
rect 2537 2752 2558 2757
rect 2569 2752 2638 2757
rect 2681 2752 2886 2757
rect 2953 2752 3006 2757
rect 3017 2752 3750 2757
rect 3769 2752 3894 2757
rect 4113 2752 4214 2757
rect 1025 2747 1198 2752
rect 81 2742 102 2747
rect 121 2742 278 2747
rect 353 2742 438 2747
rect 449 2742 478 2747
rect 521 2742 590 2747
rect 641 2742 662 2747
rect 681 2742 710 2747
rect 721 2742 774 2747
rect 785 2742 1030 2747
rect 1193 2742 3758 2747
rect 3953 2742 4054 2747
rect 4185 2742 4286 2747
rect 97 2737 102 2742
rect 449 2737 454 2742
rect 3953 2737 3958 2742
rect 97 2732 126 2737
rect 265 2732 1366 2737
rect 1409 2732 1446 2737
rect 1481 2732 2422 2737
rect 2433 2732 3134 2737
rect 3313 2732 3910 2737
rect 3929 2732 3958 2737
rect 4049 2737 4054 2742
rect 4049 2732 4086 2737
rect 4137 2732 4190 2737
rect 4201 2732 4270 2737
rect 121 2727 270 2732
rect 289 2722 742 2727
rect 753 2722 934 2727
rect 977 2722 982 2732
rect 1361 2727 1366 2732
rect 2417 2727 2422 2732
rect 3153 2727 3246 2732
rect 3313 2727 3318 2732
rect 3393 2727 3398 2732
rect 1041 2722 1102 2727
rect 1097 2717 1102 2722
rect 1153 2722 1198 2727
rect 1233 2722 1286 2727
rect 1361 2722 1382 2727
rect 1409 2722 1502 2727
rect 1625 2722 1846 2727
rect 1937 2722 1998 2727
rect 2097 2722 2190 2727
rect 2297 2722 2350 2727
rect 2417 2722 2502 2727
rect 2593 2722 2710 2727
rect 2721 2722 3062 2727
rect 3073 2722 3158 2727
rect 3241 2722 3318 2727
rect 3337 2722 3382 2727
rect 3393 2722 3422 2727
rect 3465 2722 3526 2727
rect 3569 2722 3718 2727
rect 3737 2722 3814 2727
rect 3905 2722 3910 2732
rect 4081 2727 4086 2732
rect 4081 2722 4342 2727
rect 1153 2717 1158 2722
rect 3905 2717 4062 2722
rect 121 2712 230 2717
rect 417 2712 454 2717
rect 473 2712 862 2717
rect 977 2712 1086 2717
rect 1097 2712 1134 2717
rect 1145 2712 1158 2717
rect 1217 2712 1262 2717
rect 1337 2712 2766 2717
rect 2785 2712 2822 2717
rect 2865 2712 3502 2717
rect 3665 2712 3798 2717
rect 4057 2712 4182 2717
rect 4193 2712 4278 2717
rect 4337 2712 4342 2722
rect 1145 2707 1150 2712
rect 3521 2707 3646 2712
rect 201 2702 294 2707
rect 369 2702 390 2707
rect 513 2702 542 2707
rect 553 2702 598 2707
rect 697 2702 950 2707
rect 961 2702 1062 2707
rect 1081 2702 1150 2707
rect 1161 2702 1206 2707
rect 1241 2702 1486 2707
rect 1513 2702 1606 2707
rect 1617 2702 1654 2707
rect 1665 2702 1766 2707
rect 1817 2702 1846 2707
rect 1865 2702 1950 2707
rect 2081 2702 2422 2707
rect 2433 2702 2486 2707
rect 2609 2702 2678 2707
rect 2705 2702 3014 2707
rect 3057 2702 3094 2707
rect 3209 2702 3278 2707
rect 3289 2702 3526 2707
rect 3641 2702 3974 2707
rect 3985 2702 4062 2707
rect 4121 2702 4230 2707
rect 1617 2697 1622 2702
rect 1969 2697 2062 2702
rect 281 2692 1494 2697
rect 1537 2692 1574 2697
rect 1593 2692 1622 2697
rect 1633 2692 1974 2697
rect 2057 2692 2550 2697
rect 2593 2692 2638 2697
rect 2681 2692 2990 2697
rect 3009 2687 3014 2702
rect 3969 2697 3974 2702
rect 3033 2692 3190 2697
rect 3201 2692 3302 2697
rect 3337 2692 3358 2697
rect 3369 2692 3486 2697
rect 3521 2692 3558 2697
rect 3593 2692 3662 2697
rect 3721 2692 3774 2697
rect 3817 2692 3958 2697
rect 3969 2692 4206 2697
rect 65 2682 270 2687
rect 457 2682 582 2687
rect 593 2682 654 2687
rect 689 2682 718 2687
rect 785 2682 822 2687
rect 873 2682 1126 2687
rect 1137 2682 1214 2687
rect 1265 2682 1294 2687
rect 1305 2682 1366 2687
rect 1393 2682 1502 2687
rect 1553 2682 2590 2687
rect 2737 2682 2838 2687
rect 2921 2682 2974 2687
rect 3009 2682 3102 2687
rect 3113 2682 3214 2687
rect 3265 2682 3406 2687
rect 3473 2682 3518 2687
rect 3953 2682 3990 2687
rect 4001 2682 4102 2687
rect 265 2677 462 2682
rect 1265 2677 1270 2682
rect 2609 2677 2718 2682
rect 2737 2677 2742 2682
rect 3577 2677 3702 2682
rect 3745 2677 3878 2682
rect 3953 2677 3958 2682
rect 481 2672 518 2677
rect 561 2672 766 2677
rect 865 2672 902 2677
rect 945 2672 1070 2677
rect 1105 2672 1198 2677
rect 1217 2672 1270 2677
rect 1281 2672 1718 2677
rect 1833 2672 1878 2677
rect 1889 2672 2614 2677
rect 2713 2672 2742 2677
rect 2761 2672 3398 2677
rect 3409 2672 3582 2677
rect 3697 2672 3750 2677
rect 3873 2672 3958 2677
rect 3969 2672 4014 2677
rect 161 2662 478 2667
rect 513 2662 630 2667
rect 689 2662 1998 2667
rect 2057 2662 2134 2667
rect 2145 2662 2198 2667
rect 2209 2662 2230 2667
rect 2241 2662 2446 2667
rect 2457 2662 2534 2667
rect 2585 2662 3598 2667
rect 3609 2662 3670 2667
rect 3761 2662 3950 2667
rect 4033 2662 4166 2667
rect 4185 2662 4230 2667
rect 689 2657 694 2662
rect 4033 2657 4038 2662
rect 185 2652 214 2657
rect 209 2647 214 2652
rect 425 2652 694 2657
rect 713 2652 798 2657
rect 817 2652 894 2657
rect 1017 2652 1086 2657
rect 1153 2652 1470 2657
rect 1489 2652 2518 2657
rect 2553 2652 2702 2657
rect 2753 2652 4038 2657
rect 4161 2657 4166 2662
rect 4161 2652 4198 2657
rect 4249 2652 4342 2657
rect 425 2647 430 2652
rect 889 2647 998 2652
rect 4249 2647 4254 2652
rect 209 2642 430 2647
rect 449 2642 566 2647
rect 577 2642 638 2647
rect 681 2642 766 2647
rect 825 2642 870 2647
rect 993 2642 1030 2647
rect 1073 2642 1246 2647
rect 1297 2642 2006 2647
rect 2113 2642 2686 2647
rect 2729 2642 2782 2647
rect 2849 2642 3022 2647
rect 3097 2642 3414 2647
rect 3473 2642 3710 2647
rect 3753 2642 3798 2647
rect 3809 2642 4254 2647
rect 4337 2647 4342 2652
rect 4337 2642 4366 2647
rect 577 2637 582 2642
rect 2001 2637 2118 2642
rect 449 2632 526 2637
rect 545 2632 582 2637
rect 697 2632 1014 2637
rect 1097 2632 1374 2637
rect 1425 2632 1446 2637
rect 1529 2632 1574 2637
rect 1617 2632 1646 2637
rect 1657 2632 1822 2637
rect 1921 2632 1942 2637
rect 1961 2632 1982 2637
rect 2137 2632 2358 2637
rect 2369 2632 3390 2637
rect 3489 2632 3614 2637
rect 593 2627 702 2632
rect 1009 2627 1014 2632
rect 2369 2627 2374 2632
rect 3385 2627 3494 2632
rect 3609 2627 3614 2632
rect 3721 2632 3822 2637
rect 4025 2632 4110 2637
rect 4145 2632 4222 2637
rect 3721 2627 3726 2632
rect 3817 2627 4030 2632
rect 4145 2627 4150 2632
rect 209 2622 406 2627
rect 433 2622 598 2627
rect 721 2622 990 2627
rect 1009 2622 1694 2627
rect 1713 2622 1918 2627
rect 1961 2622 2062 2627
rect 2081 2622 2374 2627
rect 2393 2622 2438 2627
rect 2505 2622 3246 2627
rect 3321 2622 3366 2627
rect 3513 2622 3590 2627
rect 3609 2622 3726 2627
rect 3745 2622 3798 2627
rect 4049 2622 4150 2627
rect 4169 2622 4342 2627
rect 2081 2617 2086 2622
rect 233 2612 446 2617
rect 489 2612 558 2617
rect 585 2612 2086 2617
rect 2105 2612 2182 2617
rect 2193 2612 2286 2617
rect 2305 2612 2334 2617
rect 2353 2612 2406 2617
rect 2497 2612 3414 2617
rect 3521 2612 3542 2617
rect 3801 2612 3846 2617
rect 3961 2612 4030 2617
rect 4057 2612 4118 2617
rect 4353 2612 4446 2617
rect 3681 2607 3782 2612
rect 3961 2607 3966 2612
rect 193 2602 326 2607
rect 353 2602 374 2607
rect 401 2602 950 2607
rect 257 2592 350 2597
rect 401 2592 406 2602
rect 945 2597 950 2602
rect 1009 2602 1678 2607
rect 1689 2602 2638 2607
rect 2673 2602 2870 2607
rect 2985 2602 3126 2607
rect 3185 2602 3222 2607
rect 3241 2602 3366 2607
rect 3385 2602 3462 2607
rect 3489 2602 3686 2607
rect 3777 2602 3966 2607
rect 4025 2607 4030 2612
rect 4113 2607 4358 2612
rect 4025 2602 4094 2607
rect 1009 2597 1014 2602
rect 441 2592 542 2597
rect 697 2592 734 2597
rect 849 2592 878 2597
rect 945 2592 1014 2597
rect 1153 2592 1182 2597
rect 1225 2592 1254 2597
rect 1273 2592 1374 2597
rect 1473 2592 2846 2597
rect 2873 2592 2926 2597
rect 2937 2592 3062 2597
rect 3089 2592 3254 2597
rect 3281 2592 3398 2597
rect 3497 2592 3606 2597
rect 3697 2592 3822 2597
rect 3977 2592 4174 2597
rect 4201 2592 4278 2597
rect 561 2587 678 2592
rect 1033 2587 1134 2592
rect 3841 2587 3958 2592
rect 329 2582 438 2587
rect 449 2582 566 2587
rect 673 2582 1038 2587
rect 1129 2582 1654 2587
rect 1673 2582 1750 2587
rect 1809 2582 1886 2587
rect 1921 2582 1990 2587
rect 2001 2582 3846 2587
rect 3953 2582 4038 2587
rect 4049 2582 4102 2587
rect 4113 2582 4222 2587
rect 4249 2582 4294 2587
rect 4049 2577 4054 2582
rect 361 2572 750 2577
rect 817 2572 846 2577
rect 857 2572 894 2577
rect 921 2572 1094 2577
rect 1145 2572 1238 2577
rect 1257 2572 1286 2577
rect 1329 2572 1366 2577
rect 1393 2572 2502 2577
rect 2513 2572 3294 2577
rect 3401 2572 3830 2577
rect 3849 2572 3926 2577
rect 3985 2572 4014 2577
rect 4025 2572 4054 2577
rect 4105 2572 4174 2577
rect 1329 2567 1334 2572
rect 3825 2567 3830 2572
rect 337 2562 494 2567
rect 505 2562 566 2567
rect 585 2562 606 2567
rect 617 2562 654 2567
rect 689 2562 902 2567
rect 913 2562 958 2567
rect 977 2562 1334 2567
rect 1345 2562 1382 2567
rect 1449 2562 1542 2567
rect 1569 2562 1686 2567
rect 1713 2562 1838 2567
rect 1849 2562 1886 2567
rect 1905 2562 2054 2567
rect 2097 2562 2182 2567
rect 2201 2562 2230 2567
rect 2249 2562 2270 2567
rect 2281 2562 2366 2567
rect 2377 2562 2398 2567
rect 2409 2562 2486 2567
rect 2529 2562 2550 2567
rect 2649 2562 2718 2567
rect 2809 2562 3014 2567
rect 3057 2562 3174 2567
rect 3185 2562 3278 2567
rect 3313 2562 3334 2567
rect 3377 2562 3454 2567
rect 3513 2562 3542 2567
rect 3649 2562 3774 2567
rect 3825 2562 4006 2567
rect 4017 2562 4102 2567
rect 4113 2562 4374 2567
rect 3185 2557 3190 2562
rect 3313 2557 3318 2562
rect 65 2552 94 2557
rect 113 2552 262 2557
rect 393 2552 702 2557
rect 809 2552 862 2557
rect 961 2552 1070 2557
rect 1177 2552 1414 2557
rect 1465 2552 2118 2557
rect 2225 2552 3190 2557
rect 3209 2552 3318 2557
rect 3337 2552 3358 2557
rect 3465 2552 3534 2557
rect 3553 2552 3646 2557
rect 3705 2552 3734 2557
rect 3761 2552 3974 2557
rect 4033 2552 4150 2557
rect 65 2527 70 2552
rect 113 2547 118 2552
rect 2113 2547 2230 2552
rect 3729 2547 3734 2552
rect 89 2542 118 2547
rect 137 2542 222 2547
rect 273 2542 422 2547
rect 457 2542 1710 2547
rect 1761 2537 1766 2547
rect 1809 2542 1998 2547
rect 2017 2542 2094 2547
rect 2249 2542 2286 2547
rect 2297 2542 2726 2547
rect 2761 2542 2790 2547
rect 2801 2542 2830 2547
rect 2913 2542 3046 2547
rect 3089 2542 3150 2547
rect 3169 2542 3190 2547
rect 3209 2542 3358 2547
rect 3393 2542 3486 2547
rect 3633 2542 3670 2547
rect 3729 2542 3790 2547
rect 3817 2542 3870 2547
rect 4041 2542 4078 2547
rect 4089 2542 4150 2547
rect 2297 2537 2302 2542
rect 3185 2537 3190 2542
rect 3393 2537 3398 2542
rect 305 2532 374 2537
rect 465 2532 494 2537
rect 569 2532 734 2537
rect 793 2532 838 2537
rect 857 2532 894 2537
rect 953 2532 982 2537
rect 1097 2532 1190 2537
rect 1201 2532 1310 2537
rect 185 2527 286 2532
rect 1201 2527 1206 2532
rect 1321 2527 1326 2537
rect 1337 2532 1398 2537
rect 1449 2532 1478 2537
rect 1537 2532 1646 2537
rect 1665 2532 1766 2537
rect 1793 2532 1878 2537
rect 1921 2532 1974 2537
rect 2009 2532 2054 2537
rect 2209 2532 2302 2537
rect 2377 2532 2438 2537
rect 2457 2532 2510 2537
rect 65 2522 190 2527
rect 281 2522 814 2527
rect 985 2522 1054 2527
rect 1121 2522 1206 2527
rect 1289 2522 1326 2527
rect 1529 2522 1566 2527
rect 1649 2522 1774 2527
rect 1828 2522 1854 2527
rect 833 2517 934 2522
rect 1121 2517 1126 2522
rect 1828 2517 1833 2522
rect 1873 2517 1878 2532
rect 2073 2527 2190 2532
rect 2545 2527 2550 2537
rect 2609 2532 3062 2537
rect 3185 2532 3398 2537
rect 3409 2532 3462 2537
rect 3473 2532 3638 2537
rect 3729 2532 3782 2537
rect 3473 2527 3478 2532
rect 4193 2527 4198 2547
rect 4217 2542 4310 2547
rect 1937 2522 2078 2527
rect 2185 2522 3478 2527
rect 3489 2522 3606 2527
rect 3625 2522 3734 2527
rect 4081 2522 4158 2527
rect 4193 2522 4222 2527
rect 3489 2517 3494 2522
rect 201 2512 710 2517
rect 721 2512 838 2517
rect 929 2512 958 2517
rect 993 2507 998 2517
rect 1033 2512 1054 2517
rect 1097 2512 1126 2517
rect 1161 2512 1214 2517
rect 1225 2512 1798 2517
rect 1817 2512 1833 2517
rect 1857 2512 1878 2517
rect 1945 2512 2470 2517
rect 2481 2512 2510 2517
rect 2625 2512 2646 2517
rect 2745 2512 2838 2517
rect 2873 2512 2990 2517
rect 3049 2512 3110 2517
rect 3129 2512 3238 2517
rect 3297 2512 3494 2517
rect 3513 2512 3590 2517
rect 3105 2507 3110 2512
rect 3601 2507 3606 2522
rect 3681 2512 3742 2517
rect 3841 2512 3918 2517
rect 3937 2512 4062 2517
rect 4081 2512 4150 2517
rect 4177 2512 4246 2517
rect 3937 2507 3942 2512
rect 121 2502 542 2507
rect 569 2502 662 2507
rect 673 2502 998 2507
rect 1009 2502 1078 2507
rect 1137 2502 1246 2507
rect 1321 2502 1358 2507
rect 1433 2502 1750 2507
rect 1761 2502 1814 2507
rect 1833 2502 1902 2507
rect 1937 2502 1974 2507
rect 1993 2502 2038 2507
rect 2081 2502 2694 2507
rect 2817 2502 2878 2507
rect 2897 2502 2942 2507
rect 2961 2502 2990 2507
rect 3033 2502 3094 2507
rect 3105 2502 3254 2507
rect 3409 2502 3574 2507
rect 3601 2502 3854 2507
rect 3913 2502 3942 2507
rect 4057 2507 4062 2512
rect 4057 2502 4190 2507
rect 527 2497 532 2502
rect 673 2497 678 2502
rect 3249 2497 3254 2502
rect 3305 2497 3414 2502
rect 209 2492 286 2497
rect 281 2487 286 2492
rect 345 2492 510 2497
rect 527 2492 678 2497
rect 769 2492 2470 2497
rect 2497 2492 3222 2497
rect 3249 2492 3310 2497
rect 3425 2492 3462 2497
rect 3473 2492 3806 2497
rect 345 2487 350 2492
rect 3473 2487 3478 2492
rect 281 2482 350 2487
rect 433 2482 502 2487
rect 545 2482 590 2487
rect 617 2482 894 2487
rect 929 2482 2582 2487
rect 2601 2482 3478 2487
rect 3489 2482 3558 2487
rect 3569 2482 3718 2487
rect 385 2472 462 2477
rect 497 2467 502 2482
rect 2577 2477 2582 2482
rect 3713 2477 3718 2482
rect 3801 2482 3830 2487
rect 3849 2482 4230 2487
rect 3801 2477 3806 2482
rect 521 2472 766 2477
rect 801 2472 902 2477
rect 913 2472 1046 2477
rect 1089 2467 1094 2477
rect 1129 2472 1182 2477
rect 1201 2472 1750 2477
rect 1817 2472 2038 2477
rect 2049 2472 2094 2477
rect 2105 2472 2198 2477
rect 2257 2472 2342 2477
rect 2425 2472 2494 2477
rect 2577 2472 2638 2477
rect 2697 2472 2790 2477
rect 2833 2472 3478 2477
rect 3513 2472 3550 2477
rect 3585 2472 3694 2477
rect 3713 2472 3806 2477
rect 3825 2467 3830 2482
rect 3865 2472 3910 2477
rect 497 2462 614 2467
rect 649 2462 694 2467
rect 737 2462 870 2467
rect 889 2462 1094 2467
rect 1105 2462 1190 2467
rect 1217 2462 1262 2467
rect 1273 2462 2454 2467
rect 2465 2462 3622 2467
rect 3825 2462 4206 2467
rect 737 2457 742 2462
rect 2449 2457 2454 2462
rect 457 2452 518 2457
rect 673 2452 742 2457
rect 753 2452 1934 2457
rect 1985 2452 2142 2457
rect 2161 2452 2214 2457
rect 2233 2452 2302 2457
rect 2313 2452 2382 2457
rect 2409 2452 2438 2457
rect 2449 2452 2934 2457
rect 2945 2452 3006 2457
rect 3025 2452 3142 2457
rect 3217 2452 3310 2457
rect 3433 2452 3470 2457
rect 3529 2452 3646 2457
rect 3665 2452 3942 2457
rect 1985 2447 1990 2452
rect 3665 2447 3670 2452
rect 249 2442 390 2447
rect 505 2442 582 2447
rect 673 2442 830 2447
rect 837 2442 854 2447
rect 865 2442 990 2447
rect 1089 2442 1198 2447
rect 1209 2442 1414 2447
rect 1473 2442 1558 2447
rect 1593 2442 1614 2447
rect 1625 2442 1990 2447
rect 2065 2442 2838 2447
rect 2937 2442 3670 2447
rect 3689 2442 3718 2447
rect 3833 2442 3958 2447
rect 3977 2442 4062 2447
rect 249 2437 254 2442
rect 65 2432 86 2437
rect 177 2432 254 2437
rect 385 2437 390 2442
rect 673 2437 678 2442
rect 837 2437 842 2442
rect 865 2437 870 2442
rect 3977 2437 3982 2442
rect 385 2432 414 2437
rect 449 2432 678 2437
rect 697 2432 822 2437
rect 833 2432 842 2437
rect 849 2432 870 2437
rect 889 2432 2222 2437
rect 2249 2432 2310 2437
rect 2321 2432 2350 2437
rect 2385 2432 2654 2437
rect 2777 2432 3286 2437
rect 3409 2432 3438 2437
rect 3449 2432 3486 2437
rect 3545 2432 3686 2437
rect 3801 2432 3982 2437
rect 4057 2437 4062 2442
rect 4057 2432 4086 2437
rect 4161 2432 4254 2437
rect 65 2397 70 2432
rect 833 2427 838 2432
rect 137 2422 222 2427
rect 385 2422 782 2427
rect 809 2422 838 2427
rect 849 2422 2566 2427
rect 2609 2422 2678 2427
rect 2769 2422 3974 2427
rect 4001 2422 4070 2427
rect 385 2417 390 2422
rect 2769 2417 2774 2422
rect 4081 2417 4086 2432
rect 4225 2422 4302 2427
rect 89 2412 118 2417
rect 65 2392 94 2397
rect 65 2377 70 2392
rect 113 2387 118 2412
rect 265 2412 390 2417
rect 399 2412 542 2417
rect 577 2412 1766 2417
rect 1849 2412 1910 2417
rect 1945 2412 1990 2417
rect 2041 2412 2774 2417
rect 2817 2412 2934 2417
rect 2977 2412 2998 2417
rect 3057 2412 3982 2417
rect 4081 2412 4142 2417
rect 265 2407 270 2412
rect 169 2402 270 2407
rect 399 2397 404 2412
rect 2817 2407 2822 2412
rect 409 2402 446 2407
rect 481 2402 622 2407
rect 665 2402 702 2407
rect 753 2402 822 2407
rect 849 2402 910 2407
rect 953 2402 1102 2407
rect 1129 2402 1182 2407
rect 1193 2402 1334 2407
rect 1361 2402 1390 2407
rect 1401 2402 1454 2407
rect 1465 2402 1558 2407
rect 1593 2402 1670 2407
rect 1745 2402 2158 2407
rect 2185 2402 2694 2407
rect 2753 2402 2774 2407
rect 2801 2402 2822 2407
rect 2841 2402 2894 2407
rect 2905 2402 2966 2407
rect 2985 2402 3094 2407
rect 3217 2402 3910 2407
rect 4009 2402 4094 2407
rect 4177 2402 4222 2407
rect 153 2392 182 2397
rect 89 2382 118 2387
rect 177 2387 182 2392
rect 257 2392 404 2397
rect 457 2392 598 2397
rect 641 2392 670 2397
rect 769 2392 2102 2397
rect 2209 2392 3590 2397
rect 3665 2392 3742 2397
rect 3777 2392 3846 2397
rect 3857 2392 3862 2402
rect 4073 2392 4358 2397
rect 257 2387 262 2392
rect 593 2387 598 2392
rect 2097 2387 2214 2392
rect 177 2382 262 2387
rect 505 2382 582 2387
rect 593 2382 726 2387
rect 857 2382 1014 2387
rect 1033 2382 1126 2387
rect 1137 2382 1158 2387
rect 1185 2382 1238 2387
rect 1273 2382 1294 2387
rect 1313 2382 1422 2387
rect 1457 2382 1486 2387
rect 1505 2382 1542 2387
rect 1569 2382 1710 2387
rect 1769 2382 1830 2387
rect 1857 2382 2078 2387
rect 2233 2382 2430 2387
rect 2449 2382 2510 2387
rect 2561 2382 2934 2387
rect 2945 2382 3006 2387
rect 3025 2382 3078 2387
rect 3121 2382 3182 2387
rect 3201 2382 3262 2387
rect 3313 2382 3502 2387
rect 3609 2382 3798 2387
rect 3905 2382 3974 2387
rect 4017 2382 4038 2387
rect 4049 2382 4110 2387
rect 385 2377 486 2382
rect 1121 2377 1126 2382
rect 1569 2377 1574 2382
rect 1857 2377 1862 2382
rect 2929 2377 2934 2382
rect 65 2372 110 2377
rect 361 2372 390 2377
rect 481 2372 518 2377
rect 529 2372 598 2377
rect 617 2372 718 2377
rect 825 2372 1070 2377
rect 1121 2372 1574 2377
rect 1585 2372 1630 2377
rect 1649 2372 1718 2377
rect 1745 2372 1862 2377
rect 1881 2372 1910 2377
rect 1921 2372 1974 2377
rect 2041 2372 2126 2377
rect 2137 2372 2390 2377
rect 2457 2372 2870 2377
rect 2929 2372 3038 2377
rect 3057 2372 3102 2377
rect 3129 2372 3270 2377
rect 3353 2372 4222 2377
rect 1585 2367 1590 2372
rect 1713 2367 1718 2372
rect 73 2362 118 2367
rect 209 2362 254 2367
rect 345 2362 806 2367
rect 897 2362 990 2367
rect 1105 2362 1150 2367
rect 1241 2362 1262 2367
rect 1369 2362 1390 2367
rect 1409 2362 1462 2367
rect 1513 2362 1590 2367
rect 1609 2362 1670 2367
rect 1713 2362 2110 2367
rect 2177 2362 2262 2367
rect 2281 2362 2910 2367
rect 2945 2362 4054 2367
rect 4097 2362 4374 2367
rect 137 2352 206 2357
rect 305 2352 366 2357
rect 385 2352 510 2357
rect 537 2352 1718 2357
rect 1729 2352 1774 2357
rect 1825 2352 1878 2357
rect 1921 2352 2014 2357
rect 2057 2352 2190 2357
rect 2313 2352 2670 2357
rect 2681 2352 3134 2357
rect 3177 2352 3790 2357
rect 3897 2352 3958 2357
rect 4073 2352 4118 2357
rect 4145 2352 4310 2357
rect 193 2342 382 2347
rect 401 2342 430 2347
rect 553 2342 598 2347
rect 641 2342 702 2347
rect 737 2342 830 2347
rect 969 2342 1022 2347
rect 1057 2342 1270 2347
rect 1305 2342 1406 2347
rect 1417 2342 1502 2347
rect 1513 2342 1558 2347
rect 1569 2342 1630 2347
rect 1721 2342 1942 2347
rect 2089 2342 2166 2347
rect 2225 2342 2326 2347
rect 2409 2342 2486 2347
rect 2513 2342 2550 2347
rect 2569 2342 2606 2347
rect 2665 2342 2694 2347
rect 2849 2342 3222 2347
rect 3233 2342 3358 2347
rect 3377 2342 3438 2347
rect 3521 2342 3566 2347
rect 3625 2342 3702 2347
rect 3777 2342 3822 2347
rect 3937 2342 4006 2347
rect 4233 2342 4318 2347
rect 2689 2337 2854 2342
rect 169 2332 222 2337
rect 369 2332 454 2337
rect 673 2332 798 2337
rect 673 2327 678 2332
rect 793 2327 798 2332
rect 921 2332 2238 2337
rect 2249 2332 2662 2337
rect 2873 2332 2918 2337
rect 2929 2332 3110 2337
rect 3177 2332 3198 2337
rect 3257 2332 3390 2337
rect 3409 2332 4094 2337
rect 4161 2332 4278 2337
rect 921 2327 926 2332
rect 2929 2327 2934 2332
rect 3409 2327 3414 2332
rect 553 2322 678 2327
rect 361 2317 494 2322
rect 769 2317 774 2327
rect 793 2322 926 2327
rect 945 2322 974 2327
rect 337 2312 366 2317
rect 489 2312 614 2317
rect 737 2312 774 2317
rect 969 2317 974 2322
rect 1073 2322 2534 2327
rect 2713 2322 2758 2327
rect 2785 2322 2934 2327
rect 2953 2322 2998 2327
rect 3009 2322 3414 2327
rect 3561 2322 3822 2327
rect 4065 2322 4150 2327
rect 4329 2322 4358 2327
rect 1073 2317 1078 2322
rect 2585 2317 2694 2322
rect 3433 2317 3542 2322
rect 3913 2317 4038 2322
rect 4145 2317 4230 2322
rect 4329 2317 4334 2322
rect 969 2312 1078 2317
rect 1097 2312 1382 2317
rect 1393 2312 1430 2317
rect 1497 2312 1654 2317
rect 1689 2312 1726 2317
rect 1793 2312 2590 2317
rect 2689 2312 3438 2317
rect 3537 2312 3790 2317
rect 3801 2312 3918 2317
rect 4033 2312 4062 2317
rect 4225 2312 4334 2317
rect 1393 2307 1398 2312
rect 161 2302 198 2307
rect 233 2302 478 2307
rect 561 2302 662 2307
rect 1105 2302 1182 2307
rect 1201 2302 1326 2307
rect 1361 2302 1398 2307
rect 1409 2302 1510 2307
rect 1537 2302 1774 2307
rect 1785 2302 1846 2307
rect 1857 2302 2126 2307
rect 2185 2302 2206 2307
rect 2281 2302 2342 2307
rect 2409 2302 2478 2307
rect 2601 2302 4142 2307
rect 153 2292 214 2297
rect 321 2292 398 2297
rect 705 2292 750 2297
rect 1153 2292 1318 2297
rect 1337 2292 1998 2297
rect 2081 2292 2150 2297
rect 2161 2292 2238 2297
rect 2273 2292 2902 2297
rect 2913 2292 3054 2297
rect 3065 2292 3534 2297
rect 4105 2292 4206 2297
rect 521 2287 630 2292
rect 1313 2287 1318 2292
rect 1993 2287 2086 2292
rect 153 2282 310 2287
rect 409 2282 526 2287
rect 625 2282 654 2287
rect 665 2282 822 2287
rect 905 2282 1070 2287
rect 1089 2282 1206 2287
rect 1217 2282 1270 2287
rect 1313 2282 1734 2287
rect 1745 2282 1974 2287
rect 2137 2282 2230 2287
rect 305 2277 414 2282
rect 905 2277 910 2282
rect 537 2272 606 2277
rect 649 2272 718 2277
rect 737 2272 814 2277
rect 881 2272 910 2277
rect 1065 2277 1070 2282
rect 2273 2277 2278 2292
rect 3553 2287 3798 2292
rect 3969 2287 4086 2292
rect 2297 2282 2446 2287
rect 2473 2282 2646 2287
rect 2657 2282 2958 2287
rect 2985 2282 3558 2287
rect 3793 2282 3822 2287
rect 3905 2282 3974 2287
rect 4081 2282 4238 2287
rect 2657 2277 2662 2282
rect 3905 2277 3910 2282
rect 1065 2272 2278 2277
rect 2289 2272 2374 2277
rect 2425 2272 2662 2277
rect 2745 2272 2918 2277
rect 2977 2272 3030 2277
rect 3049 2272 3102 2277
rect 3145 2272 3198 2277
rect 3233 2272 3278 2277
rect 3385 2272 3910 2277
rect 3977 2272 4382 2277
rect 289 2262 414 2267
rect 433 2262 798 2267
rect 833 2262 1014 2267
rect 1177 2262 1230 2267
rect 1257 2262 1318 2267
rect 1337 2262 1398 2267
rect 1409 2262 1470 2267
rect 1481 2262 1862 2267
rect 1913 2262 2014 2267
rect 2209 2262 2246 2267
rect 2513 2262 2542 2267
rect 2561 2262 3350 2267
rect 3505 2262 3774 2267
rect 3849 2262 4214 2267
rect 289 2257 294 2262
rect 177 2252 294 2257
rect 409 2257 414 2262
rect 1089 2257 1158 2262
rect 2433 2257 2518 2262
rect 3369 2257 3470 2262
rect 409 2252 582 2257
rect 761 2252 854 2257
rect 977 2252 1094 2257
rect 1153 2252 2326 2257
rect 2337 2252 2406 2257
rect 577 2247 766 2252
rect 2433 2247 2438 2257
rect 2737 2252 2854 2257
rect 2897 2252 3070 2257
rect 3105 2252 3374 2257
rect 3465 2252 3958 2257
rect 4049 2252 4166 2257
rect 2545 2247 2718 2252
rect 2897 2247 2902 2252
rect 3953 2247 4054 2252
rect 0 2242 78 2247
rect 129 2242 166 2247
rect 161 2237 166 2242
rect 305 2242 558 2247
rect 785 2242 966 2247
rect 1105 2242 1286 2247
rect 1305 2242 1478 2247
rect 1537 2242 1574 2247
rect 1585 2242 1846 2247
rect 1857 2242 1878 2247
rect 2041 2242 2438 2247
rect 2521 2242 2550 2247
rect 2713 2242 2902 2247
rect 2913 2242 3238 2247
rect 3289 2242 3318 2247
rect 3337 2242 3406 2247
rect 3417 2242 3454 2247
rect 3537 2242 3750 2247
rect 3761 2242 3830 2247
rect 3873 2242 3934 2247
rect 4073 2242 4150 2247
rect 305 2237 310 2242
rect 1897 2237 1966 2242
rect 2913 2237 2918 2242
rect 3761 2237 3766 2242
rect 161 2232 310 2237
rect 345 2232 454 2237
rect 617 2232 670 2237
rect 681 2232 702 2237
rect 761 2232 830 2237
rect 953 2232 1902 2237
rect 1961 2232 2182 2237
rect 2241 2232 2598 2237
rect 2625 2232 2854 2237
rect 2889 2232 2918 2237
rect 2937 2232 3030 2237
rect 3113 2232 3478 2237
rect 3569 2232 3766 2237
rect 3777 2232 3830 2237
rect 3889 2232 4038 2237
rect 2241 2227 2246 2232
rect 4057 2227 4190 2232
rect 329 2222 350 2227
rect 521 2222 582 2227
rect 649 2222 678 2227
rect 721 2222 750 2227
rect 769 2222 798 2227
rect 825 2222 854 2227
rect 905 2222 1094 2227
rect 1121 2222 1190 2227
rect 1217 2222 1262 2227
rect 1345 2222 1366 2227
rect 1417 2222 1454 2227
rect 1473 2222 1814 2227
rect 1881 2222 1950 2227
rect 2033 2222 2078 2227
rect 2089 2222 2246 2227
rect 2281 2222 2406 2227
rect 2537 2222 2638 2227
rect 2649 2222 2950 2227
rect 2961 2222 3102 2227
rect 3121 2222 3222 2227
rect 3233 2222 3318 2227
rect 3329 2222 3534 2227
rect 3593 2222 3870 2227
rect 4025 2222 4062 2227
rect 4185 2222 4214 2227
rect 1809 2217 1814 2222
rect 2033 2217 2038 2222
rect 2961 2217 2966 2222
rect 369 2212 454 2217
rect 681 2212 1766 2217
rect 1809 2212 1974 2217
rect 1985 2212 2038 2217
rect 2209 2212 2302 2217
rect 2809 2212 2862 2217
rect 2913 2212 2966 2217
rect 3001 2212 3454 2217
rect 3537 2212 4286 2217
rect 369 2207 374 2212
rect 305 2202 374 2207
rect 449 2207 454 2212
rect 3449 2207 3542 2212
rect 449 2202 894 2207
rect 905 2202 934 2207
rect 1009 2202 1046 2207
rect 1057 2202 1230 2207
rect 1241 2202 1998 2207
rect 2073 2202 2382 2207
rect 2409 2202 2566 2207
rect 2753 2202 2910 2207
rect 2929 2202 3134 2207
rect 3145 2202 3262 2207
rect 3297 2202 3374 2207
rect 3393 2202 3430 2207
rect 2377 2197 2382 2202
rect 2929 2197 2934 2202
rect 3425 2197 3430 2202
rect 3561 2202 3686 2207
rect 361 2192 438 2197
rect 585 2192 622 2197
rect 641 2192 750 2197
rect 793 2192 1382 2197
rect 1393 2192 2022 2197
rect 2033 2192 2134 2197
rect 2377 2192 2406 2197
rect 2609 2192 2654 2197
rect 2721 2192 2798 2197
rect 2825 2192 2934 2197
rect 2953 2192 3198 2197
rect 3209 2192 3342 2197
rect 3353 2192 3406 2197
rect 3425 2192 3462 2197
rect 3561 2192 3566 2202
rect 3681 2197 3686 2202
rect 3745 2202 3854 2207
rect 3865 2202 3982 2207
rect 3745 2197 3750 2202
rect 3585 2192 3670 2197
rect 3681 2192 3750 2197
rect 3761 2192 3902 2197
rect 3985 2192 4054 2197
rect 4065 2192 4110 2197
rect 4257 2192 4374 2197
rect 257 2182 294 2187
rect 305 2182 446 2187
rect 561 2182 598 2187
rect 305 2177 310 2182
rect 641 2177 646 2192
rect 1377 2187 1382 2192
rect 2153 2187 2286 2192
rect 2473 2187 2590 2192
rect 737 2182 838 2187
rect 873 2182 958 2187
rect 1025 2182 1102 2187
rect 1145 2182 1174 2187
rect 1185 2182 1238 2187
rect 1249 2182 1270 2187
rect 1289 2182 1326 2187
rect 1337 2182 1366 2187
rect 1377 2182 1510 2187
rect 1521 2182 1558 2187
rect 1577 2182 1630 2187
rect 1665 2182 1734 2187
rect 1761 2182 1790 2187
rect 1865 2182 1942 2187
rect 1953 2182 2006 2187
rect 2025 2182 2158 2187
rect 2281 2182 2478 2187
rect 2585 2182 2710 2187
rect 2873 2182 4102 2187
rect 2049 2177 2054 2182
rect 2705 2177 2878 2182
rect 201 2172 310 2177
rect 329 2172 358 2177
rect 489 2172 646 2177
rect 673 2172 838 2177
rect 889 2172 2054 2177
rect 2089 2172 2222 2177
rect 2281 2172 2310 2177
rect 2337 2172 2358 2177
rect 2489 2172 2678 2177
rect 2897 2172 2942 2177
rect 2961 2172 3102 2177
rect 3137 2172 3190 2177
rect 3249 2172 3278 2177
rect 3297 2172 3326 2177
rect 3337 2172 3566 2177
rect 3585 2172 3726 2177
rect 3833 2172 3974 2177
rect 4089 2172 4238 2177
rect 353 2167 358 2172
rect 2961 2167 2966 2172
rect 3249 2167 3254 2172
rect 209 2162 326 2167
rect 353 2162 382 2167
rect 569 2162 630 2167
rect 705 2162 790 2167
rect 857 2162 950 2167
rect 977 2162 1006 2167
rect 1105 2162 1126 2167
rect 1137 2162 1230 2167
rect 1241 2162 1470 2167
rect 1513 2162 1630 2167
rect 1689 2162 1718 2167
rect 1729 2162 1750 2167
rect 1833 2162 2454 2167
rect 2513 2162 2734 2167
rect 2777 2162 2966 2167
rect 2985 2162 3254 2167
rect 3265 2162 3622 2167
rect 3817 2162 3870 2167
rect 3961 2162 3998 2167
rect 321 2152 326 2162
rect 705 2157 710 2162
rect 4017 2157 4238 2162
rect 353 2152 406 2157
rect 505 2152 550 2157
rect 585 2152 710 2157
rect 721 2152 862 2157
rect 921 2152 1006 2157
rect 1081 2152 1134 2157
rect 1145 2152 1246 2157
rect 1281 2152 2422 2157
rect 2569 2152 3254 2157
rect 3313 2152 3406 2157
rect 3433 2152 3606 2157
rect 3641 2152 4022 2157
rect 4233 2152 4294 2157
rect 721 2147 726 2152
rect 2417 2147 2574 2152
rect 193 2142 238 2147
rect 497 2142 726 2147
rect 737 2142 1582 2147
rect 1665 2142 1734 2147
rect 1769 2142 1790 2147
rect 1801 2142 1894 2147
rect 2001 2142 2174 2147
rect 2193 2142 2302 2147
rect 2337 2142 2398 2147
rect 2609 2142 2662 2147
rect 2681 2142 2718 2147
rect 2785 2142 2862 2147
rect 2929 2142 3150 2147
rect 3201 2142 3262 2147
rect 3345 2142 3702 2147
rect 3761 2142 3806 2147
rect 3993 2142 4022 2147
rect 4033 2142 4222 2147
rect 4313 2142 4342 2147
rect 2337 2137 2342 2142
rect 169 2132 486 2137
rect 577 2132 1022 2137
rect 1041 2132 2014 2137
rect 2113 2132 2342 2137
rect 2393 2137 2398 2142
rect 2657 2137 2662 2142
rect 4033 2137 4038 2142
rect 4217 2137 4318 2142
rect 2393 2132 2598 2137
rect 2657 2132 2958 2137
rect 2977 2132 3094 2137
rect 3105 2132 3158 2137
rect 3193 2132 3214 2137
rect 3273 2132 3334 2137
rect 3449 2132 3934 2137
rect 3961 2132 4038 2137
rect 481 2127 582 2132
rect 2009 2127 2118 2132
rect 2593 2127 2598 2132
rect 3329 2127 3454 2132
rect 4121 2127 4198 2132
rect 73 2122 294 2127
rect 601 2122 806 2127
rect 833 2122 1046 2127
rect 1057 2122 1254 2127
rect 1265 2122 1398 2127
rect 1449 2122 1526 2127
rect 1617 2122 1678 2127
rect 1761 2122 1830 2127
rect 1849 2122 1870 2127
rect 1945 2122 1990 2127
rect 2137 2122 2286 2127
rect 2593 2122 3302 2127
rect 3473 2122 3510 2127
rect 3561 2122 3846 2127
rect 3905 2122 4030 2127
rect 4041 2122 4126 2127
rect 4193 2122 4262 2127
rect 3905 2117 3910 2122
rect 137 2112 222 2117
rect 241 2112 486 2117
rect 529 2112 590 2117
rect 649 2112 742 2117
rect 761 2112 806 2117
rect 905 2112 2062 2117
rect 2097 2112 2166 2117
rect 2193 2112 2246 2117
rect 2305 2112 2422 2117
rect 2441 2112 2534 2117
rect 2569 2112 2990 2117
rect 3001 2112 3086 2117
rect 3193 2112 3270 2117
rect 3321 2112 3390 2117
rect 3425 2112 3798 2117
rect 3849 2112 3910 2117
rect 3921 2112 3982 2117
rect 4097 2112 4182 2117
rect 2305 2107 2310 2112
rect 169 2102 206 2107
rect 441 2102 558 2107
rect 593 2102 694 2107
rect 793 2102 846 2107
rect 857 2102 998 2107
rect 1017 2102 1214 2107
rect 1281 2102 1310 2107
rect 1345 2102 1382 2107
rect 1393 2102 1470 2107
rect 1593 2102 1910 2107
rect 2081 2102 2310 2107
rect 2417 2107 2422 2112
rect 4209 2107 4302 2112
rect 2417 2102 2510 2107
rect 2625 2102 3142 2107
rect 3153 2102 3566 2107
rect 3745 2102 3790 2107
rect 3817 2102 4166 2107
rect 4185 2102 4214 2107
rect 4297 2102 4326 2107
rect 993 2097 998 2102
rect 1905 2097 2086 2102
rect 2505 2097 2630 2102
rect 3153 2097 3158 2102
rect 3585 2097 3726 2102
rect 4161 2097 4166 2102
rect 313 2092 430 2097
rect 489 2092 694 2097
rect 721 2092 798 2097
rect 809 2092 974 2097
rect 993 2092 1886 2097
rect 2105 2092 2238 2097
rect 2265 2092 2486 2097
rect 2649 2092 2702 2097
rect 2761 2092 2854 2097
rect 2969 2092 2998 2097
rect 3057 2092 3158 2097
rect 3169 2092 3590 2097
rect 3721 2092 3806 2097
rect 3929 2092 4150 2097
rect 4161 2092 4278 2097
rect 425 2087 494 2092
rect 513 2082 598 2087
rect 681 2082 726 2087
rect 769 2082 1438 2087
rect 1505 2082 1598 2087
rect 1833 2082 2006 2087
rect 2233 2082 2278 2087
rect 2297 2082 2350 2087
rect 2465 2082 2542 2087
rect 2593 2082 2830 2087
rect 2945 2082 3294 2087
rect 3305 2082 3454 2087
rect 3505 2082 3558 2087
rect 3609 2082 4046 2087
rect 4065 2082 4134 2087
rect 4241 2082 4270 2087
rect 1617 2077 1718 2082
rect 4129 2077 4246 2082
rect 337 2072 958 2077
rect 1049 2072 1078 2077
rect 1169 2072 1262 2077
rect 1281 2072 1326 2077
rect 1345 2072 1622 2077
rect 1713 2072 2574 2077
rect 2593 2072 2694 2077
rect 2705 2072 3342 2077
rect 3353 2072 3590 2077
rect 3609 2072 3950 2077
rect 2593 2067 2598 2072
rect 2705 2067 2710 2072
rect 3337 2067 3342 2072
rect 3969 2067 4078 2072
rect 449 2062 550 2067
rect 569 2062 662 2067
rect 713 2062 734 2067
rect 761 2062 822 2067
rect 841 2062 878 2067
rect 921 2062 950 2067
rect 961 2062 1038 2067
rect 1129 2062 1166 2067
rect 1177 2062 1334 2067
rect 1353 2062 1414 2067
rect 1521 2062 1550 2067
rect 1569 2062 1638 2067
rect 1649 2062 1678 2067
rect 1737 2062 1854 2067
rect 1913 2062 2014 2067
rect 2025 2062 2182 2067
rect 2273 2062 2502 2067
rect 2561 2062 2598 2067
rect 2617 2062 2662 2067
rect 2673 2062 2710 2067
rect 2729 2062 2758 2067
rect 2777 2062 3182 2067
rect 3225 2062 3326 2067
rect 3337 2062 3430 2067
rect 3441 2062 3974 2067
rect 4073 2062 4102 2067
rect 4145 2062 4286 2067
rect 1329 2057 1334 2062
rect 2657 2057 2662 2062
rect 3425 2057 3430 2062
rect 89 2052 134 2057
rect 201 2052 318 2057
rect 609 2052 630 2057
rect 649 2052 678 2057
rect 817 2052 886 2057
rect 945 2052 998 2057
rect 1105 2052 1206 2057
rect 1217 2052 1246 2057
rect 1289 2052 1318 2057
rect 1329 2052 1382 2057
rect 1529 2052 1566 2057
rect 1601 2052 1854 2057
rect 1889 2052 2110 2057
rect 2257 2052 2374 2057
rect 2449 2052 2486 2057
rect 2585 2052 2606 2057
rect 2657 2052 2702 2057
rect 2713 2052 3030 2057
rect 3089 2052 3334 2057
rect 3425 2052 3486 2057
rect 3497 2052 3534 2057
rect 3569 2052 4022 2057
rect 4049 2052 4326 2057
rect 201 2047 206 2052
rect 177 2042 206 2047
rect 313 2047 318 2052
rect 697 2047 790 2052
rect 1401 2047 1510 2052
rect 3329 2047 3334 2052
rect 4049 2047 4054 2052
rect 313 2042 702 2047
rect 785 2042 814 2047
rect 985 2042 1406 2047
rect 1505 2042 2382 2047
rect 2417 2042 2494 2047
rect 2513 2042 3318 2047
rect 3329 2042 3470 2047
rect 3497 2042 3590 2047
rect 3625 2042 3654 2047
rect 3673 2042 3838 2047
rect 3849 2042 3926 2047
rect 4001 2042 4054 2047
rect 4073 2042 4142 2047
rect 4193 2042 4390 2047
rect 833 2037 966 2042
rect 169 2032 206 2037
rect 249 2032 358 2037
rect 577 2032 838 2037
rect 961 2032 1038 2037
rect 1065 2032 1182 2037
rect 1241 2032 1606 2037
rect 1641 2032 1766 2037
rect 1793 2032 1830 2037
rect 1897 2032 2062 2037
rect 2177 2032 2270 2037
rect 2289 2032 2790 2037
rect 2801 2032 2894 2037
rect 2905 2032 3062 2037
rect 3073 2032 3102 2037
rect 3113 2032 3134 2037
rect 3145 2032 3174 2037
rect 3209 2032 3262 2037
rect 3393 2032 4374 2037
rect 577 2027 582 2032
rect 2801 2027 2806 2032
rect 193 2022 230 2027
rect 297 2022 366 2027
rect 457 2022 582 2027
rect 593 2022 686 2027
rect 785 2022 942 2027
rect 977 2022 1110 2027
rect 1233 2022 1342 2027
rect 1377 2022 1798 2027
rect 1841 2022 2014 2027
rect 2041 2022 2086 2027
rect 2193 2022 2270 2027
rect 2385 2022 2422 2027
rect 2505 2022 2534 2027
rect 2705 2022 2734 2027
rect 2753 2022 2806 2027
rect 2849 2022 3254 2027
rect 3281 2022 3374 2027
rect 3561 2022 3670 2027
rect 3705 2022 3734 2027
rect 3793 2022 3870 2027
rect 4009 2022 4198 2027
rect 4209 2022 4238 2027
rect 2529 2017 2710 2022
rect 3281 2017 3286 2022
rect 3369 2017 3526 2022
rect 3793 2017 3798 2022
rect 393 2012 678 2017
rect 105 2002 206 2007
rect 433 2002 502 2007
rect 577 2002 670 2007
rect 497 1992 574 1997
rect 769 1992 790 1997
rect 801 1992 806 2017
rect 929 2012 950 2017
rect 993 2012 1022 2017
rect 1121 2012 2430 2017
rect 2785 2012 3286 2017
rect 3521 2012 3646 2017
rect 3657 2012 3694 2017
rect 3705 2012 3798 2017
rect 3841 2012 3862 2017
rect 3897 2012 4086 2017
rect 4145 2012 4198 2017
rect 825 2002 902 2007
rect 897 1997 902 2002
rect 857 1992 886 1997
rect 897 1992 934 1997
rect 945 1992 950 2012
rect 1017 2007 1126 2012
rect 1153 2002 1270 2007
rect 1289 2002 1350 2007
rect 1473 2002 2198 2007
rect 2217 2002 2558 2007
rect 2577 2002 2598 2007
rect 2649 2002 2774 2007
rect 2873 2002 3502 2007
rect 3593 2002 3782 2007
rect 1153 1997 1158 2002
rect 2769 1997 2878 2002
rect 3497 1997 3598 2002
rect 3841 1997 3846 2012
rect 3865 2002 4038 2007
rect 4137 2002 4270 2007
rect 1009 1992 1094 1997
rect 1105 1992 1158 1997
rect 1177 1992 1422 1997
rect 1441 1992 2710 1997
rect 2897 1992 2990 1997
rect 3033 1992 3142 1997
rect 3169 1992 3222 1997
rect 3313 1992 3478 1997
rect 3617 1992 3710 1997
rect 3737 1992 3806 1997
rect 3841 1992 3862 1997
rect 3913 1992 4054 1997
rect 4081 1992 4174 1997
rect 4257 1992 4310 1997
rect 4321 1992 4326 2032
rect 4385 2027 4390 2042
rect 4369 2022 4390 2027
rect 593 1987 750 1992
rect 4257 1987 4262 1992
rect 385 1982 598 1987
rect 745 1982 830 1987
rect 865 1982 918 1987
rect 937 1982 982 1987
rect 1089 1982 2030 1987
rect 2081 1982 2206 1987
rect 2257 1982 2286 1987
rect 2345 1982 2414 1987
rect 2561 1982 2766 1987
rect 2841 1982 2982 1987
rect 3009 1982 3510 1987
rect 3521 1982 3686 1987
rect 3729 1982 3966 1987
rect 3977 1982 4262 1987
rect 4281 1982 4326 1987
rect 2449 1977 2566 1982
rect 193 1972 406 1977
rect 473 1972 1102 1977
rect 1121 1972 1206 1977
rect 1249 1972 1318 1977
rect 1329 1972 1390 1977
rect 1417 1972 1558 1977
rect 1577 1972 1598 1977
rect 1609 1972 1702 1977
rect 1329 1967 1334 1972
rect 1553 1967 1558 1972
rect 1729 1967 1734 1977
rect 1745 1972 1830 1977
rect 1881 1972 2110 1977
rect 2225 1972 2318 1977
rect 2329 1972 2366 1977
rect 2385 1972 2454 1977
rect 2577 1972 3782 1977
rect 3801 1972 4038 1977
rect 4153 1972 4222 1977
rect 2225 1967 2230 1972
rect 4033 1967 4158 1972
rect 513 1962 590 1967
rect 801 1962 878 1967
rect 969 1962 998 1967
rect 1129 1962 1302 1967
rect 1313 1962 1334 1967
rect 1417 1962 1438 1967
rect 1449 1962 1542 1967
rect 1553 1962 1662 1967
rect 1729 1962 1774 1967
rect 2169 1962 2230 1967
rect 2241 1962 2750 1967
rect 2785 1962 2854 1967
rect 2921 1962 2974 1967
rect 2985 1962 3246 1967
rect 3481 1962 3662 1967
rect 3673 1962 3734 1967
rect 3785 1962 3830 1967
rect 3873 1962 3950 1967
rect 3969 1962 4014 1967
rect 4217 1962 4254 1967
rect 329 1957 494 1962
rect 633 1957 750 1962
rect 993 1957 1134 1962
rect 3265 1957 3366 1962
rect 177 1952 334 1957
rect 489 1952 638 1957
rect 745 1952 774 1957
rect 833 1952 854 1957
rect 1153 1952 1174 1957
rect 1265 1952 1798 1957
rect 1809 1952 1910 1957
rect 1953 1952 1974 1957
rect 1993 1952 2070 1957
rect 2321 1952 2494 1957
rect 2505 1952 2582 1957
rect 2593 1952 2678 1957
rect 2705 1952 2750 1957
rect 2777 1952 3270 1957
rect 3361 1952 3390 1957
rect 3465 1952 3534 1957
rect 3593 1952 4142 1957
rect 4193 1952 4262 1957
rect 1265 1947 1270 1952
rect 1953 1947 1958 1952
rect 345 1942 470 1947
rect 529 1937 534 1947
rect 649 1942 910 1947
rect 1041 1942 1078 1947
rect 1177 1942 1270 1947
rect 1289 1942 1534 1947
rect 1545 1942 1574 1947
rect 1585 1937 1590 1947
rect 1609 1942 1654 1947
rect 1665 1942 1686 1947
rect 1721 1942 1790 1947
rect 1849 1942 1958 1947
rect 1977 1942 2014 1947
rect 2089 1942 2230 1947
rect 2249 1942 2366 1947
rect 2409 1942 2470 1947
rect 2513 1942 3070 1947
rect 3081 1942 3158 1947
rect 3193 1942 3638 1947
rect 3721 1942 3758 1947
rect 3825 1942 3942 1947
rect 3985 1942 4206 1947
rect 2089 1937 2094 1942
rect 489 1932 1510 1937
rect 1529 1932 1590 1937
rect 1641 1932 2094 1937
rect 2225 1937 2230 1942
rect 2225 1932 3222 1937
rect 3249 1932 3414 1937
rect 3425 1932 3462 1937
rect 3489 1932 3526 1937
rect 3593 1932 3798 1937
rect 3833 1932 3974 1937
rect 2129 1927 2206 1932
rect 3425 1927 3430 1932
rect 3985 1927 3990 1942
rect 4065 1932 4238 1937
rect 4065 1927 4070 1932
rect 4257 1927 4262 1952
rect 217 1922 350 1927
rect 345 1917 350 1922
rect 505 1922 534 1927
rect 665 1922 942 1927
rect 1153 1922 1718 1927
rect 1745 1922 1854 1927
rect 1873 1922 1934 1927
rect 1953 1922 1998 1927
rect 2009 1922 2134 1927
rect 2201 1922 2286 1927
rect 2465 1922 2518 1927
rect 2577 1922 2622 1927
rect 2697 1922 2894 1927
rect 2945 1922 3022 1927
rect 3041 1922 3070 1927
rect 3089 1922 3142 1927
rect 3185 1922 3430 1927
rect 3441 1922 3590 1927
rect 3673 1922 3830 1927
rect 3897 1922 3926 1927
rect 3937 1922 3990 1927
rect 4025 1922 4070 1927
rect 4089 1922 4158 1927
rect 4209 1922 4262 1927
rect 4337 1922 4382 1927
rect 505 1917 510 1922
rect 961 1917 1134 1922
rect 345 1912 510 1917
rect 553 1912 966 1917
rect 1129 1912 1454 1917
rect 1489 1912 1494 1922
rect 1873 1917 1878 1922
rect 2313 1917 2446 1922
rect 3137 1917 3142 1922
rect 1513 1912 1550 1917
rect 1561 1912 1710 1917
rect 1729 1912 1774 1917
rect 1833 1912 1878 1917
rect 1905 1912 1974 1917
rect 1985 1912 2030 1917
rect 2145 1912 2206 1917
rect 2289 1912 2318 1917
rect 2441 1912 3126 1917
rect 3137 1912 3958 1917
rect 3969 1912 4142 1917
rect 3121 1907 3126 1912
rect 3969 1907 3974 1912
rect 617 1902 670 1907
rect 705 1902 742 1907
rect 889 1902 1102 1907
rect 1153 1902 1190 1907
rect 1209 1902 2334 1907
rect 2393 1902 2510 1907
rect 2633 1902 2718 1907
rect 2849 1902 3046 1907
rect 3065 1902 3110 1907
rect 3121 1902 3150 1907
rect 3209 1902 3270 1907
rect 3321 1902 3974 1907
rect 4137 1907 4142 1912
rect 4209 1907 4214 1922
rect 4225 1912 4318 1917
rect 4337 1907 4342 1922
rect 4137 1902 4214 1907
rect 4313 1902 4342 1907
rect 761 1897 870 1902
rect 2737 1897 2830 1902
rect 577 1892 622 1897
rect 689 1892 766 1897
rect 865 1892 1814 1897
rect 1865 1892 1926 1897
rect 2009 1892 2222 1897
rect 2305 1892 2742 1897
rect 2825 1892 3158 1897
rect 3177 1892 3606 1897
rect 3625 1892 3734 1897
rect 3745 1892 3822 1897
rect 3833 1892 3854 1897
rect 3865 1892 4078 1897
rect 4265 1892 4382 1897
rect 449 1882 766 1887
rect 817 1882 910 1887
rect 921 1882 990 1887
rect 1081 1882 1646 1887
rect 1657 1882 2438 1887
rect 2465 1882 3222 1887
rect 3321 1882 3382 1887
rect 3497 1882 3534 1887
rect 3577 1882 3630 1887
rect 3689 1882 3734 1887
rect 3745 1882 3974 1887
rect 4097 1882 4246 1887
rect 4265 1882 4374 1887
rect 3217 1877 3326 1882
rect 3993 1877 4102 1882
rect 4241 1877 4246 1882
rect 281 1872 438 1877
rect 521 1872 894 1877
rect 1025 1872 1126 1877
rect 1169 1872 2014 1877
rect 2121 1872 2406 1877
rect 2537 1872 2574 1877
rect 2665 1872 2734 1877
rect 2801 1872 2982 1877
rect 3081 1872 3110 1877
rect 3121 1872 3198 1877
rect 3345 1872 3366 1877
rect 3473 1872 3502 1877
rect 3593 1872 3998 1877
rect 4241 1872 4302 1877
rect 433 1867 526 1872
rect 1121 1867 1126 1872
rect 2009 1867 2126 1872
rect 2425 1867 2518 1872
rect 3497 1867 3598 1872
rect 4121 1867 4222 1872
rect 4297 1867 4302 1872
rect 4393 1872 4446 1877
rect 4393 1867 4398 1872
rect 545 1862 750 1867
rect 809 1862 990 1867
rect 1009 1862 1110 1867
rect 1121 1862 1206 1867
rect 1233 1862 1990 1867
rect 2145 1862 2254 1867
rect 2281 1862 2358 1867
rect 2369 1862 2430 1867
rect 2513 1862 2758 1867
rect 2809 1862 3246 1867
rect 3353 1862 3406 1867
rect 3617 1862 3670 1867
rect 3681 1862 4126 1867
rect 4217 1862 4246 1867
rect 4297 1862 4398 1867
rect 2145 1857 2150 1862
rect 497 1852 1638 1857
rect 1649 1852 1734 1857
rect 1793 1852 1846 1857
rect 1889 1852 2150 1857
rect 2169 1852 3190 1857
rect 3217 1852 3262 1857
rect 3281 1852 3310 1857
rect 3409 1852 3486 1857
rect 3529 1852 3622 1857
rect 3705 1852 3774 1857
rect 3785 1852 3870 1857
rect 3897 1852 4046 1857
rect 4073 1852 4262 1857
rect 377 1842 838 1847
rect 1009 1842 2030 1847
rect 2041 1842 2302 1847
rect 2353 1842 4062 1847
rect 4105 1842 4150 1847
rect 4177 1842 4278 1847
rect 857 1837 950 1842
rect 145 1832 190 1837
rect 241 1832 398 1837
rect 465 1832 862 1837
rect 945 1832 974 1837
rect 1073 1832 1398 1837
rect 1409 1832 1494 1837
rect 1505 1832 1582 1837
rect 1609 1832 1894 1837
rect 1921 1832 1958 1837
rect 2033 1832 2086 1837
rect 2161 1832 2182 1837
rect 2289 1832 3414 1837
rect 3521 1832 4062 1837
rect 4145 1832 4254 1837
rect 4345 1832 4406 1837
rect 2033 1827 2038 1832
rect 3409 1827 3526 1832
rect 169 1822 278 1827
rect 417 1822 510 1827
rect 657 1822 710 1827
rect 721 1822 830 1827
rect 865 1822 926 1827
rect 961 1822 982 1827
rect 993 1822 1030 1827
rect 1113 1822 1150 1827
rect 1161 1822 1190 1827
rect 1217 1822 1278 1827
rect 1313 1822 1350 1827
rect 1465 1822 1494 1827
rect 1585 1822 2038 1827
rect 2065 1822 2118 1827
rect 2129 1822 2206 1827
rect 2241 1822 2278 1827
rect 2305 1822 2622 1827
rect 2665 1822 2734 1827
rect 2745 1822 2790 1827
rect 2817 1822 2902 1827
rect 2969 1822 2998 1827
rect 3057 1822 3214 1827
rect 3265 1822 3310 1827
rect 3329 1822 3390 1827
rect 3545 1822 3654 1827
rect 3681 1822 4382 1827
rect 297 1817 398 1822
rect 505 1817 662 1822
rect 113 1812 302 1817
rect 393 1812 486 1817
rect 705 1807 710 1822
rect 961 1812 966 1822
rect 993 1807 998 1822
rect 1017 1812 1046 1817
rect 1057 1812 1078 1817
rect 1113 1812 2446 1817
rect 2561 1812 2966 1817
rect 3025 1812 3430 1817
rect 3569 1812 3838 1817
rect 3865 1812 4246 1817
rect 4257 1812 4358 1817
rect 137 1802 182 1807
rect 193 1802 222 1807
rect 257 1802 590 1807
rect 705 1802 998 1807
rect 1041 1807 1046 1812
rect 3569 1807 3574 1812
rect 4401 1807 4406 1832
rect 1041 1802 1182 1807
rect 1217 1802 1318 1807
rect 1401 1802 2454 1807
rect 2465 1802 2646 1807
rect 2681 1802 2790 1807
rect 2825 1802 3246 1807
rect 3393 1802 3438 1807
rect 3489 1802 3574 1807
rect 3593 1802 3686 1807
rect 3777 1802 3902 1807
rect 3937 1802 4054 1807
rect 4209 1802 4318 1807
rect 4353 1802 4406 1807
rect 193 1782 198 1802
rect 3265 1797 3334 1802
rect 4073 1797 4214 1802
rect 225 1792 438 1797
rect 729 1792 750 1797
rect 961 1792 1046 1797
rect 1081 1792 1166 1797
rect 1201 1792 1238 1797
rect 1257 1792 1326 1797
rect 1337 1792 1382 1797
rect 1393 1792 1454 1797
rect 1465 1792 1494 1797
rect 1521 1792 1638 1797
rect 1673 1792 2190 1797
rect 2305 1792 2334 1797
rect 2585 1792 2710 1797
rect 2721 1792 2750 1797
rect 2761 1792 2958 1797
rect 2977 1792 3086 1797
rect 3185 1792 3270 1797
rect 3329 1792 4078 1797
rect 4225 1792 4310 1797
rect 633 1787 710 1792
rect 2185 1787 2310 1792
rect 3105 1787 3190 1792
rect 433 1782 638 1787
rect 705 1782 854 1787
rect 1025 1782 2070 1787
rect 2089 1782 2166 1787
rect 2393 1782 2518 1787
rect 2537 1782 3110 1787
rect 3257 1782 3318 1787
rect 3393 1782 3750 1787
rect 3785 1782 3814 1787
rect 3929 1782 4006 1787
rect 4089 1782 4350 1787
rect 289 1777 438 1782
rect 897 1777 1006 1782
rect 2513 1777 2518 1782
rect 145 1772 190 1777
rect 265 1772 294 1777
rect 649 1772 766 1777
rect 873 1772 902 1777
rect 1001 1772 2062 1777
rect 2185 1772 2302 1777
rect 2321 1772 2462 1777
rect 2513 1772 3230 1777
rect 3289 1772 3894 1777
rect 3921 1772 3990 1777
rect 4017 1772 4118 1777
rect 4185 1772 4254 1777
rect 553 1767 654 1772
rect 2089 1767 2190 1772
rect 2297 1767 2302 1772
rect 3921 1767 3926 1772
rect 249 1762 558 1767
rect 673 1762 750 1767
rect 921 1762 1030 1767
rect 1073 1762 1438 1767
rect 1521 1762 1686 1767
rect 1705 1762 1750 1767
rect 1841 1762 2006 1767
rect 2065 1762 2094 1767
rect 2297 1762 2526 1767
rect 2633 1762 3014 1767
rect 3025 1762 3174 1767
rect 3265 1762 3310 1767
rect 3353 1762 3422 1767
rect 3465 1762 3806 1767
rect 3833 1762 3926 1767
rect 4041 1762 4262 1767
rect 3169 1757 3254 1762
rect 577 1752 686 1757
rect 761 1752 854 1757
rect 873 1752 926 1757
rect 937 1752 998 1757
rect 1041 1752 1494 1757
rect 1577 1752 1622 1757
rect 1641 1752 2166 1757
rect 2217 1752 2334 1757
rect 2345 1752 3150 1757
rect 3249 1752 3286 1757
rect 3385 1752 3462 1757
rect 3505 1752 3542 1757
rect 3617 1752 3870 1757
rect 3881 1752 3918 1757
rect 3993 1752 4086 1757
rect 4097 1752 4206 1757
rect 425 1747 558 1752
rect 681 1747 766 1752
rect 137 1742 222 1747
rect 337 1742 430 1747
rect 553 1742 662 1747
rect 913 1742 958 1747
rect 1017 1742 1270 1747
rect 1361 1742 1798 1747
rect 1809 1742 1974 1747
rect 1985 1742 2030 1747
rect 2049 1742 2246 1747
rect 2337 1742 2734 1747
rect 2745 1742 2830 1747
rect 2897 1742 2950 1747
rect 2961 1742 3238 1747
rect 3297 1742 3382 1747
rect 3553 1742 3750 1747
rect 3873 1742 3950 1747
rect 4113 1742 4190 1747
rect 1265 1737 1366 1742
rect 1809 1737 1814 1742
rect 161 1732 214 1737
rect 273 1732 326 1737
rect 321 1727 326 1732
rect 441 1732 1246 1737
rect 1385 1732 1462 1737
rect 1545 1732 1814 1737
rect 1857 1732 1926 1737
rect 1937 1732 2014 1737
rect 441 1727 446 1732
rect 2049 1727 2054 1742
rect 2961 1737 2966 1742
rect 3233 1737 3302 1742
rect 2137 1732 2182 1737
rect 2313 1732 2342 1737
rect 2465 1732 2590 1737
rect 2617 1732 2726 1737
rect 2865 1732 2966 1737
rect 2977 1732 3030 1737
rect 3041 1732 3110 1737
rect 3121 1732 3182 1737
rect 3457 1732 3814 1737
rect 4369 1732 4390 1737
rect 321 1722 446 1727
rect 497 1722 710 1727
rect 721 1722 902 1727
rect 929 1722 1590 1727
rect 1833 1722 1926 1727
rect 1953 1722 2054 1727
rect 2073 1722 2494 1727
rect 2793 1722 2822 1727
rect 2873 1722 3006 1727
rect 3089 1722 3206 1727
rect 3217 1722 3246 1727
rect 3265 1722 3438 1727
rect 3569 1722 3782 1727
rect 3857 1722 4022 1727
rect 4129 1722 4238 1727
rect 1657 1717 1790 1722
rect 2513 1717 2718 1722
rect 3265 1717 3270 1722
rect 201 1712 270 1717
rect 465 1712 526 1717
rect 593 1712 1662 1717
rect 1785 1712 1982 1717
rect 2145 1712 2166 1717
rect 2385 1712 2414 1717
rect 2425 1712 2518 1717
rect 2713 1712 3270 1717
rect 3433 1717 3438 1722
rect 3857 1717 3862 1722
rect 4017 1717 4022 1722
rect 4385 1717 4390 1732
rect 3433 1712 3518 1717
rect 3569 1712 3606 1717
rect 3633 1712 3670 1717
rect 3705 1712 3862 1717
rect 3881 1712 3974 1717
rect 4017 1712 4046 1717
rect 4105 1712 4142 1717
rect 4361 1712 4390 1717
rect 2001 1707 2118 1712
rect 2161 1707 2366 1712
rect 529 1702 630 1707
rect 665 1702 790 1707
rect 913 1702 1198 1707
rect 1241 1702 1318 1707
rect 1361 1702 1526 1707
rect 1569 1702 1606 1707
rect 1673 1702 1774 1707
rect 1841 1702 2006 1707
rect 2113 1702 2142 1707
rect 2361 1702 2702 1707
rect 2865 1702 2910 1707
rect 2929 1702 2958 1707
rect 3041 1702 3070 1707
rect 3081 1702 3142 1707
rect 3169 1702 3358 1707
rect 3369 1702 3590 1707
rect 3601 1702 3686 1707
rect 3745 1702 3806 1707
rect 3897 1702 3950 1707
rect 3977 1702 4238 1707
rect 2721 1697 2846 1702
rect 2953 1697 3046 1702
rect 3169 1697 3174 1702
rect 657 1692 1022 1697
rect 1281 1692 1302 1697
rect 1329 1692 2478 1697
rect 2537 1692 2574 1697
rect 2601 1692 2726 1697
rect 2841 1692 2886 1697
rect 3089 1692 3174 1697
rect 3185 1692 4158 1697
rect 4265 1692 4294 1697
rect 1081 1687 1262 1692
rect 4153 1687 4270 1692
rect 521 1682 646 1687
rect 1057 1682 1086 1687
rect 1257 1682 2422 1687
rect 2521 1682 2638 1687
rect 2649 1682 2926 1687
rect 2993 1682 3734 1687
rect 3761 1682 3782 1687
rect 3793 1682 4070 1687
rect 665 1677 758 1682
rect 809 1677 1038 1682
rect 289 1672 510 1677
rect 505 1667 510 1672
rect 601 1672 670 1677
rect 753 1672 814 1677
rect 1033 1672 2014 1677
rect 2033 1672 2102 1677
rect 2153 1672 2182 1677
rect 2273 1672 2350 1677
rect 2433 1672 2590 1677
rect 2753 1672 4286 1677
rect 601 1667 606 1672
rect 2345 1667 2438 1672
rect 2585 1667 2758 1672
rect 505 1662 606 1667
rect 625 1662 742 1667
rect 825 1662 1582 1667
rect 1593 1662 1670 1667
rect 1681 1662 1710 1667
rect 1801 1662 2046 1667
rect 2161 1662 2326 1667
rect 2489 1662 2566 1667
rect 2777 1662 2830 1667
rect 2905 1662 3150 1667
rect 3169 1662 3278 1667
rect 3313 1662 4014 1667
rect 4217 1662 4358 1667
rect 1665 1657 1670 1662
rect 2161 1657 2166 1662
rect 4009 1657 4014 1662
rect 4113 1657 4222 1662
rect 865 1652 926 1657
rect 1009 1652 1590 1657
rect 1617 1652 1654 1657
rect 1665 1652 1686 1657
rect 1769 1652 1854 1657
rect 2025 1652 2062 1657
rect 2081 1652 2166 1657
rect 2185 1652 2294 1657
rect 2361 1652 2414 1657
rect 2569 1652 2670 1657
rect 2833 1652 3422 1657
rect 3665 1652 3830 1657
rect 3945 1652 3990 1657
rect 4009 1652 4118 1657
rect 705 1647 814 1652
rect 1873 1647 2006 1652
rect 2081 1647 2086 1652
rect 2433 1647 2550 1652
rect 2833 1647 2838 1652
rect 3441 1647 3614 1652
rect 249 1642 374 1647
rect 249 1637 254 1642
rect 225 1632 254 1637
rect 369 1637 374 1642
rect 681 1642 710 1647
rect 809 1642 838 1647
rect 681 1637 686 1642
rect 369 1632 686 1637
rect 833 1637 838 1642
rect 881 1642 1126 1647
rect 1137 1642 1198 1647
rect 1209 1642 1406 1647
rect 1457 1642 1878 1647
rect 2001 1642 2086 1647
rect 2225 1642 2438 1647
rect 2545 1642 2590 1647
rect 2681 1642 2838 1647
rect 2857 1642 2998 1647
rect 3089 1642 3446 1647
rect 3609 1642 3702 1647
rect 3737 1642 3790 1647
rect 3801 1642 3846 1647
rect 4137 1642 4222 1647
rect 881 1637 886 1642
rect 2585 1637 2686 1642
rect 2993 1637 3094 1642
rect 3697 1637 3702 1642
rect 4137 1637 4142 1642
rect 833 1632 886 1637
rect 905 1632 958 1637
rect 993 1632 1086 1637
rect 1145 1632 1246 1637
rect 1289 1632 1646 1637
rect 1657 1632 2566 1637
rect 2713 1632 2974 1637
rect 3113 1632 3342 1637
rect 3425 1632 3518 1637
rect 3545 1632 3686 1637
rect 3697 1632 4142 1637
rect 4217 1637 4222 1642
rect 4217 1632 4246 1637
rect 4329 1632 4358 1637
rect 249 1622 358 1627
rect 689 1622 822 1627
rect 985 1622 1014 1627
rect 1009 1617 1014 1622
rect 1105 1622 1758 1627
rect 1785 1622 1862 1627
rect 1905 1622 2510 1627
rect 2529 1622 2726 1627
rect 2761 1622 3798 1627
rect 3817 1622 3902 1627
rect 4153 1622 4190 1627
rect 4225 1622 4334 1627
rect 1105 1617 1110 1622
rect 2529 1617 2534 1622
rect 4225 1617 4230 1622
rect 745 1612 774 1617
rect 769 1607 774 1612
rect 833 1612 982 1617
rect 1009 1612 1110 1617
rect 1169 1612 2310 1617
rect 2321 1612 2534 1617
rect 2545 1612 2662 1617
rect 2769 1612 2886 1617
rect 2929 1612 2990 1617
rect 3057 1612 3454 1617
rect 3561 1612 3638 1617
rect 3679 1612 3726 1617
rect 3737 1612 3830 1617
rect 833 1607 838 1612
rect 2305 1607 2310 1612
rect 2545 1607 2550 1612
rect 2657 1607 2758 1612
rect 417 1602 534 1607
rect 769 1602 838 1607
rect 1129 1602 1166 1607
rect 1217 1602 1286 1607
rect 1329 1602 1558 1607
rect 1569 1602 2278 1607
rect 2305 1602 2342 1607
rect 2417 1602 2550 1607
rect 2601 1602 2638 1607
rect 2753 1602 2942 1607
rect 2953 1602 3126 1607
rect 3137 1602 3206 1607
rect 3217 1602 3390 1607
rect 3497 1602 3574 1607
rect 3585 1602 3670 1607
rect 1553 1597 1558 1602
rect 2337 1597 2342 1602
rect 3679 1597 3684 1612
rect 3689 1602 3734 1607
rect 3769 1602 3814 1607
rect 3825 1602 3830 1612
rect 3953 1612 4030 1617
rect 4145 1612 4230 1617
rect 3953 1597 3958 1612
rect 4353 1607 4358 1632
rect 3969 1602 4094 1607
rect 4177 1602 4254 1607
rect 4329 1602 4358 1607
rect 137 1592 206 1597
rect 1129 1592 1486 1597
rect 1505 1592 1526 1597
rect 1553 1592 1982 1597
rect 2017 1592 2062 1597
rect 2097 1592 2206 1597
rect 2289 1592 2326 1597
rect 2337 1592 2358 1597
rect 2481 1592 3684 1597
rect 3721 1592 3742 1597
rect 3769 1592 3990 1597
rect 4017 1592 4078 1597
rect 4121 1592 4214 1597
rect 4297 1592 4326 1597
rect 689 1582 918 1587
rect 937 1582 1022 1587
rect 1145 1582 1926 1587
rect 1977 1582 2014 1587
rect 2033 1582 2110 1587
rect 2297 1582 2614 1587
rect 2633 1582 3214 1587
rect 3257 1582 3326 1587
rect 3385 1582 3486 1587
rect 3529 1582 3566 1587
rect 3585 1582 3646 1587
rect 3665 1582 3926 1587
rect 3961 1582 4118 1587
rect 689 1577 694 1582
rect 665 1572 694 1577
rect 913 1577 918 1582
rect 913 1572 942 1577
rect 1033 1572 1974 1577
rect 2017 1572 2310 1577
rect 2321 1572 2462 1577
rect 2513 1572 3126 1577
rect 3153 1572 3414 1577
rect 3425 1572 3598 1577
rect 3617 1572 3686 1577
rect 3697 1572 3726 1577
rect 3745 1572 3958 1577
rect 3977 1572 4302 1577
rect 777 1567 878 1572
rect 937 1567 1038 1572
rect 2305 1567 2310 1572
rect 3409 1567 3414 1572
rect 313 1562 374 1567
rect 625 1562 782 1567
rect 873 1562 902 1567
rect 1097 1562 1142 1567
rect 1153 1562 1326 1567
rect 1337 1562 1374 1567
rect 1385 1562 1430 1567
rect 1489 1562 1534 1567
rect 1577 1562 1702 1567
rect 1721 1562 1830 1567
rect 1953 1562 2054 1567
rect 2145 1562 2190 1567
rect 2305 1562 2678 1567
rect 2721 1562 2862 1567
rect 2881 1562 3174 1567
rect 3297 1562 3382 1567
rect 3409 1562 3542 1567
rect 3561 1562 3950 1567
rect 4001 1562 4150 1567
rect 209 1552 510 1557
rect 761 1552 886 1557
rect 897 1552 1022 1557
rect 1097 1552 1126 1557
rect 1217 1552 1342 1557
rect 1393 1552 1670 1557
rect 1769 1552 2406 1557
rect 2425 1552 2838 1557
rect 2889 1552 2966 1557
rect 2985 1552 3598 1557
rect 3633 1552 3798 1557
rect 4049 1552 4158 1557
rect 4217 1552 4310 1557
rect 881 1547 886 1552
rect 1665 1547 1774 1552
rect 2961 1547 2966 1552
rect 3817 1547 3894 1552
rect 3945 1547 4022 1552
rect 129 1542 302 1547
rect 329 1542 670 1547
rect 881 1542 1262 1547
rect 1481 1542 1646 1547
rect 1921 1542 2142 1547
rect 2177 1542 2222 1547
rect 721 1537 862 1542
rect 1257 1537 1350 1542
rect 1481 1537 1486 1542
rect 1793 1537 1926 1542
rect 2289 1537 2294 1547
rect 2401 1542 2446 1547
rect 2457 1542 2534 1547
rect 2593 1542 2918 1547
rect 2961 1542 3062 1547
rect 3089 1542 3142 1547
rect 3217 1542 3310 1547
rect 3353 1542 3822 1547
rect 3889 1542 3950 1547
rect 4017 1542 4094 1547
rect 2593 1537 2598 1542
rect 4081 1537 4102 1538
rect 201 1532 334 1537
rect 441 1532 470 1537
rect 649 1532 726 1537
rect 857 1532 1174 1537
rect 1209 1532 1238 1537
rect 1345 1532 1486 1537
rect 1505 1532 1662 1537
rect 1713 1532 1798 1537
rect 1945 1532 1982 1537
rect 1993 1532 2046 1537
rect 2145 1532 2214 1537
rect 2289 1532 2598 1537
rect 2617 1532 3750 1537
rect 3833 1532 3878 1537
rect 3961 1532 4070 1537
rect 4081 1533 4142 1537
rect 4097 1532 4142 1533
rect 329 1527 446 1532
rect 513 1522 638 1527
rect 129 1512 230 1517
rect 241 1512 502 1517
rect 513 1507 518 1522
rect 633 1517 638 1522
rect 737 1522 1326 1527
rect 1505 1522 1510 1532
rect 1545 1522 1670 1527
rect 1729 1522 1774 1527
rect 1873 1522 3342 1527
rect 3425 1522 3510 1527
rect 3537 1522 4070 1527
rect 4265 1522 4366 1527
rect 737 1517 742 1522
rect 4065 1517 4070 1522
rect 633 1512 742 1517
rect 761 1512 790 1517
rect 881 1512 934 1517
rect 993 1512 1022 1517
rect 1033 1512 1222 1517
rect 1257 1512 1318 1517
rect 1345 1512 1462 1517
rect 1481 1512 3046 1517
rect 3057 1512 3078 1517
rect 3097 1512 3134 1517
rect 3153 1512 3294 1517
rect 3329 1512 3430 1517
rect 3465 1512 3742 1517
rect 3817 1512 3894 1517
rect 3937 1512 4014 1517
rect 4065 1512 4166 1517
rect 4225 1512 4318 1517
rect 785 1507 886 1512
rect 1345 1507 1350 1512
rect 121 1502 150 1507
rect 145 1497 150 1502
rect 217 1502 518 1507
rect 905 1502 1350 1507
rect 1457 1507 1462 1512
rect 3073 1507 3078 1512
rect 1457 1502 2166 1507
rect 2201 1502 2342 1507
rect 2369 1502 3054 1507
rect 3073 1502 3110 1507
rect 3121 1502 3150 1507
rect 3209 1502 3326 1507
rect 3337 1502 3502 1507
rect 3521 1502 3694 1507
rect 3705 1502 3918 1507
rect 4025 1502 4198 1507
rect 4209 1502 4238 1507
rect 217 1497 222 1502
rect 73 1492 110 1497
rect 145 1492 222 1497
rect 529 1492 926 1497
rect 953 1492 998 1497
rect 1081 1492 1262 1497
rect 1281 1492 1742 1497
rect 1769 1492 2718 1497
rect 2801 1492 3078 1497
rect 3089 1492 3134 1497
rect 3169 1492 3222 1497
rect 3241 1492 3286 1497
rect 3297 1492 3406 1497
rect 3417 1492 3854 1497
rect 105 1477 110 1492
rect 529 1487 534 1492
rect 2713 1487 2806 1492
rect 3281 1487 3286 1492
rect 3849 1487 3854 1492
rect 3929 1492 4102 1497
rect 4249 1492 4278 1497
rect 3929 1487 3934 1492
rect 4097 1487 4254 1492
rect 281 1482 534 1487
rect 737 1482 766 1487
rect 1009 1482 1694 1487
rect 1737 1482 2118 1487
rect 2297 1482 2518 1487
rect 2545 1482 2630 1487
rect 2657 1482 2694 1487
rect 2945 1482 3270 1487
rect 3281 1482 3606 1487
rect 3617 1482 3638 1487
rect 3713 1482 3798 1487
rect 3849 1482 3934 1487
rect 3961 1482 4078 1487
rect 281 1477 286 1482
rect 761 1477 1014 1482
rect 2201 1477 2278 1482
rect 2825 1477 2926 1482
rect 3713 1477 3718 1482
rect 105 1472 286 1477
rect 1041 1472 1286 1477
rect 1513 1472 2206 1477
rect 2273 1472 2422 1477
rect 2433 1472 2614 1477
rect 2649 1472 2830 1477
rect 2921 1472 3718 1477
rect 3777 1472 3830 1477
rect 4041 1472 4206 1477
rect 1305 1467 1494 1472
rect 3825 1467 3830 1472
rect 313 1462 382 1467
rect 401 1462 702 1467
rect 721 1462 782 1467
rect 793 1462 1310 1467
rect 1489 1462 1926 1467
rect 2049 1462 2134 1467
rect 2217 1462 2558 1467
rect 2577 1462 2846 1467
rect 2865 1462 2934 1467
rect 2953 1462 3062 1467
rect 3097 1462 3118 1467
rect 3169 1462 3214 1467
rect 3233 1462 3286 1467
rect 3345 1462 3542 1467
rect 3561 1462 3670 1467
rect 3825 1462 4174 1467
rect 401 1457 406 1462
rect 305 1452 406 1457
rect 697 1457 702 1462
rect 3345 1457 3350 1462
rect 3689 1457 3806 1462
rect 697 1452 742 1457
rect 1009 1452 2070 1457
rect 2137 1452 2926 1457
rect 2945 1452 3350 1457
rect 3369 1452 3422 1457
rect 3457 1452 3694 1457
rect 3801 1452 3846 1457
rect 4049 1452 4158 1457
rect 2945 1447 2950 1452
rect 257 1442 366 1447
rect 601 1442 678 1447
rect 705 1442 742 1447
rect 777 1442 862 1447
rect 905 1442 1086 1447
rect 1161 1442 1230 1447
rect 1249 1442 1286 1447
rect 1337 1442 2102 1447
rect 2113 1442 2142 1447
rect 2153 1442 2214 1447
rect 2241 1442 2438 1447
rect 2457 1442 2838 1447
rect 2905 1442 2950 1447
rect 2969 1442 3070 1447
rect 3105 1442 3190 1447
rect 3217 1442 3302 1447
rect 3353 1442 3518 1447
rect 3545 1442 3590 1447
rect 3689 1442 3822 1447
rect 3873 1442 3974 1447
rect 3993 1442 4038 1447
rect 4081 1442 4246 1447
rect 601 1437 606 1442
rect 321 1432 606 1437
rect 673 1437 678 1442
rect 737 1437 742 1442
rect 2433 1437 2438 1442
rect 673 1432 726 1437
rect 737 1432 774 1437
rect 833 1432 902 1437
rect 929 1432 1374 1437
rect 1481 1432 1902 1437
rect 1913 1432 2070 1437
rect 2105 1432 2198 1437
rect 2321 1432 2374 1437
rect 2433 1432 2478 1437
rect 2537 1432 2558 1437
rect 2569 1432 2606 1437
rect 2617 1432 2654 1437
rect 2705 1432 2758 1437
rect 2889 1432 3006 1437
rect 3145 1432 3366 1437
rect 3401 1432 3462 1437
rect 3497 1432 3798 1437
rect 193 1422 294 1427
rect 321 1417 326 1432
rect 721 1427 726 1432
rect 1369 1427 1486 1432
rect 2065 1427 2070 1432
rect 2369 1427 2374 1432
rect 2777 1427 2870 1432
rect 3873 1427 3878 1442
rect 3969 1437 3974 1442
rect 3969 1432 4246 1437
rect 617 1422 710 1427
rect 721 1422 1350 1427
rect 1505 1417 1510 1427
rect 1537 1422 2046 1427
rect 2065 1422 2358 1427
rect 2369 1422 2470 1427
rect 2489 1422 2534 1427
rect 2641 1422 2782 1427
rect 2865 1422 3270 1427
rect 3409 1422 3542 1427
rect 3641 1422 3718 1427
rect 3785 1422 3902 1427
rect 3929 1422 4030 1427
rect 4097 1422 4230 1427
rect 2465 1417 2470 1422
rect 89 1412 182 1417
rect 177 1407 182 1412
rect 249 1412 326 1417
rect 425 1412 598 1417
rect 673 1412 942 1417
rect 961 1412 1046 1417
rect 1097 1412 1190 1417
rect 1289 1412 1414 1417
rect 1505 1412 1550 1417
rect 1665 1412 2206 1417
rect 2305 1412 2454 1417
rect 2465 1412 2886 1417
rect 3105 1412 3150 1417
rect 3281 1412 3326 1417
rect 3369 1412 3462 1417
rect 3513 1412 3862 1417
rect 4041 1412 4086 1417
rect 249 1407 254 1412
rect 425 1407 430 1412
rect 177 1402 254 1407
rect 401 1402 430 1407
rect 593 1407 598 1412
rect 2201 1407 2310 1412
rect 2449 1407 2454 1412
rect 2905 1407 3110 1412
rect 3169 1407 3262 1412
rect 3857 1407 4046 1412
rect 4081 1407 4198 1412
rect 593 1402 1806 1407
rect 1849 1402 1902 1407
rect 1921 1402 1982 1407
rect 2025 1402 2182 1407
rect 2329 1402 2382 1407
rect 2449 1402 2534 1407
rect 2545 1402 2910 1407
rect 3129 1402 3174 1407
rect 3257 1402 3470 1407
rect 3569 1402 3646 1407
rect 2529 1397 2534 1402
rect 3729 1397 3838 1402
rect 441 1392 646 1397
rect 657 1392 998 1397
rect 1049 1392 1078 1397
rect 1161 1392 1222 1397
rect 1249 1392 1462 1397
rect 1585 1392 1662 1397
rect 1673 1392 1710 1397
rect 1721 1392 1750 1397
rect 1761 1392 1862 1397
rect 1921 1392 1958 1397
rect 1969 1392 1998 1397
rect 2009 1392 2054 1397
rect 2121 1392 2166 1397
rect 2241 1392 2294 1397
rect 2305 1392 2350 1397
rect 2529 1392 2670 1397
rect 2793 1392 2822 1397
rect 2849 1392 2950 1397
rect 2993 1392 3014 1397
rect 3081 1392 3462 1397
rect 3513 1392 3542 1397
rect 3617 1392 3734 1397
rect 3833 1392 3862 1397
rect 3921 1392 4022 1397
rect 4041 1392 4158 1397
rect 2289 1387 2294 1392
rect 2665 1387 2798 1392
rect 3617 1387 3622 1392
rect 3921 1387 3926 1392
rect 393 1382 422 1387
rect 513 1382 702 1387
rect 817 1382 838 1387
rect 961 1382 990 1387
rect 1265 1382 2246 1387
rect 2289 1382 2310 1387
rect 2337 1382 2406 1387
rect 2417 1382 2598 1387
rect 2625 1382 2646 1387
rect 2817 1382 2862 1387
rect 2881 1382 3110 1387
rect 3161 1382 3254 1387
rect 3289 1382 3622 1387
rect 3745 1382 3926 1387
rect 4017 1387 4022 1392
rect 4177 1387 4182 1397
rect 4017 1382 4182 1387
rect 4193 1387 4198 1407
rect 4225 1402 4230 1422
rect 4257 1402 4366 1407
rect 4217 1392 4310 1397
rect 4193 1382 4270 1387
rect 417 1377 518 1382
rect 1009 1377 1246 1382
rect 2337 1377 2342 1382
rect 537 1372 622 1377
rect 641 1372 1014 1377
rect 1241 1372 1598 1377
rect 1609 1372 1878 1377
rect 1889 1372 1950 1377
rect 1993 1372 2206 1377
rect 2233 1372 2342 1377
rect 2369 1372 2398 1377
rect 2489 1372 2662 1377
rect 2673 1372 3190 1377
rect 3265 1372 3454 1377
rect 3489 1372 3566 1377
rect 3633 1372 3718 1377
rect 3769 1372 3990 1377
rect 4281 1372 4358 1377
rect 1873 1367 1878 1372
rect 2393 1367 2494 1372
rect 2657 1367 2662 1372
rect 3985 1367 4070 1372
rect 4153 1367 4286 1372
rect 113 1362 286 1367
rect 465 1362 526 1367
rect 809 1362 870 1367
rect 1017 1362 1174 1367
rect 1185 1362 1262 1367
rect 1377 1362 1422 1367
rect 1449 1362 1534 1367
rect 1585 1362 1638 1367
rect 1825 1362 1854 1367
rect 1873 1362 2022 1367
rect 2049 1362 2070 1367
rect 2161 1362 2254 1367
rect 2265 1362 2374 1367
rect 2513 1362 2542 1367
rect 2585 1362 2630 1367
rect 2657 1362 2798 1367
rect 2857 1362 3086 1367
rect 3169 1362 3838 1367
rect 4065 1362 4158 1367
rect 465 1357 470 1362
rect 521 1357 790 1362
rect 1169 1357 1174 1362
rect 1257 1357 1382 1362
rect 1721 1357 1806 1362
rect 2161 1357 2166 1362
rect 209 1352 470 1357
rect 785 1352 1134 1357
rect 1169 1352 1238 1357
rect 1513 1352 1534 1357
rect 1577 1352 1726 1357
rect 1801 1352 2166 1357
rect 2177 1352 3454 1357
rect 3465 1352 3590 1357
rect 3769 1352 3790 1357
rect 3921 1352 4046 1357
rect 4177 1352 4286 1357
rect 1233 1347 1238 1352
rect 1401 1347 1494 1352
rect 3609 1347 3750 1352
rect 3809 1347 3902 1352
rect 121 1342 222 1347
rect 481 1342 598 1347
rect 689 1342 726 1347
rect 785 1342 870 1347
rect 953 1342 1046 1347
rect 1185 1342 1222 1347
rect 1233 1342 1406 1347
rect 1489 1342 1630 1347
rect 1737 1342 2110 1347
rect 2353 1342 2398 1347
rect 2473 1342 2758 1347
rect 2785 1342 2822 1347
rect 2833 1342 3310 1347
rect 3377 1342 3406 1347
rect 3489 1342 3614 1347
rect 3745 1342 3814 1347
rect 3897 1342 4206 1347
rect 4217 1342 4310 1347
rect 593 1337 598 1342
rect 1625 1337 1742 1342
rect 2169 1337 2326 1342
rect 497 1332 582 1337
rect 593 1332 686 1337
rect 697 1332 782 1337
rect 873 1332 966 1337
rect 1065 1332 1166 1337
rect 1241 1332 1398 1337
rect 1417 1332 1486 1337
rect 1505 1332 1606 1337
rect 1761 1332 1846 1337
rect 1913 1332 1942 1337
rect 2009 1332 2046 1337
rect 2145 1332 2174 1337
rect 2321 1332 2990 1337
rect 3057 1332 3166 1337
rect 3201 1332 3238 1337
rect 3361 1332 3414 1337
rect 3425 1332 4110 1337
rect 4257 1332 4366 1337
rect 985 1327 1070 1332
rect 1161 1327 1166 1332
rect 3361 1327 3366 1332
rect 369 1322 990 1327
rect 1161 1322 1358 1327
rect 1569 1322 2134 1327
rect 2153 1322 2310 1327
rect 2409 1322 2790 1327
rect 2809 1322 2870 1327
rect 3041 1322 3062 1327
rect 3089 1322 3182 1327
rect 3209 1322 3366 1327
rect 3417 1322 3934 1327
rect 3969 1322 4030 1327
rect 4049 1322 4126 1327
rect 4193 1322 4222 1327
rect 2865 1317 2870 1322
rect 4049 1317 4054 1322
rect 201 1312 238 1317
rect 545 1312 590 1317
rect 641 1312 670 1317
rect 729 1312 1222 1317
rect 1345 1312 1478 1317
rect 1713 1312 1854 1317
rect 1889 1312 2190 1317
rect 2201 1312 2606 1317
rect 2777 1312 2854 1317
rect 2865 1312 2918 1317
rect 2977 1312 3094 1317
rect 3105 1312 3230 1317
rect 3313 1312 3862 1317
rect 3889 1312 4054 1317
rect 3225 1307 3318 1312
rect 3889 1307 3894 1312
rect 545 1302 622 1307
rect 657 1302 742 1307
rect 833 1302 902 1307
rect 1017 1302 1158 1307
rect 1177 1302 1214 1307
rect 1233 1302 1374 1307
rect 1489 1302 3206 1307
rect 3337 1302 3414 1307
rect 3641 1302 3894 1307
rect 3913 1302 3998 1307
rect 1369 1297 1494 1302
rect 3537 1297 3646 1302
rect 4193 1297 4198 1322
rect 409 1292 1174 1297
rect 1265 1292 1350 1297
rect 1705 1292 1790 1297
rect 1801 1292 2126 1297
rect 2249 1292 3230 1297
rect 3265 1292 3542 1297
rect 3665 1292 4254 1297
rect 1169 1287 1270 1292
rect 377 1282 454 1287
rect 521 1282 630 1287
rect 657 1282 718 1287
rect 713 1277 718 1282
rect 801 1282 830 1287
rect 889 1282 966 1287
rect 985 1282 1150 1287
rect 1433 1282 1942 1287
rect 1953 1282 2038 1287
rect 2089 1282 2254 1287
rect 2401 1282 2518 1287
rect 2529 1282 2726 1287
rect 2753 1282 3950 1287
rect 4009 1282 4038 1287
rect 4169 1282 4270 1287
rect 801 1277 806 1282
rect 1937 1277 1942 1282
rect 2249 1277 2406 1282
rect 585 1272 694 1277
rect 713 1272 806 1277
rect 929 1272 1406 1277
rect 1489 1272 1830 1277
rect 1865 1272 1902 1277
rect 1937 1272 2046 1277
rect 2065 1272 2166 1277
rect 2185 1272 2230 1277
rect 2425 1272 2462 1277
rect 1489 1267 1494 1272
rect 2513 1267 2518 1282
rect 2537 1272 3302 1277
rect 3345 1272 3446 1277
rect 3457 1272 3502 1277
rect 3697 1272 3726 1277
rect 3809 1272 3838 1277
rect 4129 1272 4150 1277
rect 3721 1267 3814 1272
rect 4009 1267 4102 1272
rect 529 1262 574 1267
rect 873 1262 1094 1267
rect 1153 1262 1190 1267
rect 1353 1262 1494 1267
rect 1529 1262 2294 1267
rect 2329 1262 2382 1267
rect 2513 1262 3550 1267
rect 3857 1262 3966 1267
rect 3985 1262 4014 1267
rect 4097 1262 4126 1267
rect 593 1257 758 1262
rect 3857 1257 3862 1262
rect 273 1252 334 1257
rect 457 1252 598 1257
rect 753 1252 910 1257
rect 961 1252 1054 1257
rect 1217 1252 1254 1257
rect 1313 1252 1382 1257
rect 1457 1252 1614 1257
rect 1633 1252 1974 1257
rect 2001 1252 2118 1257
rect 2137 1252 2310 1257
rect 2321 1252 2470 1257
rect 2521 1252 2950 1257
rect 3001 1252 3030 1257
rect 3049 1252 3118 1257
rect 3145 1252 3174 1257
rect 3297 1252 3646 1257
rect 3697 1252 3862 1257
rect 3961 1257 3966 1262
rect 3961 1252 4190 1257
rect 1073 1247 1182 1252
rect 3025 1247 3030 1252
rect 473 1242 1078 1247
rect 1177 1242 1734 1247
rect 1761 1242 1878 1247
rect 1977 1242 1998 1247
rect 2033 1242 2182 1247
rect 2201 1242 2254 1247
rect 2265 1242 2430 1247
rect 2449 1242 2534 1247
rect 1761 1237 1766 1242
rect 2577 1237 2582 1247
rect 2601 1242 2662 1247
rect 2705 1242 2814 1247
rect 2993 1237 2998 1247
rect 3025 1242 3046 1247
rect 3057 1242 3134 1247
rect 3385 1242 3510 1247
rect 3625 1242 3766 1247
rect 3873 1242 4150 1247
rect 305 1232 502 1237
rect 601 1232 638 1237
rect 665 1232 926 1237
rect 961 1232 1166 1237
rect 1257 1232 1766 1237
rect 1785 1232 2838 1237
rect 2881 1232 2958 1237
rect 2993 1232 3070 1237
rect 3121 1232 3174 1237
rect 3233 1232 3270 1237
rect 3369 1232 3494 1237
rect 305 1227 310 1232
rect 2881 1227 2886 1232
rect 3121 1227 3126 1232
rect 3505 1227 3510 1242
rect 3761 1237 3878 1242
rect 4145 1237 4150 1242
rect 3545 1232 3662 1237
rect 3713 1232 3742 1237
rect 3921 1232 4078 1237
rect 4145 1232 4294 1237
rect 145 1222 198 1227
rect 225 1222 334 1227
rect 345 1222 430 1227
rect 425 1217 430 1222
rect 513 1222 846 1227
rect 889 1222 926 1227
rect 937 1222 1078 1227
rect 1097 1222 1126 1227
rect 1145 1222 1238 1227
rect 1273 1222 1302 1227
rect 1321 1222 1534 1227
rect 1577 1222 1974 1227
rect 1993 1222 2366 1227
rect 2433 1222 2470 1227
rect 2489 1222 2526 1227
rect 2545 1222 2654 1227
rect 2705 1222 2782 1227
rect 2793 1222 2886 1227
rect 2905 1222 3126 1227
rect 3193 1222 3270 1227
rect 3337 1222 3398 1227
rect 3417 1222 3454 1227
rect 3505 1222 3942 1227
rect 513 1217 518 1222
rect 2465 1217 2470 1222
rect 425 1212 518 1217
rect 569 1212 1742 1217
rect 1801 1212 1902 1217
rect 1937 1212 2006 1217
rect 2313 1212 2358 1217
rect 2401 1212 2446 1217
rect 2465 1212 2510 1217
rect 2561 1212 2614 1217
rect 2753 1212 2966 1217
rect 3097 1212 3310 1217
rect 3441 1212 3494 1217
rect 3537 1212 3574 1217
rect 3649 1212 3726 1217
rect 3953 1212 4070 1217
rect 2025 1207 2174 1212
rect 2217 1207 2294 1212
rect 2609 1207 2614 1212
rect 3329 1207 3422 1212
rect 3721 1207 3958 1212
rect 193 1202 406 1207
rect 601 1202 638 1207
rect 921 1202 958 1207
rect 1049 1202 2030 1207
rect 2169 1202 2222 1207
rect 2289 1202 2398 1207
rect 2409 1202 2486 1207
rect 2513 1202 2598 1207
rect 2609 1202 2742 1207
rect 2833 1202 3334 1207
rect 3417 1202 3702 1207
rect 713 1197 902 1202
rect 2593 1197 2598 1202
rect 2737 1197 2838 1202
rect 521 1192 590 1197
rect 625 1192 678 1197
rect 689 1192 718 1197
rect 897 1192 1710 1197
rect 1817 1192 1862 1197
rect 1881 1192 1926 1197
rect 1977 1192 2022 1197
rect 2073 1192 2158 1197
rect 2233 1192 2310 1197
rect 2449 1192 2502 1197
rect 2593 1192 2654 1197
rect 2857 1192 3030 1197
rect 3153 1192 3182 1197
rect 3193 1192 3238 1197
rect 3273 1192 3382 1197
rect 3393 1192 3414 1197
rect 3425 1192 3478 1197
rect 3521 1192 3566 1197
rect 3593 1192 3638 1197
rect 3665 1192 3742 1197
rect 3761 1192 3806 1197
rect 3857 1192 3918 1197
rect 3929 1192 4030 1197
rect 2329 1187 2430 1192
rect 3857 1187 3862 1192
rect 177 1182 910 1187
rect 929 1182 1102 1187
rect 1161 1182 1222 1187
rect 1281 1182 1382 1187
rect 1393 1182 1438 1187
rect 1481 1182 1582 1187
rect 1753 1182 1846 1187
rect 1897 1182 2070 1187
rect 2225 1182 2334 1187
rect 2425 1182 3230 1187
rect 3273 1182 3302 1187
rect 3361 1182 3862 1187
rect 3881 1182 4118 1187
rect 4289 1182 4358 1187
rect 929 1177 934 1182
rect 2225 1177 2230 1182
rect 465 1172 494 1177
rect 569 1172 614 1177
rect 625 1172 654 1177
rect 665 1172 702 1177
rect 721 1172 742 1177
rect 801 1172 934 1177
rect 985 1172 1006 1177
rect 1033 1172 1374 1177
rect 1401 1172 1502 1177
rect 1521 1172 2230 1177
rect 2241 1172 2270 1177
rect 2337 1172 2542 1177
rect 2577 1172 2598 1177
rect 2633 1172 2678 1177
rect 2753 1172 2798 1177
rect 2841 1172 2926 1177
rect 2945 1172 3014 1177
rect 3025 1172 3046 1177
rect 3073 1172 3134 1177
rect 3161 1172 3206 1177
rect 3265 1172 3430 1177
rect 3441 1172 3494 1177
rect 3537 1172 3678 1177
rect 3705 1172 3726 1177
rect 3833 1172 3862 1177
rect 3913 1172 3974 1177
rect 4089 1172 4286 1177
rect 1521 1167 1526 1172
rect 161 1162 206 1167
rect 449 1162 734 1167
rect 881 1162 1006 1167
rect 1017 1162 1302 1167
rect 729 1157 886 1162
rect 169 1152 246 1157
rect 361 1152 710 1157
rect 905 1152 958 1157
rect 985 1152 1054 1157
rect 1145 1152 1206 1157
rect 1217 1152 1286 1157
rect 241 1147 246 1152
rect 1201 1147 1206 1152
rect 1297 1147 1302 1162
rect 1321 1162 1350 1167
rect 1401 1162 1526 1167
rect 1545 1162 1614 1167
rect 1737 1162 3126 1167
rect 3145 1162 3198 1167
rect 3385 1162 3414 1167
rect 3545 1162 3590 1167
rect 3601 1162 3654 1167
rect 3713 1162 3774 1167
rect 3841 1162 4166 1167
rect 4225 1162 4318 1167
rect 1321 1152 1326 1162
rect 3121 1157 3126 1162
rect 3217 1157 3366 1162
rect 3433 1157 3526 1162
rect 1337 1152 1422 1157
rect 1441 1152 1574 1157
rect 1633 1152 1798 1157
rect 1817 1152 1918 1157
rect 2033 1152 2182 1157
rect 2289 1152 2838 1157
rect 2865 1152 3102 1157
rect 3121 1152 3222 1157
rect 3361 1152 3438 1157
rect 3521 1152 3958 1157
rect 4097 1152 4142 1157
rect 1441 1147 1446 1152
rect 2033 1147 2038 1152
rect 3977 1147 4078 1152
rect 4161 1147 4286 1152
rect 177 1142 222 1147
rect 241 1142 374 1147
rect 385 1142 478 1147
rect 577 1142 646 1147
rect 673 1142 806 1147
rect 889 1142 958 1147
rect 985 1142 1094 1147
rect 1105 1142 1166 1147
rect 1201 1142 1246 1147
rect 1297 1142 1446 1147
rect 417 1132 670 1137
rect 857 1132 918 1137
rect 929 1132 998 1137
rect 1025 1132 1030 1142
rect 1089 1137 1094 1142
rect 1457 1137 1462 1147
rect 1497 1142 1558 1147
rect 1585 1142 1606 1147
rect 1705 1142 1734 1147
rect 1809 1142 1838 1147
rect 1921 1142 1974 1147
rect 2009 1142 2038 1147
rect 2049 1142 2110 1147
rect 2281 1142 2326 1147
rect 2393 1142 3254 1147
rect 3305 1142 3366 1147
rect 3377 1142 3510 1147
rect 3609 1142 3662 1147
rect 3681 1142 3726 1147
rect 3737 1142 3854 1147
rect 3873 1142 3982 1147
rect 4073 1142 4166 1147
rect 4281 1142 4310 1147
rect 2129 1137 2246 1142
rect 1041 1132 1078 1137
rect 1089 1132 1478 1137
rect 1585 1132 1638 1137
rect 1721 1132 2134 1137
rect 2241 1132 3606 1137
rect 993 1127 998 1132
rect 1073 1127 1078 1132
rect 169 1122 350 1127
rect 369 1122 430 1127
rect 697 1122 966 1127
rect 993 1122 1062 1127
rect 1073 1122 1406 1127
rect 1553 1122 1654 1127
rect 1713 1122 1758 1127
rect 1817 1122 1854 1127
rect 1913 1122 1982 1127
rect 2025 1122 2230 1127
rect 2321 1122 2686 1127
rect 2713 1122 2790 1127
rect 3145 1122 3182 1127
rect 3233 1122 3270 1127
rect 3337 1122 3358 1127
rect 3385 1122 3446 1127
rect 169 1117 174 1122
rect 145 1112 174 1117
rect 345 1117 350 1122
rect 449 1117 606 1122
rect 1057 1117 1062 1122
rect 2809 1117 3126 1122
rect 3465 1117 3566 1122
rect 3601 1117 3606 1132
rect 3681 1127 3686 1142
rect 3745 1132 3790 1137
rect 3865 1132 4366 1137
rect 3681 1122 3710 1127
rect 3777 1122 3806 1127
rect 3849 1122 3894 1127
rect 3945 1122 4054 1127
rect 4137 1122 4198 1127
rect 4193 1117 4198 1122
rect 345 1112 454 1117
rect 601 1112 790 1117
rect 913 1112 958 1117
rect 977 1112 1030 1117
rect 1057 1112 2406 1117
rect 2521 1112 2670 1117
rect 2681 1112 2814 1117
rect 3121 1112 3470 1117
rect 3561 1112 3590 1117
rect 3601 1112 3982 1117
rect 3993 1112 4086 1117
rect 4193 1112 4222 1117
rect 2401 1107 2502 1112
rect 153 1102 590 1107
rect 769 1102 822 1107
rect 849 1102 1174 1107
rect 1209 1102 1254 1107
rect 1353 1102 1422 1107
rect 1521 1102 2206 1107
rect 2217 1102 2350 1107
rect 2361 1102 2382 1107
rect 2497 1102 3110 1107
rect 3145 1102 3190 1107
rect 3225 1102 3326 1107
rect 3353 1102 3374 1107
rect 3417 1102 3566 1107
rect 3585 1102 3590 1112
rect 3697 1102 3790 1107
rect 3809 1102 4182 1107
rect 4241 1102 4270 1107
rect 4361 1102 4390 1107
rect 3105 1097 3110 1102
rect 4177 1097 4246 1102
rect 193 1092 238 1097
rect 305 1092 382 1097
rect 809 1092 878 1097
rect 889 1092 1870 1097
rect 1993 1092 2022 1097
rect 2081 1092 2126 1097
rect 2145 1092 2678 1097
rect 2705 1092 2758 1097
rect 2769 1092 2814 1097
rect 2841 1092 2918 1097
rect 2961 1092 3094 1097
rect 3105 1092 3158 1097
rect 2145 1087 2150 1092
rect 3233 1087 3238 1097
rect 3249 1092 3310 1097
rect 3329 1092 3838 1097
rect 3953 1092 4022 1097
rect 4385 1087 4390 1102
rect 265 1082 366 1087
rect 361 1077 366 1082
rect 457 1082 486 1087
rect 609 1082 750 1087
rect 785 1082 926 1087
rect 937 1082 982 1087
rect 1001 1082 1118 1087
rect 1305 1082 1334 1087
rect 1409 1082 2150 1087
rect 2201 1082 3078 1087
rect 3089 1082 3118 1087
rect 3233 1082 3382 1087
rect 3393 1082 3470 1087
rect 3545 1082 3598 1087
rect 3657 1082 4150 1087
rect 4225 1082 4390 1087
rect 457 1077 462 1082
rect 609 1077 614 1082
rect 161 1072 190 1077
rect 185 1067 190 1072
rect 297 1072 342 1077
rect 361 1072 462 1077
rect 569 1072 614 1077
rect 745 1077 750 1082
rect 1209 1077 1286 1082
rect 4225 1077 4230 1082
rect 745 1072 1214 1077
rect 1281 1072 1526 1077
rect 1585 1072 1606 1077
rect 1625 1072 1766 1077
rect 1833 1072 1926 1077
rect 1961 1072 3262 1077
rect 3305 1072 3878 1077
rect 3897 1072 3918 1077
rect 3977 1072 4230 1077
rect 297 1067 302 1072
rect 185 1062 302 1067
rect 817 1062 998 1067
rect 1009 1062 1030 1067
rect 1225 1062 1462 1067
rect 1545 1062 2222 1067
rect 2233 1062 2558 1067
rect 2585 1062 2630 1067
rect 2689 1062 2854 1067
rect 2881 1062 2990 1067
rect 3009 1062 3142 1067
rect 3153 1062 3294 1067
rect 3313 1062 3382 1067
rect 3401 1062 4182 1067
rect 689 1057 798 1062
rect 1057 1057 1182 1062
rect 2881 1057 2886 1062
rect 3313 1057 3318 1062
rect 4177 1057 4182 1062
rect 513 1052 694 1057
rect 793 1052 958 1057
rect 1033 1052 1062 1057
rect 1177 1052 2150 1057
rect 2313 1052 2766 1057
rect 2825 1052 2886 1057
rect 3017 1052 3158 1057
rect 3193 1052 3262 1057
rect 3297 1052 3318 1057
rect 3337 1052 3518 1057
rect 3641 1052 3670 1057
rect 3681 1052 3766 1057
rect 3793 1052 3862 1057
rect 3945 1052 4006 1057
rect 4177 1052 4238 1057
rect 2169 1047 2294 1052
rect 2905 1047 2998 1052
rect 4001 1047 4006 1052
rect 321 1042 494 1047
rect 705 1042 1622 1047
rect 1697 1042 1758 1047
rect 1841 1042 2174 1047
rect 2289 1042 2910 1047
rect 2993 1042 3990 1047
rect 4001 1042 4166 1047
rect 321 1037 326 1042
rect 297 1032 326 1037
rect 489 1037 494 1042
rect 1841 1037 1846 1042
rect 4161 1037 4166 1042
rect 4249 1042 4326 1047
rect 4249 1037 4254 1042
rect 489 1032 574 1037
rect 593 1032 1550 1037
rect 1633 1032 1678 1037
rect 1705 1032 1750 1037
rect 1761 1032 1814 1037
rect 1825 1032 1846 1037
rect 1865 1032 4006 1037
rect 4161 1032 4254 1037
rect 4369 1032 4374 1082
rect 369 1027 470 1032
rect 1825 1027 1830 1032
rect 73 1022 118 1027
rect 177 1022 326 1027
rect 345 1022 374 1027
rect 465 1022 806 1027
rect 921 1022 950 1027
rect 961 1022 1022 1027
rect 1113 1022 1254 1027
rect 1265 1022 1286 1027
rect 1393 1022 1614 1027
rect 1697 1022 1830 1027
rect 1841 1022 2158 1027
rect 2273 1022 2726 1027
rect 2737 1022 2862 1027
rect 2953 1022 3014 1027
rect 3113 1022 3230 1027
rect 3273 1022 3326 1027
rect 3377 1022 3422 1027
rect 3441 1022 3782 1027
rect 3865 1022 3934 1027
rect 3985 1022 4030 1027
rect 321 1017 326 1022
rect 1697 1017 1702 1022
rect 321 1012 470 1017
rect 817 1012 846 1017
rect 881 1012 1702 1017
rect 1745 1012 1782 1017
rect 465 1007 822 1012
rect 1841 1007 1846 1022
rect 2153 1017 2158 1022
rect 3441 1017 3446 1022
rect 1921 1012 1974 1017
rect 1993 1012 2078 1017
rect 2153 1012 2342 1017
rect 2369 1012 3254 1017
rect 3273 1012 3310 1017
rect 3377 1012 3446 1017
rect 3473 1012 3910 1017
rect 4033 1012 4062 1017
rect 4089 1012 4206 1017
rect 281 1002 374 1007
rect 417 1002 446 1007
rect 865 1002 966 1007
rect 1009 1002 1846 1007
rect 2041 1002 2062 1007
rect 2369 997 2374 1012
rect 4089 1007 4094 1012
rect 2401 1002 2486 1007
rect 2521 1002 2686 1007
rect 2705 1002 2854 1007
rect 2945 1002 2974 1007
rect 3073 1002 3110 1007
rect 3241 1002 3486 1007
rect 3505 1002 3718 1007
rect 3745 1002 3894 1007
rect 4001 1002 4094 1007
rect 4201 1007 4206 1012
rect 4201 1002 4350 1007
rect 2401 997 2406 1002
rect 3505 997 3510 1002
rect 113 992 214 997
rect 249 992 302 997
rect 329 992 414 997
rect 425 992 550 997
rect 585 992 654 997
rect 729 992 806 997
rect 881 992 958 997
rect 977 992 1966 997
rect 2009 992 2054 997
rect 2209 992 2278 997
rect 2305 992 2374 997
rect 2385 992 2406 997
rect 2425 992 2694 997
rect 2713 992 2766 997
rect 3001 992 3510 997
rect 3593 992 3630 997
rect 3689 992 3758 997
rect 3785 992 3830 997
rect 4137 992 4182 997
rect 2785 987 2942 992
rect 3849 987 3966 992
rect 273 982 310 987
rect 377 982 398 987
rect 721 982 878 987
rect 889 982 974 987
rect 1041 982 1097 987
rect 1105 982 1350 987
rect 1393 982 2022 987
rect 2081 982 2190 987
rect 2217 982 2790 987
rect 2937 982 2966 987
rect 2985 982 3046 987
rect 3073 982 3118 987
rect 3217 982 3262 987
rect 3313 982 3342 987
rect 3377 982 3414 987
rect 3673 982 3750 987
rect 3777 982 3854 987
rect 3961 982 4190 987
rect 4249 982 4342 987
rect 417 977 606 982
rect 1092 977 1097 982
rect 2081 977 2086 982
rect 257 972 278 977
rect 313 972 422 977
rect 601 972 710 977
rect 761 972 902 977
rect 929 972 1014 977
rect 1033 972 1086 977
rect 1092 972 1126 977
rect 1169 972 1238 977
rect 1249 972 1374 977
rect 1401 972 1446 977
rect 1489 972 2086 977
rect 2185 977 2190 982
rect 2185 972 3446 977
rect 3585 972 3670 977
rect 1009 967 1014 972
rect 3745 967 3750 982
rect 4249 977 4254 982
rect 3769 972 3822 977
rect 3833 972 3862 977
rect 3913 972 3950 977
rect 4049 972 4102 977
rect 4153 972 4254 977
rect 4337 977 4342 982
rect 4337 972 4382 977
rect 425 962 590 967
rect 673 962 702 967
rect 713 962 942 967
rect 1009 962 1094 967
rect 1201 962 1294 967
rect 1329 962 1422 967
rect 1433 962 1806 967
rect 1825 962 1918 967
rect 1945 962 2038 967
rect 2361 962 2902 967
rect 2913 962 2990 967
rect 3033 962 3102 967
rect 3201 962 3326 967
rect 3353 962 3406 967
rect 3449 962 3502 967
rect 3745 962 3838 967
rect 4257 962 4326 967
rect 585 957 678 962
rect 1825 957 1830 962
rect 2201 957 2342 962
rect 3521 957 3726 962
rect 3985 957 4238 962
rect 321 952 350 957
rect 385 952 502 957
rect 529 952 566 957
rect 721 952 846 957
rect 961 952 1158 957
rect 1241 952 1830 957
rect 1841 952 2206 957
rect 2337 952 3526 957
rect 3721 952 3990 957
rect 4233 952 4334 957
rect 145 942 254 947
rect 321 942 510 947
rect 321 937 326 942
rect 177 932 326 937
rect 337 932 414 937
rect 529 932 534 952
rect 1841 947 1846 952
rect 545 942 614 947
rect 737 942 774 947
rect 793 942 934 947
rect 969 942 1182 947
rect 1201 942 1470 947
rect 1569 942 1622 947
rect 1697 942 1766 947
rect 1785 942 1846 947
rect 1897 942 1950 947
rect 1961 942 1990 947
rect 2217 942 2358 947
rect 2441 942 2478 947
rect 2513 942 2534 947
rect 2561 942 2630 947
rect 2641 942 3150 947
rect 3257 942 3286 947
rect 3305 942 3398 947
rect 3417 942 3550 947
rect 3569 942 3598 947
rect 3609 942 3806 947
rect 3897 942 3958 947
rect 3977 942 4230 947
rect 4249 942 4318 947
rect 1201 937 1206 942
rect 2513 937 2518 942
rect 2641 937 2646 942
rect 3281 937 3286 942
rect 3801 937 3902 942
rect 3953 937 3958 942
rect 4225 937 4230 942
rect 577 932 758 937
rect 769 932 1118 937
rect 1153 932 1206 937
rect 1217 932 1270 937
rect 1497 932 1526 937
rect 1625 932 1958 937
rect 2009 932 2102 937
rect 2145 932 2518 937
rect 2625 932 2646 937
rect 2673 932 2726 937
rect 2849 932 2982 937
rect 3025 932 3150 937
rect 3281 932 3350 937
rect 3375 932 3390 937
rect 3585 932 3654 937
rect 3697 932 3782 937
rect 3921 932 3942 937
rect 3953 932 4190 937
rect 4225 932 4374 937
rect 441 927 534 932
rect 1385 927 1478 932
rect 2009 927 2014 932
rect 97 922 134 927
rect 417 922 446 927
rect 569 922 814 927
rect 873 922 1014 927
rect 1073 922 1110 927
rect 1121 922 1390 927
rect 1473 922 2014 927
rect 2097 927 2102 932
rect 2097 922 2134 927
rect 225 917 342 922
rect 2129 917 2134 922
rect 2225 922 2390 927
rect 2409 922 2438 927
rect 2449 922 2590 927
rect 2225 917 2230 922
rect 2625 917 2630 932
rect 2673 927 2678 932
rect 3025 927 3030 932
rect 3375 927 3380 932
rect 3937 927 3942 932
rect 2660 922 2678 927
rect 2713 922 2878 927
rect 2905 922 2942 927
rect 2953 922 3030 927
rect 3041 922 3070 927
rect 3089 922 3118 927
rect 3201 922 3380 927
rect 3433 922 3478 927
rect 3529 922 3638 927
rect 3657 922 3718 927
rect 3873 922 3926 927
rect 3937 922 4022 927
rect 4177 922 4382 927
rect 2660 917 2665 922
rect 3737 917 3854 922
rect 4177 917 4182 922
rect 177 912 230 917
rect 337 912 366 917
rect 481 912 558 917
rect 625 912 854 917
rect 881 912 926 917
rect 1025 912 1158 917
rect 1233 912 1286 917
rect 1401 912 1446 917
rect 1457 912 1638 917
rect 1697 912 1830 917
rect 1849 912 1910 917
rect 2009 912 2086 917
rect 2129 912 2230 917
rect 2249 912 2286 917
rect 2433 912 2630 917
rect 2649 912 2665 917
rect 2673 912 3038 917
rect 3185 912 3742 917
rect 3849 912 3878 917
rect 3913 912 4182 917
rect 4193 912 4270 917
rect 1457 907 1462 912
rect 257 902 398 907
rect 537 902 710 907
rect 817 902 902 907
rect 929 902 1126 907
rect 1161 902 1262 907
rect 1329 902 1430 907
rect 1457 902 1478 907
rect 1521 902 1566 907
rect 1729 902 1878 907
rect 1969 902 2030 907
rect 2273 902 2406 907
rect 2425 902 2486 907
rect 2505 902 2566 907
rect 2585 902 2838 907
rect 2897 902 2958 907
rect 2977 902 3102 907
rect 3161 902 3262 907
rect 3289 902 3670 907
rect 3681 902 3750 907
rect 3801 902 3846 907
rect 3865 902 3902 907
rect 4217 902 4358 907
rect 417 897 518 902
rect 2401 897 2406 902
rect 2833 897 2838 902
rect 3665 897 3670 902
rect 329 892 422 897
rect 513 892 558 897
rect 585 892 686 897
rect 705 892 1502 897
rect 1529 892 1934 897
rect 1961 892 2022 897
rect 2105 892 2230 897
rect 2297 892 2366 897
rect 2401 892 2502 897
rect 2553 892 2646 897
rect 2673 892 2822 897
rect 2833 892 3390 897
rect 3465 892 3622 897
rect 3665 892 4070 897
rect 2105 887 2110 892
rect 289 882 982 887
rect 1113 882 1374 887
rect 1729 882 2110 887
rect 2225 887 2230 892
rect 3617 887 3622 892
rect 4065 887 4070 892
rect 2225 882 2870 887
rect 2881 882 3198 887
rect 3241 882 3606 887
rect 3617 882 3702 887
rect 4065 882 4278 887
rect 1025 877 1094 882
rect 1449 877 1686 882
rect 185 872 606 877
rect 769 872 1030 877
rect 1089 872 1454 877
rect 1681 872 1710 877
rect 625 867 750 872
rect 1729 867 1734 882
rect 2865 877 2870 882
rect 3721 877 3934 882
rect 1809 872 1966 877
rect 2201 872 2294 877
rect 2305 872 2470 877
rect 2521 872 2702 877
rect 2777 872 2814 877
rect 2865 872 3358 877
rect 3497 872 3726 877
rect 3929 872 3958 877
rect 2305 867 2310 872
rect 297 862 462 867
rect 545 862 630 867
rect 745 862 974 867
rect 1041 862 1230 867
rect 1257 862 1326 867
rect 1465 862 1734 867
rect 1817 862 2174 867
rect 2233 862 2310 867
rect 2329 862 2614 867
rect 2665 862 2694 867
rect 2761 862 2870 867
rect 2889 862 2926 867
rect 2969 862 3142 867
rect 3169 862 3206 867
rect 3265 862 3334 867
rect 3385 862 3910 867
rect 4089 862 4286 867
rect 1345 857 1446 862
rect 3201 857 3206 862
rect 377 852 398 857
rect 409 852 486 857
rect 513 852 902 857
rect 921 852 1030 857
rect 1137 852 1350 857
rect 1441 852 1534 857
rect 1713 852 1766 857
rect 1865 852 1910 857
rect 1937 852 2030 857
rect 2241 852 2278 857
rect 2329 852 3174 857
rect 3201 852 3342 857
rect 3361 852 3918 857
rect 4289 852 4366 857
rect 1553 847 1694 852
rect 305 842 446 847
rect 441 837 446 842
rect 561 842 662 847
rect 745 842 806 847
rect 817 842 1006 847
rect 1121 842 1166 847
rect 1249 842 1558 847
rect 1689 842 2094 847
rect 2137 842 2206 847
rect 2225 842 2350 847
rect 2449 842 2478 847
rect 2513 842 2542 847
rect 2585 842 2638 847
rect 2777 842 2830 847
rect 2905 842 2982 847
rect 3057 842 3102 847
rect 3121 842 3214 847
rect 3273 842 3326 847
rect 3361 842 3942 847
rect 3969 842 4246 847
rect 561 837 566 842
rect 1161 837 1254 842
rect 2137 837 2142 842
rect 289 832 318 837
rect 353 832 422 837
rect 441 832 566 837
rect 585 832 662 837
rect 857 832 934 837
rect 1025 832 1142 837
rect 1393 832 1606 837
rect 1617 832 1750 837
rect 1769 832 1798 837
rect 1929 832 2142 837
rect 2201 837 2206 842
rect 2657 837 2758 842
rect 2201 832 2662 837
rect 2753 832 3438 837
rect 3545 832 3830 837
rect 3905 832 4062 837
rect 4289 832 4374 837
rect 289 827 294 832
rect 761 827 838 832
rect 1273 827 1374 832
rect 3433 827 3550 832
rect 4289 827 4294 832
rect 185 822 294 827
rect 313 822 382 827
rect 633 822 766 827
rect 833 822 1278 827
rect 1369 822 1790 827
rect 1913 822 1974 827
rect 1985 822 2334 827
rect 2385 822 3414 827
rect 3569 822 3590 827
rect 3689 822 3894 827
rect 4009 822 4294 827
rect 1985 817 1990 822
rect 3585 817 3662 822
rect 3889 817 4014 822
rect 4305 817 4310 827
rect 433 812 518 817
rect 553 812 670 817
rect 777 812 830 817
rect 881 812 1158 817
rect 1289 812 1326 817
rect 1361 812 1990 817
rect 2225 812 3134 817
rect 881 807 886 812
rect 2009 807 2230 812
rect 3145 807 3150 817
rect 3273 812 3462 817
rect 3657 812 3774 817
rect 4033 812 4086 817
rect 4129 812 4182 817
rect 4233 812 4310 817
rect 337 802 358 807
rect 385 802 454 807
rect 489 802 718 807
rect 753 802 886 807
rect 905 802 1206 807
rect 1217 802 1358 807
rect 1369 802 2014 807
rect 2241 802 2534 807
rect 2545 802 2566 807
rect 2585 802 2662 807
rect 2713 802 2814 807
rect 2889 802 2990 807
rect 3009 802 3062 807
rect 3121 802 3150 807
rect 3161 802 3310 807
rect 3337 802 3390 807
rect 3441 802 3502 807
rect 3585 802 3646 807
rect 3737 802 3878 807
rect 3937 802 3974 807
rect 4033 802 4038 812
rect 4129 802 4134 812
rect 4225 802 4310 807
rect 1201 797 1206 802
rect 137 792 214 797
rect 225 792 286 797
rect 465 792 486 797
rect 497 792 518 797
rect 761 792 862 797
rect 1009 792 1126 797
rect 1201 792 1454 797
rect 1649 792 1918 797
rect 1977 792 2142 797
rect 2169 792 2198 797
rect 2257 792 2342 797
rect 2361 792 3470 797
rect 3537 792 3638 797
rect 3665 792 3766 797
rect 3801 792 3902 797
rect 4033 792 4070 797
rect 4145 792 4182 797
rect 537 787 742 792
rect 1449 787 1542 792
rect 1649 787 1654 792
rect 393 782 542 787
rect 737 782 838 787
rect 865 782 894 787
rect 953 782 982 787
rect 993 782 1046 787
rect 1169 782 1206 787
rect 1329 782 1430 787
rect 1537 782 1654 787
rect 1673 782 1758 787
rect 1785 782 1902 787
rect 1945 782 2030 787
rect 2097 782 2366 787
rect 2385 782 2486 787
rect 2521 782 2606 787
rect 2673 782 2710 787
rect 2785 782 2870 787
rect 2953 782 3014 787
rect 3025 782 3142 787
rect 3185 782 3358 787
rect 3377 782 3478 787
rect 3521 782 3710 787
rect 3745 782 4134 787
rect 4193 782 4262 787
rect 4129 777 4198 782
rect 297 772 838 777
rect 849 772 1038 777
rect 1153 772 1182 777
rect 1193 772 1374 777
rect 1449 772 1518 777
rect 1769 772 1886 777
rect 1969 772 2342 777
rect 2425 772 2486 777
rect 2577 772 3142 777
rect 3249 772 3550 777
rect 3705 772 3870 777
rect 849 767 854 772
rect 1449 767 1454 772
rect 257 762 854 767
rect 873 762 1454 767
rect 1513 767 1518 772
rect 3137 767 3254 772
rect 3569 767 3686 772
rect 3921 767 4070 772
rect 1513 762 1758 767
rect 1817 762 2494 767
rect 2505 762 2830 767
rect 2985 762 3078 767
rect 3089 762 3118 767
rect 3273 762 3326 767
rect 3353 762 3574 767
rect 3681 762 3878 767
rect 3897 762 3926 767
rect 4065 762 4214 767
rect 1753 757 1822 762
rect 2849 757 2966 762
rect 3873 757 3878 762
rect 65 752 782 757
rect 801 752 918 757
rect 929 752 1006 757
rect 1113 752 1238 757
rect 1249 752 1286 757
rect 1321 752 1502 757
rect 1841 752 1894 757
rect 1937 752 2126 757
rect 2177 752 2246 757
rect 2289 752 2358 757
rect 2449 752 2606 757
rect 2617 752 2854 757
rect 2961 752 3246 757
rect 3297 752 3414 757
rect 3505 752 3654 757
rect 3697 752 3798 757
rect 3873 752 4070 757
rect 289 742 374 747
rect 385 742 542 747
rect 601 742 670 747
rect 713 742 1022 747
rect 1153 742 1270 747
rect 1313 742 1374 747
rect 1401 742 1470 747
rect 1713 742 1742 747
rect 1833 742 1854 747
rect 1897 742 2022 747
rect 2121 742 2206 747
rect 2289 742 2982 747
rect 3009 742 3070 747
rect 3081 742 3198 747
rect 3225 742 3430 747
rect 3609 742 3894 747
rect 3929 742 4006 747
rect 4249 742 4358 747
rect 289 712 294 742
rect 321 732 342 737
rect 361 732 430 737
rect 473 732 1070 737
rect 1273 732 1590 737
rect 1697 732 1750 737
rect 1761 732 1910 737
rect 2033 732 2254 737
rect 1089 727 1254 732
rect 2033 727 2038 732
rect 2289 727 2294 742
rect 2337 727 2430 732
rect 2449 727 2454 737
rect 2481 732 2558 737
rect 2577 732 2750 737
rect 2761 732 3062 737
rect 3089 732 3190 737
rect 3289 732 3334 737
rect 3393 732 3550 737
rect 3569 732 3742 737
rect 3569 727 3574 732
rect 3889 727 3894 742
rect 3905 732 3966 737
rect 4089 732 4206 737
rect 4089 727 4094 732
rect 529 722 614 727
rect 697 722 766 727
rect 785 722 1094 727
rect 1249 722 2038 727
rect 2185 722 2294 727
rect 2313 722 2342 727
rect 2425 722 2454 727
rect 2505 722 3294 727
rect 3441 722 3574 727
rect 3617 722 3862 727
rect 3889 722 4094 727
rect 4201 727 4206 732
rect 4249 727 4254 742
rect 4201 722 4254 727
rect 4353 727 4358 742
rect 4353 722 4374 727
rect 785 717 790 722
rect 3289 717 3446 722
rect 3617 717 3622 722
rect 321 712 374 717
rect 577 712 686 717
rect 761 712 790 717
rect 809 712 878 717
rect 937 712 1894 717
rect 681 707 766 712
rect 1889 707 1894 712
rect 2049 712 2646 717
rect 2665 712 2806 717
rect 2905 712 2966 717
rect 3017 712 3270 717
rect 3465 712 3622 717
rect 3689 712 3766 717
rect 3833 712 3926 717
rect 4265 712 4350 717
rect 4369 712 4374 722
rect 2049 707 2054 712
rect 2641 707 2646 712
rect 3945 707 4054 712
rect 521 702 598 707
rect 801 702 966 707
rect 1001 702 1198 707
rect 1241 702 1782 707
rect 1793 702 1854 707
rect 1889 702 2054 707
rect 2193 702 2286 707
rect 2313 702 2462 707
rect 2497 702 2526 707
rect 2553 702 2614 707
rect 2641 702 3134 707
rect 3225 702 3254 707
rect 3321 702 3950 707
rect 4049 702 4286 707
rect 1777 697 1782 702
rect 2609 697 2614 702
rect 3129 697 3230 702
rect 377 692 406 697
rect 569 692 718 697
rect 809 692 910 697
rect 945 692 1558 697
rect 1577 692 1750 697
rect 1777 692 1870 697
rect 2241 692 2374 697
rect 2537 692 2590 697
rect 2609 692 2670 697
rect 2753 692 2854 697
rect 2865 692 2910 697
rect 2921 692 3110 697
rect 3489 692 3734 697
rect 3817 692 4038 697
rect 2393 687 2518 692
rect 3729 687 3822 692
rect 4153 687 4222 692
rect 281 682 494 687
rect 529 682 566 687
rect 585 682 646 687
rect 769 682 854 687
rect 865 682 2198 687
rect 2209 682 2398 687
rect 2513 682 2766 687
rect 2777 682 2958 687
rect 2977 682 3070 687
rect 3113 682 3230 687
rect 3369 682 3470 687
rect 3489 682 3710 687
rect 3841 682 4158 687
rect 4217 682 4294 687
rect 345 672 462 677
rect 513 672 550 677
rect 801 672 934 677
rect 985 672 1366 677
rect 1377 672 1534 677
rect 1553 672 1654 677
rect 1745 672 1822 677
rect 1881 672 1902 677
rect 1921 667 2022 672
rect 241 662 438 667
rect 489 662 582 667
rect 665 662 686 667
rect 921 662 950 667
rect 1281 662 1926 667
rect 2017 662 2046 667
rect 2065 662 2134 667
rect 993 657 1086 662
rect 1161 657 1262 662
rect 2065 657 2070 662
rect 169 652 342 657
rect 593 652 758 657
rect 777 652 798 657
rect 881 652 918 657
rect 969 652 998 657
rect 1081 652 1110 657
rect 1137 652 1166 657
rect 1257 652 1582 657
rect 1729 652 2070 657
rect 2129 657 2134 662
rect 2193 657 2198 682
rect 3369 677 3374 682
rect 2241 672 2406 677
rect 2457 672 2838 677
rect 2849 672 2998 677
rect 3041 672 3086 677
rect 3097 672 3150 677
rect 3345 672 3374 677
rect 3465 677 3470 682
rect 3465 672 4030 677
rect 4177 672 4206 677
rect 4025 667 4182 672
rect 2249 662 3030 667
rect 3345 662 3606 667
rect 3785 662 3878 667
rect 3105 657 3214 662
rect 3345 657 3350 662
rect 3601 657 3790 662
rect 3897 657 4006 662
rect 2129 652 2158 657
rect 2193 652 2678 657
rect 2745 652 2846 657
rect 2889 652 2966 657
rect 2985 652 3110 657
rect 3209 652 3350 657
rect 3457 652 3582 657
rect 3809 652 3902 657
rect 4001 652 4110 657
rect 337 647 598 652
rect 881 647 886 652
rect 177 642 302 647
rect 689 642 886 647
rect 961 642 1118 647
rect 689 637 694 642
rect 1137 637 1142 652
rect 1577 647 1734 652
rect 305 632 342 637
rect 369 632 478 637
rect 537 632 694 637
rect 785 632 830 637
rect 849 632 1142 637
rect 1153 642 1558 647
rect 1753 642 1806 647
rect 1817 642 2582 647
rect 2673 642 2902 647
rect 2913 642 3038 647
rect 3065 642 3198 647
rect 3401 642 3678 647
rect 3697 642 3806 647
rect 3857 642 3990 647
rect 4057 642 4126 647
rect 1153 627 1158 642
rect 2673 637 2678 642
rect 1169 632 1238 637
rect 1305 632 1982 637
rect 2017 632 2054 637
rect 2113 632 2206 637
rect 2305 632 2678 637
rect 2689 632 3294 637
rect 3385 632 3534 637
rect 3681 632 3750 637
rect 3953 632 3982 637
rect 2689 627 2694 632
rect 3681 627 3686 632
rect 3745 627 3958 632
rect 185 622 262 627
rect 305 617 310 627
rect 393 622 598 627
rect 737 622 846 627
rect 945 622 1158 627
rect 1241 622 1326 627
rect 1345 622 1582 627
rect 1649 622 2446 627
rect 2553 622 2694 627
rect 2705 622 2790 627
rect 2873 622 3062 627
rect 3441 622 3686 627
rect 3705 622 3726 627
rect 4073 622 4126 627
rect 945 617 950 622
rect 2441 617 2558 622
rect 3081 617 3406 622
rect 233 612 310 617
rect 505 612 718 617
rect 753 612 782 617
rect 825 612 950 617
rect 1289 612 1374 617
rect 1625 612 1750 617
rect 1937 612 2030 617
rect 2153 612 2246 617
rect 2265 612 2422 617
rect 329 607 486 612
rect 969 607 1070 612
rect 1761 607 1942 612
rect 2241 607 2246 612
rect 2577 607 2582 617
rect 2593 612 2638 617
rect 2721 612 3086 617
rect 3401 612 3630 617
rect 3729 612 3846 617
rect 3953 612 4102 617
rect 3729 607 3734 612
rect 121 602 334 607
rect 481 602 678 607
rect 673 597 678 602
rect 705 602 846 607
rect 929 602 974 607
rect 1065 602 1766 607
rect 1961 602 2022 607
rect 2049 602 2134 607
rect 2177 602 2214 607
rect 2241 602 2326 607
rect 2401 602 2454 607
rect 2481 602 3318 607
rect 3345 602 3390 607
rect 3449 602 3734 607
rect 3817 602 4342 607
rect 705 597 710 602
rect 2017 597 2022 602
rect 2321 597 2326 602
rect 137 592 214 597
rect 305 592 470 597
rect 489 592 622 597
rect 649 592 710 597
rect 721 592 830 597
rect 977 592 1046 597
rect 1089 592 1166 597
rect 1193 592 1262 597
rect 1297 592 1350 597
rect 1433 592 1494 597
rect 1577 592 1974 597
rect 2017 592 2038 597
rect 2177 592 2246 597
rect 2281 592 2302 597
rect 2321 592 2598 597
rect 2673 592 3238 597
rect 3297 592 3742 597
rect 3785 592 3870 597
rect 3953 592 3990 597
rect 4001 592 4102 597
rect 4153 592 4230 597
rect 465 587 470 592
rect 265 582 294 587
rect 385 582 446 587
rect 465 582 566 587
rect 681 582 838 587
rect 1081 582 1270 587
rect 1361 582 1462 587
rect 1473 582 1798 587
rect 1833 582 1878 587
rect 1953 582 2062 587
rect 2249 582 2318 587
rect 2329 582 2454 587
rect 2505 582 2806 587
rect 2825 582 2870 587
rect 2881 582 2950 587
rect 2961 582 2998 587
rect 3033 582 3126 587
rect 3193 582 3222 587
rect 3241 582 3326 587
rect 3361 582 3750 587
rect 3953 582 3998 587
rect 289 577 390 582
rect 561 577 686 582
rect 1473 577 1478 582
rect 2113 577 2230 582
rect 3217 577 3222 582
rect 409 572 542 577
rect 705 572 750 577
rect 857 572 958 577
rect 1001 572 1038 577
rect 1081 572 1110 577
rect 1129 572 1198 577
rect 1241 572 1310 577
rect 1417 572 1478 577
rect 1537 572 2118 577
rect 2225 572 2926 577
rect 2977 572 3078 577
rect 3217 572 3254 577
rect 3337 572 3774 577
rect 3969 572 4022 577
rect 4113 572 4198 577
rect 769 567 862 572
rect 953 567 958 572
rect 1537 567 1542 572
rect 249 562 270 567
rect 377 562 430 567
rect 457 562 542 567
rect 625 562 774 567
rect 953 562 1542 567
rect 1553 562 2046 567
rect 2041 557 2046 562
rect 2129 562 2486 567
rect 2593 562 2710 567
rect 2729 562 2798 567
rect 2809 562 2910 567
rect 2921 562 2926 572
rect 3217 562 3310 567
rect 3361 562 3390 567
rect 3417 562 3470 567
rect 3505 562 3574 567
rect 4121 562 4310 567
rect 2129 557 2134 562
rect 2497 557 2598 562
rect 2705 557 2710 562
rect 2945 557 3126 562
rect 193 552 918 557
rect 945 552 966 557
rect 1001 552 1062 557
rect 1105 552 1158 557
rect 1193 552 1406 557
rect 1537 552 1590 557
rect 1617 552 1646 557
rect 1745 552 1878 557
rect 1937 552 2022 557
rect 2041 552 2134 557
rect 2201 552 2278 557
rect 2353 552 2438 557
rect 913 547 918 552
rect 1401 547 1542 552
rect 1585 547 1590 552
rect 2497 547 2502 557
rect 2617 552 2662 557
rect 2705 552 2950 557
rect 3121 552 3478 557
rect 3625 552 3686 557
rect 3937 552 3974 557
rect 4153 552 4318 557
rect 225 542 246 547
rect 345 542 390 547
rect 473 542 598 547
rect 777 542 854 547
rect 913 542 942 547
rect 225 537 230 542
rect 937 537 942 542
rect 1049 542 1358 547
rect 1585 542 1638 547
rect 1681 542 1774 547
rect 1793 542 1814 547
rect 2153 542 2302 547
rect 2425 542 2502 547
rect 2545 542 2966 547
rect 3009 542 3110 547
rect 3233 542 3582 547
rect 3617 542 3662 547
rect 3905 542 3950 547
rect 1049 537 1054 542
rect 2545 537 2550 542
rect 3969 537 3974 552
rect 4089 542 4198 547
rect 4225 542 4318 547
rect 193 532 230 537
rect 377 532 462 537
rect 521 532 550 537
rect 617 532 766 537
rect 937 532 1054 537
rect 1073 532 1118 537
rect 1137 532 1334 537
rect 1473 532 1582 537
rect 1609 532 1798 537
rect 1929 532 1974 537
rect 2345 532 2430 537
rect 2529 532 2550 537
rect 2593 532 2646 537
rect 457 527 526 532
rect 1969 527 1974 532
rect 2217 527 2326 532
rect 2529 527 2534 532
rect 569 522 734 527
rect 833 522 910 527
rect 1097 522 1198 527
rect 1361 522 1454 527
rect 1641 522 1958 527
rect 1969 522 2182 527
rect 2193 522 2222 527
rect 2321 522 2382 527
rect 2417 522 2534 527
rect 1001 517 1078 522
rect 1953 517 1958 522
rect 2177 517 2182 522
rect 2641 517 2646 532
rect 2665 527 2670 537
rect 2713 532 2838 537
rect 3001 532 3118 537
rect 3193 532 3398 537
rect 3585 532 3614 537
rect 3657 532 3774 537
rect 3873 532 3942 537
rect 3969 532 4070 537
rect 2865 527 2982 532
rect 2665 522 2726 527
rect 2745 522 2806 527
rect 2841 522 2870 527
rect 2977 522 3030 527
rect 3249 522 3374 527
rect 3393 522 3398 532
rect 4065 527 4070 532
rect 3529 522 3798 527
rect 4065 522 4118 527
rect 145 512 246 517
rect 417 512 502 517
rect 513 512 830 517
rect 513 507 518 512
rect 825 507 830 512
rect 921 512 1006 517
rect 1073 512 1310 517
rect 1433 512 1534 517
rect 1609 512 1702 517
rect 1721 512 1830 517
rect 1953 512 1990 517
rect 2177 512 2566 517
rect 2577 512 2622 517
rect 2641 512 2814 517
rect 2857 512 2902 517
rect 2937 512 2958 517
rect 2977 512 3062 517
rect 3209 512 3294 517
rect 3337 512 3470 517
rect 3513 512 3550 517
rect 3609 512 3766 517
rect 3865 512 3902 517
rect 3961 512 4086 517
rect 4257 512 4374 517
rect 921 507 926 512
rect 2561 507 2566 512
rect 217 502 342 507
rect 433 502 542 507
rect 553 502 582 507
rect 665 502 702 507
rect 825 502 926 507
rect 1017 502 1126 507
rect 1161 502 1622 507
rect 1633 502 1958 507
rect 2209 502 2238 507
rect 577 497 670 502
rect 1617 497 1622 502
rect 2233 497 2238 502
rect 2313 502 2342 507
rect 2393 502 2478 507
rect 2561 502 2774 507
rect 2785 502 2814 507
rect 2897 502 3022 507
rect 3041 502 3158 507
rect 3201 502 3238 507
rect 3297 502 3638 507
rect 3665 502 3966 507
rect 4081 502 4142 507
rect 4313 502 4358 507
rect 2313 497 2318 502
rect 321 492 406 497
rect 401 487 406 492
rect 689 492 806 497
rect 1025 492 1086 497
rect 1193 492 1214 497
rect 1257 492 1310 497
rect 1481 492 1550 497
rect 1617 492 1654 497
rect 1809 492 1902 497
rect 1945 492 2078 497
rect 2233 492 2318 497
rect 689 487 694 492
rect 1649 487 1814 492
rect 401 482 694 487
rect 865 482 902 487
rect 1121 482 1390 487
rect 1505 482 1630 487
rect 737 477 846 482
rect 921 477 1102 482
rect 2337 477 2342 502
rect 2369 492 2454 497
rect 2505 492 2686 497
rect 2713 492 2742 497
rect 2769 487 2774 502
rect 2809 497 2902 502
rect 3201 497 3206 502
rect 2921 492 3206 497
rect 3225 492 3390 497
rect 3409 492 3494 497
rect 3505 492 3670 497
rect 3777 492 3918 497
rect 3977 492 4014 497
rect 3505 487 3510 492
rect 3665 487 3758 492
rect 2353 482 2494 487
rect 2569 482 2606 487
rect 2769 482 3510 487
rect 3753 482 3822 487
rect 3529 477 3646 482
rect 713 472 742 477
rect 841 472 926 477
rect 1097 472 1774 477
rect 1769 467 1774 472
rect 2089 472 2310 477
rect 2337 472 2462 477
rect 2697 472 2766 477
rect 2865 472 3062 477
rect 3497 472 3534 477
rect 3641 472 3910 477
rect 3929 472 4206 477
rect 2089 467 2094 472
rect 3057 467 3502 472
rect 3929 467 3934 472
rect 521 462 694 467
rect 729 462 1750 467
rect 1769 462 2094 467
rect 2273 462 2414 467
rect 2449 462 2510 467
rect 2529 462 2694 467
rect 2769 462 2798 467
rect 2905 462 3038 467
rect 3521 462 3638 467
rect 3729 462 3934 467
rect 4201 467 4206 472
rect 4201 462 4246 467
rect 521 457 526 462
rect 297 452 382 457
rect 497 452 526 457
rect 689 457 694 462
rect 2529 457 2534 462
rect 689 452 1214 457
rect 1233 452 1606 457
rect 2513 452 2534 457
rect 2641 452 3414 457
rect 3449 452 3550 457
rect 3665 452 3702 457
rect 3753 452 4190 457
rect 2249 447 2518 452
rect 2641 447 2646 452
rect 465 442 1734 447
rect 2225 442 2254 447
rect 2529 442 2558 447
rect 2593 442 2646 447
rect 2769 442 2974 447
rect 3385 442 3894 447
rect 225 432 502 437
rect 697 432 734 437
rect 1033 432 1942 437
rect 753 427 1006 432
rect 2225 427 2230 442
rect 2769 437 2774 442
rect 3889 437 3894 442
rect 3977 442 4102 447
rect 3977 437 3982 442
rect 2265 432 2774 437
rect 2809 432 2878 437
rect 2889 432 2950 437
rect 3185 432 3270 437
rect 3321 432 3406 437
rect 3513 432 3558 437
rect 3737 432 3758 437
rect 3801 432 3870 437
rect 3889 432 3982 437
rect 4001 432 4062 437
rect 4145 432 4182 437
rect 3185 427 3190 432
rect 185 422 462 427
rect 681 422 758 427
rect 1001 422 1030 427
rect 1129 422 1446 427
rect 1529 422 2230 427
rect 2249 422 2790 427
rect 2817 422 2838 427
rect 2865 422 2926 427
rect 2937 422 3030 427
rect 3049 422 3142 427
rect 3161 422 3190 427
rect 3265 427 3270 432
rect 3553 427 3718 432
rect 3265 422 3366 427
rect 3457 422 3534 427
rect 3713 422 3830 427
rect 4025 422 4238 427
rect 4257 422 4374 427
rect 1025 417 1030 422
rect 1441 417 1534 422
rect 2817 417 2822 422
rect 3049 417 3054 422
rect 169 412 278 417
rect 369 412 398 417
rect 393 407 398 412
rect 465 412 1014 417
rect 1025 412 1422 417
rect 1553 412 1886 417
rect 2225 412 2270 417
rect 2305 412 2414 417
rect 2537 412 2614 417
rect 2633 412 3054 417
rect 3137 417 3142 422
rect 3137 412 3254 417
rect 3345 412 3798 417
rect 3937 412 4198 417
rect 465 407 470 412
rect 1553 407 1558 412
rect 2409 407 2542 412
rect 2609 407 2614 412
rect 145 402 182 407
rect 393 402 470 407
rect 753 402 846 407
rect 1305 402 1342 407
rect 1385 402 1558 407
rect 1569 402 1662 407
rect 1785 402 1814 407
rect 1905 402 1942 407
rect 2217 402 2390 407
rect 2561 402 2582 407
rect 2609 402 2790 407
rect 2801 402 2862 407
rect 2873 402 3326 407
rect 3353 402 4062 407
rect 4169 402 4270 407
rect 177 397 182 402
rect 609 397 734 402
rect 865 397 1030 402
rect 1169 397 1286 402
rect 1809 397 1910 402
rect 2561 397 2566 402
rect 177 392 214 397
rect 249 392 286 397
rect 585 392 614 397
rect 729 392 870 397
rect 1025 392 1054 397
rect 1145 392 1174 397
rect 1281 392 1670 397
rect 1929 392 2022 397
rect 2145 392 2246 397
rect 2305 392 2382 397
rect 2401 392 2502 397
rect 2521 392 2566 397
rect 2785 397 2790 402
rect 2785 392 2870 397
rect 2881 392 2934 397
rect 2969 392 3086 397
rect 3369 392 3806 397
rect 3985 392 4046 397
rect 4225 392 4310 397
rect 2561 387 2766 392
rect 3161 387 3246 392
rect 249 382 318 387
rect 489 382 542 387
rect 617 382 710 387
rect 721 382 1046 387
rect 1057 382 1166 387
rect 1209 382 1278 387
rect 1289 382 1422 387
rect 1705 382 1774 387
rect 1825 382 1846 387
rect 2281 382 2342 387
rect 2353 382 2462 387
rect 2497 382 2550 387
rect 2761 382 3166 387
rect 3241 382 3406 387
rect 3497 382 3526 387
rect 3561 382 3646 387
rect 3681 382 3710 387
rect 3729 382 4158 387
rect 721 377 726 382
rect 1705 377 1710 382
rect 97 372 238 377
rect 233 367 238 372
rect 329 372 478 377
rect 329 367 334 372
rect 233 362 334 367
rect 473 367 478 372
rect 553 372 606 377
rect 553 367 558 372
rect 473 362 558 367
rect 601 367 606 372
rect 697 372 726 377
rect 777 372 822 377
rect 937 372 974 377
rect 1153 372 1294 377
rect 1305 372 1358 377
rect 1497 372 1558 377
rect 1681 372 1710 377
rect 1769 377 1774 382
rect 3401 377 3502 382
rect 4153 377 4158 382
rect 4257 382 4326 387
rect 4257 377 4262 382
rect 1769 372 1798 377
rect 1873 372 2054 377
rect 697 367 702 372
rect 1385 367 1478 372
rect 1873 367 1878 372
rect 601 362 702 367
rect 1041 362 1270 367
rect 1369 362 1390 367
rect 1473 362 1742 367
rect 1809 362 1878 367
rect 2049 367 2054 372
rect 2321 372 2886 377
rect 2921 372 2950 377
rect 3177 372 3230 377
rect 3529 372 3862 377
rect 3969 372 4134 377
rect 4153 372 4262 377
rect 4281 372 4366 377
rect 2321 367 2326 372
rect 2945 367 3182 372
rect 3225 367 3382 372
rect 3529 367 3534 372
rect 2049 362 2126 367
rect 2225 362 2342 367
rect 2433 362 2822 367
rect 3377 362 3534 367
rect 3553 362 3774 367
rect 3785 362 3894 367
rect 1041 357 1046 362
rect 1265 357 1374 362
rect 1737 357 1814 362
rect 1913 357 2014 362
rect 2817 357 2918 362
rect 721 352 814 357
rect 977 352 1046 357
rect 1097 352 1158 357
rect 1401 352 1502 357
rect 1889 352 1918 357
rect 2009 352 2038 357
rect 2249 352 2550 357
rect 2577 352 2678 357
rect 2721 352 2774 357
rect 2913 352 2942 357
rect 2993 352 3118 357
rect 3177 352 3358 357
rect 3593 352 3854 357
rect 1545 347 1718 352
rect 1889 347 1894 352
rect 185 342 310 347
rect 329 342 406 347
rect 529 342 590 347
rect 617 342 662 347
rect 801 342 846 347
rect 1025 342 1134 347
rect 1241 342 1334 347
rect 1521 342 1550 347
rect 1713 342 1894 347
rect 1905 342 2014 347
rect 2145 342 2310 347
rect 2449 342 3366 347
rect 3417 342 3558 347
rect 3577 342 3614 347
rect 3633 342 3750 347
rect 3769 342 3814 347
rect 3993 342 4078 347
rect 1889 337 1894 342
rect 2449 337 2454 342
rect 3553 337 3558 342
rect 201 332 534 337
rect 529 327 534 332
rect 641 332 1678 337
rect 1889 332 1918 337
rect 1953 332 2070 337
rect 2345 332 2454 337
rect 2465 332 2526 337
rect 641 327 646 332
rect 1673 327 1678 332
rect 305 322 390 327
rect 457 322 510 327
rect 529 322 646 327
rect 665 322 750 327
rect 809 322 862 327
rect 1297 322 1430 327
rect 1569 322 1654 327
rect 1673 322 1846 327
rect 2217 322 2262 327
rect 2497 322 2502 332
rect 2521 327 2526 332
rect 2593 332 2654 337
rect 2681 332 2750 337
rect 2977 332 3062 337
rect 3185 332 3270 337
rect 3393 332 3462 337
rect 3553 332 3630 337
rect 3657 332 3734 337
rect 2593 327 2598 332
rect 2769 327 2950 332
rect 2521 322 2598 327
rect 2649 322 2774 327
rect 2945 322 3126 327
rect 3225 322 3294 327
rect 1169 317 1278 322
rect 1449 317 1550 322
rect 1841 317 1846 322
rect 3729 317 3734 332
rect 3745 327 3750 342
rect 3809 337 3814 342
rect 3809 332 3854 337
rect 3913 332 4022 337
rect 4113 332 4246 337
rect 3745 322 3950 327
rect 793 312 1174 317
rect 1273 312 1454 317
rect 1545 312 1598 317
rect 1841 312 1886 317
rect 2721 312 2918 317
rect 2937 312 2998 317
rect 3337 312 3414 317
rect 3537 312 3718 317
rect 3729 312 4006 317
rect 4265 312 4326 317
rect 2913 307 2918 312
rect 553 302 726 307
rect 777 302 806 307
rect 1185 302 1382 307
rect 1417 302 1454 307
rect 1505 302 1710 307
rect 1793 302 1878 307
rect 1969 302 2198 307
rect 2225 302 2326 307
rect 2345 302 2478 307
rect 2593 302 2630 307
rect 2697 302 2830 307
rect 2913 302 3142 307
rect 1793 297 1798 302
rect 1969 297 1974 302
rect 609 292 638 297
rect 633 277 638 292
rect 793 292 846 297
rect 793 277 798 292
rect 265 272 294 277
rect 633 272 798 277
rect 841 277 846 292
rect 1017 292 1350 297
rect 1401 292 1598 297
rect 1017 277 1022 292
rect 1593 287 1598 292
rect 1665 292 1798 297
rect 1809 292 1838 297
rect 1665 287 1670 292
rect 1041 282 1070 287
rect 841 272 1022 277
rect 1065 277 1070 282
rect 1545 282 1574 287
rect 1593 282 1670 287
rect 1833 287 1838 292
rect 1897 292 1974 297
rect 2193 297 2198 302
rect 2345 297 2350 302
rect 2193 292 2350 297
rect 2473 297 2478 302
rect 3409 297 3414 312
rect 3825 302 3958 307
rect 2473 292 3102 297
rect 3409 292 3454 297
rect 1897 287 1902 292
rect 1833 282 1902 287
rect 1985 282 2358 287
rect 2649 282 2710 287
rect 2817 282 2870 287
rect 2953 282 3094 287
rect 3313 282 3390 287
rect 3561 282 3614 287
rect 1545 277 1550 282
rect 2473 277 2582 282
rect 2865 277 2958 282
rect 3313 277 3318 282
rect 1065 272 1550 277
rect 2289 272 2478 277
rect 2577 272 2606 277
rect 3121 272 3270 277
rect 3289 272 3318 277
rect 3385 277 3390 282
rect 3385 272 3590 277
rect 3785 272 3886 277
rect 2129 267 2262 272
rect 2625 267 2846 272
rect 3121 267 3126 272
rect 1969 262 1998 267
rect 1993 257 1998 262
rect 2105 262 2134 267
rect 2257 262 2278 267
rect 2489 262 2518 267
rect 2537 262 2630 267
rect 2841 262 3126 267
rect 3265 267 3270 272
rect 3785 267 3790 272
rect 3265 262 3334 267
rect 2105 257 2110 262
rect 2273 257 2494 262
rect 3329 257 3334 262
rect 3457 262 3486 267
rect 3673 262 3742 267
rect 3761 262 3790 267
rect 3881 267 3886 272
rect 3881 262 3910 267
rect 3977 262 4102 267
rect 3457 257 3462 262
rect 3673 257 3678 262
rect 497 252 582 257
rect 497 247 502 252
rect 145 242 214 247
rect 393 242 502 247
rect 577 247 582 252
rect 921 252 1118 257
rect 577 242 614 247
rect 761 242 830 247
rect 921 237 926 252
rect 441 232 566 237
rect 897 232 926 237
rect 1113 237 1118 252
rect 1153 252 1374 257
rect 1993 252 2110 257
rect 2129 252 2246 257
rect 2601 252 2830 257
rect 3137 252 3310 257
rect 3329 252 3462 257
rect 3617 252 3678 257
rect 3737 257 3742 262
rect 3977 257 3982 262
rect 3737 252 3862 257
rect 3881 252 3982 257
rect 4097 257 4102 262
rect 4097 252 4126 257
rect 4193 252 4246 257
rect 1153 237 1158 252
rect 1369 247 1374 252
rect 2825 247 3142 252
rect 1369 242 1454 247
rect 2313 242 2694 247
rect 1201 237 1350 242
rect 2689 237 2806 242
rect 3209 237 3286 242
rect 3857 237 3862 252
rect 3929 242 4174 247
rect 1113 232 1158 237
rect 1177 232 1206 237
rect 1345 232 1486 237
rect 2225 232 2294 237
rect 2801 232 2830 237
rect 2921 232 3054 237
rect 801 227 878 232
rect 2225 227 2230 232
rect 193 222 374 227
rect 401 222 486 227
rect 617 222 702 227
rect 617 217 622 222
rect 305 212 422 217
rect 457 212 622 217
rect 697 217 702 222
rect 737 222 806 227
rect 873 222 998 227
rect 1073 222 1134 227
rect 1217 222 1390 227
rect 1441 222 1478 227
rect 737 217 742 222
rect 993 217 998 222
rect 1537 217 1542 227
rect 1561 222 1638 227
rect 1561 217 1566 222
rect 697 212 742 217
rect 817 212 894 217
rect 993 212 1254 217
rect 1337 212 1566 217
rect 1633 217 1638 222
rect 1785 222 1854 227
rect 2201 222 2230 227
rect 2289 227 2294 232
rect 2921 227 2926 232
rect 2289 222 2398 227
rect 2625 222 2774 227
rect 2809 222 2926 227
rect 3049 227 3054 232
rect 3089 232 3214 237
rect 3281 232 3310 237
rect 3689 232 3774 237
rect 3857 232 3926 237
rect 4009 232 4238 237
rect 3089 227 3094 232
rect 3921 227 4014 232
rect 3049 222 3094 227
rect 3225 222 3326 227
rect 3377 222 3678 227
rect 3753 222 3782 227
rect 3825 222 3902 227
rect 4153 222 4310 227
rect 1785 217 1790 222
rect 1633 212 1790 217
rect 1849 217 1854 222
rect 2625 217 2630 222
rect 3673 217 3758 222
rect 4033 217 4158 222
rect 1849 212 1878 217
rect 2217 212 2342 217
rect 2409 212 2630 217
rect 2865 212 2934 217
rect 2993 212 3070 217
rect 3817 212 4038 217
rect 305 207 310 212
rect 2337 207 2414 212
rect 2865 207 2870 212
rect 2929 207 2934 212
rect 217 202 310 207
rect 321 202 902 207
rect 937 202 1006 207
rect 1025 202 1110 207
rect 1377 202 1702 207
rect 1697 197 1702 202
rect 1785 202 1910 207
rect 1953 202 2062 207
rect 2249 202 2318 207
rect 2609 202 2870 207
rect 1785 197 1790 202
rect 2913 197 2918 207
rect 2929 202 3038 207
rect 3049 202 3110 207
rect 3321 202 3374 207
rect 3745 202 3870 207
rect 249 192 278 197
rect 273 177 278 192
rect 505 192 566 197
rect 505 187 510 192
rect 425 182 510 187
rect 561 187 566 192
rect 785 192 838 197
rect 785 187 790 192
rect 561 182 790 187
rect 833 187 838 192
rect 1121 192 1206 197
rect 1297 192 1374 197
rect 1417 192 1462 197
rect 1697 192 1790 197
rect 1897 192 2006 197
rect 2137 192 2310 197
rect 2353 192 2470 197
rect 2545 192 2918 197
rect 3009 197 3014 202
rect 3865 197 3870 202
rect 3961 202 4222 207
rect 3961 197 3966 202
rect 3009 192 3174 197
rect 3793 192 3846 197
rect 3865 192 3966 197
rect 4225 192 4302 197
rect 1121 187 1126 192
rect 833 182 1126 187
rect 425 177 430 182
rect 273 172 430 177
rect 1201 177 1206 192
rect 1217 182 1334 187
rect 1481 182 1662 187
rect 3297 182 3398 187
rect 4033 182 4118 187
rect 1353 177 1486 182
rect 1657 177 1662 182
rect 2697 177 2790 182
rect 3137 177 3222 182
rect 1201 172 1358 177
rect 1657 172 1878 177
rect 2257 172 2350 177
rect 2257 167 2262 172
rect 529 162 686 167
rect 1081 162 1174 167
rect 1329 162 1702 167
rect 1193 157 1334 162
rect 1697 157 1702 162
rect 1761 162 1790 167
rect 1969 162 2038 167
rect 2225 162 2262 167
rect 2345 167 2350 172
rect 2673 172 2702 177
rect 2785 172 3142 177
rect 3217 172 3286 177
rect 3377 172 3406 177
rect 3425 172 3662 177
rect 2673 167 2678 172
rect 3281 167 3382 172
rect 2345 162 2678 167
rect 2697 162 2774 167
rect 3153 162 3206 167
rect 1761 157 1766 162
rect 1969 157 1974 162
rect 449 152 1070 157
rect 449 147 454 152
rect 1065 147 1070 152
rect 1153 152 1198 157
rect 1537 152 1654 157
rect 1697 152 1766 157
rect 1945 152 1974 157
rect 2033 157 2038 162
rect 3425 157 3430 172
rect 2033 152 2062 157
rect 2273 152 2334 157
rect 2793 152 3430 157
rect 3657 157 3662 172
rect 3681 172 3766 177
rect 3681 157 3686 172
rect 3761 167 3766 172
rect 3761 162 3782 167
rect 3777 157 3782 162
rect 3657 152 3686 157
rect 3705 152 3766 157
rect 3777 152 4142 157
rect 1153 147 1158 152
rect 169 142 454 147
rect 473 142 550 147
rect 641 142 718 147
rect 1065 142 1158 147
rect 1177 142 1198 147
rect 1217 142 1326 147
rect 1409 142 1462 147
rect 1497 142 1598 147
rect 1905 142 2006 147
rect 2025 142 2262 147
rect 2345 142 2542 147
rect 2689 142 2806 147
rect 2257 137 2350 142
rect 1329 132 1510 137
rect 2801 127 2806 142
rect 2985 142 3038 147
rect 2985 127 2990 142
rect 305 122 334 127
rect 329 117 334 122
rect 561 122 1166 127
rect 561 117 566 122
rect 1161 117 1166 122
rect 1273 122 1574 127
rect 1977 122 2006 127
rect 1273 117 1278 122
rect 2001 117 2006 122
rect 2065 122 2118 127
rect 2065 117 2070 122
rect 329 112 566 117
rect 625 112 662 117
rect 1161 112 1278 117
rect 1297 112 1470 117
rect 2001 112 2070 117
rect 2113 117 2118 122
rect 2201 122 2254 127
rect 2201 117 2206 122
rect 2113 112 2206 117
rect 2249 117 2254 122
rect 2329 122 2358 127
rect 2433 122 2510 127
rect 2553 122 2694 127
rect 2801 122 2990 127
rect 3033 127 3038 142
rect 3209 142 3262 147
rect 3209 127 3214 142
rect 3033 122 3214 127
rect 3257 127 3262 142
rect 3433 142 3686 147
rect 3993 142 4062 147
rect 4105 142 4222 147
rect 4241 142 4358 147
rect 3433 127 3438 142
rect 3257 122 3438 127
rect 3457 122 3486 127
rect 2329 117 2334 122
rect 2433 117 2438 122
rect 2249 112 2334 117
rect 2401 112 2438 117
rect 3481 117 3486 122
rect 3697 122 3982 127
rect 3697 117 3702 122
rect 3481 112 3702 117
rect 3977 117 3982 122
rect 4041 122 4094 127
rect 4041 117 4046 122
rect 3977 112 4046 117
rect 4089 107 4094 122
rect 4249 122 4278 127
rect 4249 107 4254 122
rect 609 102 774 107
rect 4089 102 4254 107
rect 1281 82 3870 87
rect 1601 62 1630 67
rect 1625 57 1630 62
rect 2153 62 2182 67
rect 2153 57 2158 62
rect 1625 52 2158 57
use AND2X2  AND2X2_0
timestamp 1745462530
transform 1 0 2544 0 1 3570
box -8 -3 40 105
use AND2X2  AND2X2_1
timestamp 1745462530
transform 1 0 2536 0 -1 3770
box -8 -3 40 105
use AND2X2  AND2X2_2
timestamp 1745462530
transform 1 0 2632 0 1 3570
box -8 -3 40 105
use AND2X2  AND2X2_3
timestamp 1745462530
transform 1 0 2576 0 -1 3770
box -8 -3 40 105
use AND2X2  AND2X2_4
timestamp 1745462530
transform 1 0 2616 0 -1 3770
box -8 -3 40 105
use AND2X2  AND2X2_5
timestamp 1745462530
transform 1 0 1864 0 1 3570
box -8 -3 40 105
use AND2X2  AND2X2_6
timestamp 1745462530
transform 1 0 2656 0 -1 3770
box -8 -3 40 105
use AND2X2  AND2X2_7
timestamp 1745462530
transform 1 0 1768 0 1 3570
box -8 -3 40 105
use AND2X2  AND2X2_8
timestamp 1745462530
transform 1 0 2496 0 -1 2570
box -8 -3 40 105
use AND2X2  AND2X2_9
timestamp 1745462530
transform 1 0 2464 0 1 2570
box -8 -3 40 105
use AND2X2  AND2X2_10
timestamp 1745462530
transform 1 0 1600 0 -1 3570
box -8 -3 40 105
use AND2X2  AND2X2_11
timestamp 1745462530
transform 1 0 3760 0 1 2170
box -8 -3 40 105
use AND2X2  AND2X2_12
timestamp 1745462530
transform 1 0 3000 0 1 1570
box -8 -3 40 105
use AND2X2  AND2X2_13
timestamp 1745462530
transform 1 0 3056 0 1 1570
box -8 -3 40 105
use AND2X2  AND2X2_14
timestamp 1745462530
transform 1 0 3552 0 -1 1770
box -8 -3 40 105
use AND2X2  AND2X2_15
timestamp 1745462530
transform 1 0 3200 0 -1 2170
box -8 -3 40 105
use AND2X2  AND2X2_16
timestamp 1745462530
transform 1 0 3112 0 -1 2170
box -8 -3 40 105
use AND2X2  AND2X2_17
timestamp 1745462530
transform 1 0 2016 0 1 2970
box -8 -3 40 105
use AND2X2  AND2X2_18
timestamp 1745462530
transform 1 0 384 0 1 3970
box -8 -3 40 105
use AND2X2  AND2X2_19
timestamp 1745462530
transform 1 0 1832 0 -1 4170
box -8 -3 40 105
use AND2X2  AND2X2_20
timestamp 1745462530
transform 1 0 1880 0 1 4170
box -8 -3 40 105
use AND2X2  AND2X2_21
timestamp 1745462530
transform 1 0 4008 0 -1 4170
box -8 -3 40 105
use AND2X2  AND2X2_22
timestamp 1745462530
transform 1 0 4032 0 -1 3970
box -8 -3 40 105
use AND2X2  AND2X2_23
timestamp 1745462530
transform 1 0 4128 0 1 4170
box -8 -3 40 105
use AND2X2  AND2X2_24
timestamp 1745462530
transform 1 0 4048 0 1 3970
box -8 -3 40 105
use AND2X2  AND2X2_25
timestamp 1745462530
transform 1 0 2848 0 1 4170
box -8 -3 40 105
use AND2X2  AND2X2_26
timestamp 1745462530
transform 1 0 776 0 1 3770
box -8 -3 40 105
use AND2X2  AND2X2_27
timestamp 1745462530
transform 1 0 2528 0 1 4170
box -8 -3 40 105
use AND2X2  AND2X2_28
timestamp 1745462530
transform 1 0 1200 0 1 3970
box -8 -3 40 105
use AND2X2  AND2X2_29
timestamp 1745462530
transform 1 0 1248 0 1 3970
box -8 -3 40 105
use AOI21X1  AOI21X1_0
timestamp 1745462530
transform 1 0 2336 0 1 2570
box -7 -3 39 105
use AOI21X1  AOI21X1_1
timestamp 1745462530
transform 1 0 320 0 1 3570
box -7 -3 39 105
use AOI21X1  AOI21X1_2
timestamp 1745462530
transform 1 0 248 0 1 3570
box -7 -3 39 105
use AOI21X1  AOI21X1_3
timestamp 1745462530
transform 1 0 176 0 -1 3570
box -7 -3 39 105
use AOI21X1  AOI21X1_4
timestamp 1745462530
transform 1 0 224 0 -1 3570
box -7 -3 39 105
use AOI21X1  AOI21X1_5
timestamp 1745462530
transform 1 0 2480 0 -1 1770
box -7 -3 39 105
use AOI21X1  AOI21X1_6
timestamp 1745462530
transform 1 0 2496 0 1 1570
box -7 -3 39 105
use AOI21X1  AOI21X1_7
timestamp 1745462530
transform 1 0 2424 0 -1 1770
box -7 -3 39 105
use AOI21X1  AOI21X1_8
timestamp 1745462530
transform 1 0 2424 0 1 1570
box -7 -3 39 105
use AOI21X1  AOI21X1_9
timestamp 1745462530
transform 1 0 2464 0 1 1770
box -7 -3 39 105
use AOI21X1  AOI21X1_10
timestamp 1745462530
transform 1 0 2392 0 -1 1970
box -7 -3 39 105
use AOI21X1  AOI21X1_11
timestamp 1745462530
transform 1 0 2360 0 1 1770
box -7 -3 39 105
use AOI21X1  AOI21X1_12
timestamp 1745462530
transform 1 0 2288 0 -1 1970
box -7 -3 39 105
use AOI21X1  AOI21X1_13
timestamp 1745462530
transform 1 0 2288 0 -1 1770
box -7 -3 39 105
use AOI21X1  AOI21X1_14
timestamp 1745462530
transform 1 0 2256 0 1 1570
box -7 -3 39 105
use AOI21X1  AOI21X1_15
timestamp 1745462530
transform 1 0 2344 0 -1 1770
box -7 -3 39 105
use AOI21X1  AOI21X1_16
timestamp 1745462530
transform 1 0 2360 0 1 1570
box -7 -3 39 105
use AOI21X1  AOI21X1_17
timestamp 1745462530
transform 1 0 920 0 1 3370
box -7 -3 39 105
use AOI21X1  AOI21X1_18
timestamp 1745462530
transform 1 0 888 0 -1 3570
box -7 -3 39 105
use AOI21X1  AOI21X1_19
timestamp 1745462530
transform 1 0 928 0 -1 3570
box -7 -3 39 105
use AOI21X1  AOI21X1_20
timestamp 1745462530
transform 1 0 880 0 1 3370
box -7 -3 39 105
use AOI21X1  AOI21X1_21
timestamp 1745462530
transform 1 0 1264 0 -1 3370
box -7 -3 39 105
use AOI21X1  AOI21X1_22
timestamp 1745462530
transform 1 0 1376 0 -1 3170
box -7 -3 39 105
use AOI21X1  AOI21X1_23
timestamp 1745462530
transform 1 0 1312 0 1 3170
box -7 -3 39 105
use AOI21X1  AOI21X1_24
timestamp 1745462530
transform 1 0 4072 0 1 2570
box -7 -3 39 105
use AOI21X1  AOI21X1_25
timestamp 1745462530
transform 1 0 3160 0 -1 2570
box -7 -3 39 105
use AOI21X1  AOI21X1_26
timestamp 1745462530
transform 1 0 4048 0 -1 2570
box -7 -3 39 105
use AOI21X1  AOI21X1_27
timestamp 1745462530
transform 1 0 3824 0 1 2570
box -7 -3 39 105
use AOI21X1  AOI21X1_28
timestamp 1745462530
transform 1 0 3328 0 1 2570
box -7 -3 39 105
use AOI21X1  AOI21X1_29
timestamp 1745462530
transform 1 0 1464 0 1 2770
box -7 -3 39 105
use AOI21X1  AOI21X1_30
timestamp 1745462530
transform 1 0 1504 0 -1 2370
box -7 -3 39 105
use AOI21X1  AOI21X1_31
timestamp 1745462530
transform 1 0 1456 0 -1 2570
box -7 -3 39 105
use AOI21X1  AOI21X1_32
timestamp 1745462530
transform 1 0 528 0 -1 2170
box -7 -3 39 105
use AOI21X1  AOI21X1_33
timestamp 1745462530
transform 1 0 632 0 1 1970
box -7 -3 39 105
use AOI21X1  AOI21X1_34
timestamp 1745462530
transform 1 0 704 0 -1 1970
box -7 -3 39 105
use AOI21X1  AOI21X1_35
timestamp 1745462530
transform 1 0 472 0 -1 1970
box -7 -3 39 105
use AOI21X1  AOI21X1_36
timestamp 1745462530
transform 1 0 920 0 1 970
box -7 -3 39 105
use AOI21X1  AOI21X1_37
timestamp 1745462530
transform 1 0 976 0 -1 1170
box -7 -3 39 105
use AOI21X1  AOI21X1_38
timestamp 1745462530
transform 1 0 1048 0 1 1170
box -7 -3 39 105
use AOI21X1  AOI21X1_39
timestamp 1745462530
transform 1 0 1096 0 1 970
box -7 -3 39 105
use AOI21X1  AOI21X1_40
timestamp 1745462530
transform 1 0 1464 0 1 970
box -7 -3 39 105
use AOI21X1  AOI21X1_41
timestamp 1745462530
transform 1 0 1448 0 -1 1170
box -7 -3 39 105
use AOI21X1  AOI21X1_42
timestamp 1745462530
transform 1 0 1528 0 -1 1370
box -7 -3 39 105
use AOI21X1  AOI21X1_43
timestamp 1745462530
transform 1 0 2296 0 1 970
box -7 -3 39 105
use AOI21X1  AOI21X1_44
timestamp 1745462530
transform 1 0 2840 0 1 970
box -7 -3 39 105
use AOI21X1  AOI21X1_45
timestamp 1745462530
transform 1 0 2792 0 1 970
box -7 -3 39 105
use AOI21X1  AOI21X1_46
timestamp 1745462530
transform 1 0 2728 0 -1 1370
box -7 -3 39 105
use AOI21X1  AOI21X1_47
timestamp 1745462530
transform 1 0 3152 0 1 970
box -7 -3 39 105
use AOI21X1  AOI21X1_48
timestamp 1745462530
transform 1 0 3240 0 1 970
box -7 -3 39 105
use AOI21X1  AOI21X1_49
timestamp 1745462530
transform 1 0 3376 0 -1 1170
box -7 -3 39 105
use AOI21X1  AOI21X1_50
timestamp 1745462530
transform 1 0 3432 0 -1 1170
box -7 -3 39 105
use AOI21X1  AOI21X1_51
timestamp 1745462530
transform 1 0 3440 0 -1 1370
box -7 -3 39 105
use AOI21X1  AOI21X1_52
timestamp 1745462530
transform 1 0 3168 0 -1 2170
box -7 -3 39 105
use AOI21X1  AOI21X1_53
timestamp 1745462530
transform 1 0 3056 0 -1 2170
box -7 -3 39 105
use AOI21X1  AOI21X1_54
timestamp 1745462530
transform 1 0 2920 0 -1 2170
box -7 -3 39 105
use AOI21X1  AOI21X1_55
timestamp 1745462530
transform 1 0 3032 0 1 2570
box -7 -3 39 105
use AOI21X1  AOI21X1_56
timestamp 1745462530
transform 1 0 3064 0 -1 2770
box -7 -3 39 105
use AOI21X1  AOI21X1_57
timestamp 1745462530
transform 1 0 3104 0 -1 2770
box -7 -3 39 105
use AOI21X1  AOI21X1_58
timestamp 1745462530
transform 1 0 2952 0 1 2770
box -7 -3 39 105
use AOI21X1  AOI21X1_59
timestamp 1745462530
transform 1 0 3016 0 -1 2770
box -7 -3 39 105
use AOI21X1  AOI21X1_60
timestamp 1745462530
transform 1 0 2992 0 1 2570
box -7 -3 39 105
use AOI21X1  AOI21X1_61
timestamp 1745462530
transform 1 0 3472 0 1 2570
box -7 -3 39 105
use AOI21X1  AOI21X1_62
timestamp 1745462530
transform 1 0 2392 0 -1 2770
box -7 -3 39 105
use AOI21X1  AOI21X1_63
timestamp 1745462530
transform 1 0 1456 0 1 3570
box -7 -3 39 105
use AOI21X1  AOI21X1_64
timestamp 1745462530
transform 1 0 1456 0 -1 3370
box -7 -3 39 105
use AOI21X1  AOI21X1_65
timestamp 1745462530
transform 1 0 1368 0 -1 3370
box -7 -3 39 105
use AOI21X1  AOI21X1_66
timestamp 1745462530
transform 1 0 656 0 1 4170
box -7 -3 39 105
use AOI21X1  AOI21X1_67
timestamp 1745462530
transform 1 0 504 0 -1 3970
box -7 -3 39 105
use AOI21X1  AOI21X1_68
timestamp 1745462530
transform 1 0 152 0 1 3770
box -7 -3 39 105
use AOI21X1  AOI21X1_69
timestamp 1745462530
transform 1 0 104 0 1 3770
box -7 -3 39 105
use AOI22X1  AOI22X1_0
timestamp 1745462530
transform 1 0 3032 0 1 3370
box -8 -3 46 105
use AOI22X1  AOI22X1_1
timestamp 1745462530
transform 1 0 3168 0 -1 3370
box -8 -3 46 105
use AOI22X1  AOI22X1_2
timestamp 1745462530
transform 1 0 3192 0 1 3370
box -8 -3 46 105
use AOI22X1  AOI22X1_3
timestamp 1745462530
transform 1 0 3216 0 -1 3370
box -8 -3 46 105
use AOI22X1  AOI22X1_4
timestamp 1745462530
transform 1 0 3112 0 1 3370
box -8 -3 46 105
use AOI22X1  AOI22X1_5
timestamp 1745462530
transform 1 0 2632 0 1 3370
box -8 -3 46 105
use AOI22X1  AOI22X1_6
timestamp 1745462530
transform 1 0 2584 0 1 3370
box -8 -3 46 105
use AOI22X1  AOI22X1_7
timestamp 1745462530
transform 1 0 2872 0 -1 3570
box -8 -3 46 105
use AOI22X1  AOI22X1_8
timestamp 1745462530
transform 1 0 3048 0 -1 3570
box -8 -3 46 105
use AOI22X1  AOI22X1_9
timestamp 1745462530
transform 1 0 3328 0 -1 3570
box -8 -3 46 105
use AOI22X1  AOI22X1_10
timestamp 1745462530
transform 1 0 3376 0 -1 3570
box -8 -3 46 105
use AOI22X1  AOI22X1_11
timestamp 1745462530
transform 1 0 3352 0 1 3370
box -8 -3 46 105
use AOI22X1  AOI22X1_12
timestamp 1745462530
transform 1 0 3096 0 -1 3570
box -8 -3 46 105
use AOI22X1  AOI22X1_13
timestamp 1745462530
transform 1 0 2488 0 -1 3570
box -8 -3 46 105
use AOI22X1  AOI22X1_14
timestamp 1745462530
transform 1 0 2432 0 -1 3570
box -8 -3 46 105
use AOI22X1  AOI22X1_15
timestamp 1745462530
transform 1 0 2784 0 -1 3570
box -8 -3 46 105
use AOI22X1  AOI22X1_16
timestamp 1745462530
transform 1 0 3000 0 -1 3570
box -8 -3 46 105
use AOI22X1  AOI22X1_17
timestamp 1745462530
transform 1 0 3256 0 -1 3570
box -8 -3 46 105
use AOI22X1  AOI22X1_18
timestamp 1745462530
transform 1 0 3248 0 1 3570
box -8 -3 46 105
use AOI22X1  AOI22X1_19
timestamp 1745462530
transform 1 0 3272 0 1 3370
box -8 -3 46 105
use AOI22X1  AOI22X1_20
timestamp 1745462530
transform 1 0 3176 0 -1 3570
box -8 -3 46 105
use AOI22X1  AOI22X1_21
timestamp 1745462530
transform 1 0 2456 0 1 3570
box -8 -3 46 105
use AOI22X1  AOI22X1_22
timestamp 1745462530
transform 1 0 2384 0 -1 3570
box -8 -3 46 105
use AOI22X1  AOI22X1_23
timestamp 1745462530
transform 1 0 2688 0 -1 3570
box -8 -3 46 105
use AOI22X1  AOI22X1_24
timestamp 1745462530
transform 1 0 2960 0 -1 3570
box -8 -3 46 105
use AOI22X1  AOI22X1_25
timestamp 1745462530
transform 1 0 3544 0 -1 3570
box -8 -3 46 105
use AOI22X1  AOI22X1_26
timestamp 1745462530
transform 1 0 3552 0 1 3570
box -8 -3 46 105
use AOI22X1  AOI22X1_27
timestamp 1745462530
transform 1 0 3496 0 -1 3570
box -8 -3 46 105
use AOI22X1  AOI22X1_28
timestamp 1745462530
transform 1 0 3456 0 -1 3570
box -8 -3 46 105
use AOI22X1  AOI22X1_29
timestamp 1745462530
transform 1 0 2600 0 -1 3570
box -8 -3 46 105
use AOI22X1  AOI22X1_30
timestamp 1745462530
transform 1 0 2544 0 -1 3570
box -8 -3 46 105
use AOI22X1  AOI22X1_31
timestamp 1745462530
transform 1 0 2720 0 1 3370
box -8 -3 46 105
use AOI22X1  AOI22X1_32
timestamp 1745462530
transform 1 0 2888 0 1 3370
box -8 -3 46 105
use AOI22X1  AOI22X1_33
timestamp 1745462530
transform 1 0 3512 0 1 3370
box -8 -3 46 105
use AOI22X1  AOI22X1_34
timestamp 1745462530
transform 1 0 3552 0 1 3370
box -8 -3 46 105
use AOI22X1  AOI22X1_35
timestamp 1745462530
transform 1 0 3472 0 1 3370
box -8 -3 46 105
use AOI22X1  AOI22X1_36
timestamp 1745462530
transform 1 0 3424 0 1 3370
box -8 -3 46 105
use AOI22X1  AOI22X1_37
timestamp 1745462530
transform 1 0 2480 0 1 3370
box -8 -3 46 105
use AOI22X1  AOI22X1_38
timestamp 1745462530
transform 1 0 2528 0 1 3370
box -8 -3 46 105
use AOI22X1  AOI22X1_39
timestamp 1745462530
transform 1 0 2752 0 -1 3370
box -8 -3 46 105
use AOI22X1  AOI22X1_40
timestamp 1745462530
transform 1 0 2928 0 -1 3370
box -8 -3 46 105
use AOI22X1  AOI22X1_41
timestamp 1745462530
transform 1 0 3440 0 -1 3370
box -8 -3 46 105
use AOI22X1  AOI22X1_42
timestamp 1745462530
transform 1 0 3488 0 -1 3370
box -8 -3 46 105
use AOI22X1  AOI22X1_43
timestamp 1745462530
transform 1 0 3392 0 -1 3370
box -8 -3 46 105
use AOI22X1  AOI22X1_44
timestamp 1745462530
transform 1 0 3344 0 -1 3370
box -8 -3 46 105
use AOI22X1  AOI22X1_45
timestamp 1745462530
transform 1 0 2496 0 -1 3370
box -8 -3 46 105
use AOI22X1  AOI22X1_46
timestamp 1745462530
transform 1 0 2560 0 -1 3370
box -8 -3 46 105
use AOI22X1  AOI22X1_47
timestamp 1745462530
transform 1 0 2760 0 1 3170
box -8 -3 46 105
use AOI22X1  AOI22X1_48
timestamp 1745462530
transform 1 0 2840 0 -1 3170
box -8 -3 46 105
use AOI22X1  AOI22X1_49
timestamp 1745462530
transform 1 0 3480 0 -1 3170
box -8 -3 46 105
use AOI22X1  AOI22X1_50
timestamp 1745462530
transform 1 0 3472 0 1 3170
box -8 -3 46 105
use AOI22X1  AOI22X1_51
timestamp 1745462530
transform 1 0 3424 0 -1 3170
box -8 -3 46 105
use AOI22X1  AOI22X1_52
timestamp 1745462530
transform 1 0 3368 0 -1 3170
box -8 -3 46 105
use AOI22X1  AOI22X1_53
timestamp 1745462530
transform 1 0 2536 0 1 3170
box -8 -3 46 105
use AOI22X1  AOI22X1_54
timestamp 1745462530
transform 1 0 2504 0 -1 3170
box -8 -3 46 105
use AOI22X1  AOI22X1_55
timestamp 1745462530
transform 1 0 2704 0 1 3170
box -8 -3 46 105
use AOI22X1  AOI22X1_56
timestamp 1745462530
transform 1 0 2872 0 1 3170
box -8 -3 46 105
use AOI22X1  AOI22X1_57
timestamp 1745462530
transform 1 0 3264 0 -1 3170
box -8 -3 46 105
use AOI22X1  AOI22X1_58
timestamp 1745462530
transform 1 0 3336 0 1 3170
box -8 -3 46 105
use AOI22X1  AOI22X1_59
timestamp 1745462530
transform 1 0 3288 0 1 3170
box -8 -3 46 105
use AOI22X1  AOI22X1_60
timestamp 1745462530
transform 1 0 3208 0 -1 3170
box -8 -3 46 105
use AOI22X1  AOI22X1_61
timestamp 1745462530
transform 1 0 2416 0 1 3170
box -8 -3 46 105
use AOI22X1  AOI22X1_62
timestamp 1745462530
transform 1 0 2864 0 -1 3370
box -8 -3 46 105
use AOI22X1  AOI22X1_63
timestamp 1745462530
transform 1 0 2424 0 -1 3170
box -8 -3 46 105
use AOI22X1  AOI22X1_64
timestamp 1745462530
transform 1 0 2048 0 -1 1770
box -8 -3 46 105
use AOI22X1  AOI22X1_65
timestamp 1745462530
transform 1 0 2000 0 1 570
box -8 -3 46 105
use AOI22X1  AOI22X1_66
timestamp 1745462530
transform 1 0 784 0 -1 2770
box -8 -3 46 105
use AOI22X1  AOI22X1_67
timestamp 1745462530
transform 1 0 3704 0 -1 1770
box -8 -3 46 105
use AOI22X1  AOI22X1_68
timestamp 1745462530
transform 1 0 3760 0 -1 2770
box -8 -3 46 105
use AOI22X1  AOI22X1_69
timestamp 1745462530
transform 1 0 3672 0 -1 770
box -8 -3 46 105
use AOI22X1  AOI22X1_70
timestamp 1745462530
transform 1 0 1888 0 1 1570
box -8 -3 46 105
use AOI22X1  AOI22X1_71
timestamp 1745462530
transform 1 0 768 0 1 570
box -8 -3 46 105
use AOI22X1  AOI22X1_72
timestamp 1745462530
transform 1 0 1816 0 -1 2770
box -8 -3 46 105
use AOI22X1  AOI22X1_73
timestamp 1745462530
transform 1 0 2488 0 1 1370
box -8 -3 46 105
use AOI22X1  AOI22X1_74
timestamp 1745462530
transform 1 0 3736 0 1 1370
box -8 -3 46 105
use AOI22X1  AOI22X1_75
timestamp 1745462530
transform 1 0 2512 0 1 570
box -8 -3 46 105
use AOI22X1  AOI22X1_76
timestamp 1745462530
transform 1 0 1040 0 1 1570
box -8 -3 46 105
use AOI22X1  AOI22X1_77
timestamp 1745462530
transform 1 0 1056 0 1 570
box -8 -3 46 105
use AOI22X1  AOI22X1_78
timestamp 1745462530
transform 1 0 744 0 -1 2770
box -8 -3 46 105
use AOI22X1  AOI22X1_79
timestamp 1745462530
transform 1 0 3496 0 -1 1770
box -8 -3 46 105
use AOI22X1  AOI22X1_80
timestamp 1745462530
transform 1 0 3576 0 -1 2770
box -8 -3 46 105
use AOI22X1  AOI22X1_81
timestamp 1745462530
transform 1 0 3616 0 1 570
box -8 -3 46 105
use AOI22X1  AOI22X1_82
timestamp 1745462530
transform 1 0 1376 0 -1 1570
box -8 -3 46 105
use AOI22X1  AOI22X1_83
timestamp 1745462530
transform 1 0 544 0 -1 970
box -8 -3 46 105
use AOI22X1  AOI22X1_84
timestamp 1745462530
transform 1 0 1512 0 1 2770
box -8 -3 46 105
use AOI22X1  AOI22X1_85
timestamp 1745462530
transform 1 0 2792 0 -1 1570
box -8 -3 46 105
use AOI22X1  AOI22X1_86
timestamp 1745462530
transform 1 0 3576 0 -1 1970
box -8 -3 46 105
use AOI22X1  AOI22X1_87
timestamp 1745462530
transform 1 0 2696 0 1 570
box -8 -3 46 105
use AOI22X1  AOI22X1_88
timestamp 1745462530
transform 1 0 1088 0 -1 1770
box -8 -3 46 105
use AOI22X1  AOI22X1_89
timestamp 1745462530
transform 1 0 1112 0 1 570
box -8 -3 46 105
use AOI22X1  AOI22X1_90
timestamp 1745462530
transform 1 0 832 0 -1 2770
box -8 -3 46 105
use AOI22X1  AOI22X1_91
timestamp 1745462530
transform 1 0 3360 0 1 1970
box -8 -3 46 105
use AOI22X1  AOI22X1_92
timestamp 1745462530
transform 1 0 3512 0 -1 2770
box -8 -3 46 105
use AOI22X1  AOI22X1_93
timestamp 1745462530
transform 1 0 3416 0 1 570
box -8 -3 46 105
use AOI22X1  AOI22X1_94
timestamp 1745462530
transform 1 0 1168 0 -1 1770
box -8 -3 46 105
use AOI22X1  AOI22X1_95
timestamp 1745462530
transform 1 0 608 0 -1 970
box -8 -3 46 105
use AOI22X1  AOI22X1_96
timestamp 1745462530
transform 1 0 1176 0 1 2770
box -8 -3 46 105
use AOI22X1  AOI22X1_97
timestamp 1745462530
transform 1 0 2488 0 -1 1970
box -8 -3 46 105
use AOI22X1  AOI22X1_98
timestamp 1745462530
transform 1 0 3568 0 1 1970
box -8 -3 46 105
use AOI22X1  AOI22X1_99
timestamp 1745462530
transform 1 0 2368 0 1 570
box -8 -3 46 105
use AOI22X1  AOI22X1_100
timestamp 1745462530
transform 1 0 1656 0 1 1770
box -8 -3 46 105
use AOI22X1  AOI22X1_101
timestamp 1745462530
transform 1 0 1616 0 1 570
box -8 -3 46 105
use AOI22X1  AOI22X1_102
timestamp 1745462530
transform 1 0 616 0 -1 2570
box -8 -3 46 105
use AOI22X1  AOI22X1_103
timestamp 1745462530
transform 1 0 4040 0 -1 1970
box -8 -3 46 105
use AOI22X1  AOI22X1_104
timestamp 1745462530
transform 1 0 4104 0 -1 2770
box -8 -3 46 105
use AOI22X1  AOI22X1_105
timestamp 1745462530
transform 1 0 3904 0 -1 570
box -8 -3 46 105
use AOI22X1  AOI22X1_106
timestamp 1745462530
transform 1 0 1984 0 -1 1970
box -8 -3 46 105
use AOI22X1  AOI22X1_107
timestamp 1745462530
transform 1 0 568 0 1 770
box -8 -3 46 105
use AOI22X1  AOI22X1_108
timestamp 1745462530
transform 1 0 1944 0 1 2570
box -8 -3 46 105
use AOI22X1  AOI22X1_109
timestamp 1745462530
transform 1 0 3128 0 -1 1970
box -8 -3 46 105
use AOI22X1  AOI22X1_110
timestamp 1745462530
transform 1 0 4040 0 -1 2170
box -8 -3 46 105
use AOI22X1  AOI22X1_111
timestamp 1745462530
transform 1 0 2952 0 1 570
box -8 -3 46 105
use AOI22X1  AOI22X1_112
timestamp 1745462530
transform 1 0 1784 0 1 1570
box -8 -3 46 105
use AOI22X1  AOI22X1_113
timestamp 1745462530
transform 1 0 1736 0 1 570
box -8 -3 46 105
use AOI22X1  AOI22X1_114
timestamp 1745462530
transform 1 0 576 0 1 2570
box -8 -3 46 105
use AOI22X1  AOI22X1_115
timestamp 1745462530
transform 1 0 4048 0 -1 1770
box -8 -3 46 105
use AOI22X1  AOI22X1_116
timestamp 1745462530
transform 1 0 4112 0 1 2570
box -8 -3 46 105
use AOI22X1  AOI22X1_117
timestamp 1745462530
transform 1 0 3840 0 -1 570
box -8 -3 46 105
use AOI22X1  AOI22X1_118
timestamp 1745462530
transform 1 0 1552 0 1 1570
box -8 -3 46 105
use AOI22X1  AOI22X1_119
timestamp 1745462530
transform 1 0 504 0 -1 770
box -8 -3 46 105
use AOI22X1  AOI22X1_120
timestamp 1745462530
transform 1 0 1656 0 1 2770
box -8 -3 46 105
use AOI22X1  AOI22X1_121
timestamp 1745462530
transform 1 0 2264 0 -1 1570
box -8 -3 46 105
use AOI22X1  AOI22X1_122
timestamp 1745462530
transform 1 0 3384 0 -1 1570
box -8 -3 46 105
use AOI22X1  AOI22X1_123
timestamp 1745462530
transform 1 0 2216 0 -1 570
box -8 -3 46 105
use AOI22X1  AOI22X1_124
timestamp 1745462530
transform 1 0 1440 0 -1 1770
box -8 -3 46 105
use AOI22X1  AOI22X1_125
timestamp 1745462530
transform 1 0 1360 0 1 570
box -8 -3 46 105
use AOI22X1  AOI22X1_126
timestamp 1745462530
transform 1 0 576 0 1 2770
box -8 -3 46 105
use AOI22X1  AOI22X1_127
timestamp 1745462530
transform 1 0 3128 0 -1 1770
box -8 -3 46 105
use AOI22X1  AOI22X1_128
timestamp 1745462530
transform 1 0 3208 0 1 2570
box -8 -3 46 105
use AOI22X1  AOI22X1_129
timestamp 1745462530
transform 1 0 3200 0 -1 570
box -8 -3 46 105
use AOI22X1  AOI22X1_130
timestamp 1745462530
transform 1 0 1144 0 1 1570
box -8 -3 46 105
use AOI22X1  AOI22X1_131
timestamp 1745462530
transform 1 0 568 0 1 570
box -8 -3 46 105
use AOI22X1  AOI22X1_132
timestamp 1745462530
transform 1 0 1336 0 1 2770
box -8 -3 46 105
use AOI22X1  AOI22X1_133
timestamp 1745462530
transform 1 0 3032 0 1 1370
box -8 -3 46 105
use AOI22X1  AOI22X1_134
timestamp 1745462530
transform 1 0 3304 0 -1 1570
box -8 -3 46 105
use AOI22X1  AOI22X1_135
timestamp 1745462530
transform 1 0 2872 0 -1 570
box -8 -3 46 105
use AOI22X1  AOI22X1_136
timestamp 1745462530
transform 1 0 3456 0 -1 3770
box -8 -3 46 105
use AOI22X1  AOI22X1_137
timestamp 1745462530
transform 1 0 3240 0 -1 3970
box -8 -3 46 105
use AOI22X1  AOI22X1_138
timestamp 1745462530
transform 1 0 3424 0 -1 4170
box -8 -3 46 105
use AOI22X1  AOI22X1_139
timestamp 1745462530
transform 1 0 3520 0 1 3770
box -8 -3 46 105
use AOI22X1  AOI22X1_140
timestamp 1745462530
transform 1 0 3544 0 -1 3970
box -8 -3 46 105
use AOI22X1  AOI22X1_141
timestamp 1745462530
transform 1 0 2048 0 -1 3770
box -8 -3 46 105
use AOI22X1  AOI22X1_142
timestamp 1745462530
transform 1 0 1696 0 -1 3770
box -8 -3 46 105
use AOI22X1  AOI22X1_143
timestamp 1745462530
transform 1 0 2320 0 -1 3970
box -8 -3 46 105
use AOI22X1  AOI22X1_144
timestamp 1745462530
transform 1 0 2336 0 -1 4170
box -8 -3 46 105
use AOI22X1  AOI22X1_145
timestamp 1745462530
transform 1 0 2016 0 1 3770
box -8 -3 46 105
use AOI22X1  AOI22X1_146
timestamp 1745462530
transform 1 0 1720 0 1 3770
box -8 -3 46 105
use AOI22X1  AOI22X1_147
timestamp 1745462530
transform 1 0 2152 0 1 3970
box -8 -3 46 105
use AOI22X1  AOI22X1_148
timestamp 1745462530
transform 1 0 2224 0 -1 4170
box -8 -3 46 105
use AOI22X1  AOI22X1_149
timestamp 1745462530
transform 1 0 3504 0 -1 3770
box -8 -3 46 105
use AOI22X1  AOI22X1_150
timestamp 1745462530
transform 1 0 3456 0 -1 3970
box -8 -3 46 105
use AOI22X1  AOI22X1_151
timestamp 1745462530
transform 1 0 3520 0 -1 4170
box -8 -3 46 105
use AOI22X1  AOI22X1_152
timestamp 1745462530
transform 1 0 3472 0 1 3770
box -8 -3 46 105
use AOI22X1  AOI22X1_153
timestamp 1745462530
transform 1 0 3544 0 1 3970
box -8 -3 46 105
use AOI22X1  AOI22X1_154
timestamp 1745462530
transform 1 0 2536 0 1 3770
box -8 -3 46 105
use AOI22X1  AOI22X1_155
timestamp 1745462530
transform 1 0 1824 0 1 3770
box -8 -3 46 105
use AOI22X1  AOI22X1_156
timestamp 1745462530
transform 1 0 2760 0 -1 3970
box -8 -3 46 105
use AOI22X1  AOI22X1_157
timestamp 1745462530
transform 1 0 2664 0 1 3970
box -8 -3 46 105
use AOI22X1  AOI22X1_158
timestamp 1745462530
transform 1 0 2616 0 1 3770
box -8 -3 46 105
use AOI22X1  AOI22X1_159
timestamp 1745462530
transform 1 0 1776 0 1 3770
box -8 -3 46 105
use AOI22X1  AOI22X1_160
timestamp 1745462530
transform 1 0 3032 0 -1 3970
box -8 -3 46 105
use AOI22X1  AOI22X1_161
timestamp 1745462530
transform 1 0 3040 0 1 3970
box -8 -3 46 105
use AOI22X1  AOI22X1_162
timestamp 1745462530
transform 1 0 968 0 -1 3370
box -8 -3 46 105
use AOI22X1  AOI22X1_163
timestamp 1745462530
transform 1 0 1120 0 -1 3570
box -8 -3 46 105
use AOI22X1  AOI22X1_164
timestamp 1745462530
transform 1 0 3912 0 1 970
box -8 -3 46 105
use AOI22X1  AOI22X1_165
timestamp 1745462530
transform 1 0 3808 0 -1 1170
box -8 -3 46 105
use AOI22X1  AOI22X1_166
timestamp 1745462530
transform 1 0 3056 0 -1 970
box -8 -3 46 105
use AOI22X1  AOI22X1_167
timestamp 1745462530
transform 1 0 2920 0 1 1170
box -8 -3 46 105
use AOI22X1  AOI22X1_168
timestamp 1745462530
transform 1 0 3928 0 -1 2770
box -8 -3 46 105
use AOI22X1  AOI22X1_169
timestamp 1745462530
transform 1 0 4040 0 -1 2770
box -8 -3 46 105
use AOI22X1  AOI22X1_170
timestamp 1745462530
transform 1 0 3816 0 -1 2170
box -8 -3 46 105
use AOI22X1  AOI22X1_171
timestamp 1745462530
transform 1 0 2984 0 -1 2170
box -8 -3 46 105
use AOI22X1  AOI22X1_172
timestamp 1745462530
transform 1 0 600 0 1 2170
box -8 -3 46 105
use AOI22X1  AOI22X1_173
timestamp 1745462530
transform 1 0 712 0 1 1970
box -8 -3 46 105
use AOI22X1  AOI22X1_174
timestamp 1745462530
transform 1 0 1976 0 -1 2970
box -8 -3 46 105
use AOI22X1  AOI22X1_175
timestamp 1745462530
transform 1 0 1960 0 1 2370
box -8 -3 46 105
use AOI22X1  AOI22X1_176
timestamp 1745462530
transform 1 0 1648 0 -1 970
box -8 -3 46 105
use AOI22X1  AOI22X1_177
timestamp 1745462530
transform 1 0 1640 0 1 1170
box -8 -3 46 105
use AOI22X1  AOI22X1_178
timestamp 1745462530
transform 1 0 672 0 -1 970
box -8 -3 46 105
use AOI22X1  AOI22X1_179
timestamp 1745462530
transform 1 0 616 0 1 1170
box -8 -3 46 105
use AOI22X1  AOI22X1_180
timestamp 1745462530
transform 1 0 3320 0 1 770
box -8 -3 46 105
use AOI22X1  AOI22X1_181
timestamp 1745462530
transform 1 0 3312 0 1 970
box -8 -3 46 105
use AOI22X1  AOI22X1_182
timestamp 1745462530
transform 1 0 3040 0 1 770
box -8 -3 46 105
use AOI22X1  AOI22X1_183
timestamp 1745462530
transform 1 0 2984 0 -1 1170
box -8 -3 46 105
use AOI22X1  AOI22X1_184
timestamp 1745462530
transform 1 0 3088 0 1 2570
box -8 -3 46 105
use AOI22X1  AOI22X1_185
timestamp 1745462530
transform 1 0 3000 0 1 2770
box -8 -3 46 105
use AOI22X1  AOI22X1_186
timestamp 1745462530
transform 1 0 3192 0 -1 1770
box -8 -3 46 105
use AOI22X1  AOI22X1_187
timestamp 1745462530
transform 1 0 2912 0 -1 1770
box -8 -3 46 105
use AOI22X1  AOI22X1_188
timestamp 1745462530
transform 1 0 632 0 -1 2170
box -8 -3 46 105
use AOI22X1  AOI22X1_189
timestamp 1745462530
transform 1 0 776 0 1 1970
box -8 -3 46 105
use AOI22X1  AOI22X1_190
timestamp 1745462530
transform 1 0 1416 0 1 2770
box -8 -3 46 105
use AOI22X1  AOI22X1_191
timestamp 1745462530
transform 1 0 1344 0 1 2370
box -8 -3 46 105
use AOI22X1  AOI22X1_192
timestamp 1745462530
transform 1 0 1464 0 1 770
box -8 -3 46 105
use AOI22X1  AOI22X1_193
timestamp 1745462530
transform 1 0 1480 0 1 1170
box -8 -3 46 105
use AOI22X1  AOI22X1_194
timestamp 1745462530
transform 1 0 672 0 -1 770
box -8 -3 46 105
use AOI22X1  AOI22X1_195
timestamp 1745462530
transform 1 0 672 0 -1 1170
box -8 -3 46 105
use AOI22X1  AOI22X1_196
timestamp 1745462530
transform 1 0 3912 0 -1 970
box -8 -3 46 105
use AOI22X1  AOI22X1_197
timestamp 1745462530
transform 1 0 3864 0 -1 1170
box -8 -3 46 105
use AOI22X1  AOI22X1_198
timestamp 1745462530
transform 1 0 2464 0 -1 970
box -8 -3 46 105
use AOI22X1  AOI22X1_199
timestamp 1745462530
transform 1 0 2432 0 1 1170
box -8 -3 46 105
use AOI22X1  AOI22X1_200
timestamp 1745462530
transform 1 0 3976 0 1 2570
box -8 -3 46 105
use AOI22X1  AOI22X1_201
timestamp 1745462530
transform 1 0 4024 0 1 2770
box -8 -3 46 105
use AOI22X1  AOI22X1_202
timestamp 1745462530
transform 1 0 3336 0 -1 1770
box -8 -3 46 105
use AOI22X1  AOI22X1_203
timestamp 1745462530
transform 1 0 2848 0 -1 1770
box -8 -3 46 105
use AOI22X1  AOI22X1_204
timestamp 1745462530
transform 1 0 576 0 -1 2170
box -8 -3 46 105
use AOI22X1  AOI22X1_205
timestamp 1745462530
transform 1 0 640 0 -1 1970
box -8 -3 46 105
use AOI22X1  AOI22X1_206
timestamp 1745462530
transform 1 0 1648 0 -1 2970
box -8 -3 46 105
use AOI22X1  AOI22X1_207
timestamp 1745462530
transform 1 0 1648 0 1 2370
box -8 -3 46 105
use AOI22X1  AOI22X1_208
timestamp 1745462530
transform 1 0 1888 0 -1 970
box -8 -3 46 105
use AOI22X1  AOI22X1_209
timestamp 1745462530
transform 1 0 1888 0 1 1170
box -8 -3 46 105
use AOI22X1  AOI22X1_210
timestamp 1745462530
transform 1 0 736 0 -1 770
box -8 -3 46 105
use AOI22X1  AOI22X1_211
timestamp 1745462530
transform 1 0 736 0 -1 1170
box -8 -3 46 105
use AOI22X1  AOI22X1_212
timestamp 1745462530
transform 1 0 3856 0 1 770
box -8 -3 46 105
use AOI22X1  AOI22X1_213
timestamp 1745462530
transform 1 0 3664 0 1 970
box -8 -3 46 105
use AOI22X1  AOI22X1_214
timestamp 1745462530
transform 1 0 2496 0 1 770
box -8 -3 46 105
use AOI22X1  AOI22X1_215
timestamp 1745462530
transform 1 0 2520 0 -1 1170
box -8 -3 46 105
use AOI22X1  AOI22X1_216
timestamp 1745462530
transform 1 0 3736 0 1 2570
box -8 -3 46 105
use AOI22X1  AOI22X1_217
timestamp 1745462530
transform 1 0 3784 0 1 2770
box -8 -3 46 105
use AOI22X1  AOI22X1_218
timestamp 1745462530
transform 1 0 3792 0 -1 1770
box -8 -3 46 105
use AOI22X1  AOI22X1_219
timestamp 1745462530
transform 1 0 2976 0 -1 1770
box -8 -3 46 105
use AOI22X1  AOI22X1_220
timestamp 1745462530
transform 1 0 776 0 -1 2170
box -8 -3 46 105
use AOI22X1  AOI22X1_221
timestamp 1745462530
transform 1 0 832 0 -1 1970
box -8 -3 46 105
use AOI22X1  AOI22X1_222
timestamp 1745462530
transform 1 0 1920 0 -1 2970
box -8 -3 46 105
use AOI22X1  AOI22X1_223
timestamp 1745462530
transform 1 0 1896 0 1 2370
box -8 -3 46 105
use AOI22X1  AOI22X1_224
timestamp 1745462530
transform 1 0 1944 0 1 770
box -8 -3 46 105
use AOI22X1  AOI22X1_225
timestamp 1745462530
transform 1 0 2056 0 -1 1170
box -8 -3 46 105
use AOI22X1  AOI22X1_226
timestamp 1745462530
transform 1 0 912 0 1 770
box -8 -3 46 105
use AOI22X1  AOI22X1_227
timestamp 1745462530
transform 1 0 808 0 -1 1170
box -8 -3 46 105
use AOI22X1  AOI22X1_228
timestamp 1745462530
transform 1 0 3480 0 1 770
box -8 -3 46 105
use AOI22X1  AOI22X1_229
timestamp 1745462530
transform 1 0 3528 0 1 970
box -8 -3 46 105
use AOI22X1  AOI22X1_230
timestamp 1745462530
transform 1 0 2624 0 1 770
box -8 -3 46 105
use AOI22X1  AOI22X1_231
timestamp 1745462530
transform 1 0 2496 0 1 1170
box -8 -3 46 105
use AOI22X1  AOI22X1_232
timestamp 1745462530
transform 1 0 3368 0 -1 2770
box -8 -3 46 105
use AOI22X1  AOI22X1_233
timestamp 1745462530
transform 1 0 3312 0 1 2770
box -8 -3 46 105
use AOI22X1  AOI22X1_234
timestamp 1745462530
transform 1 0 3432 0 -1 2170
box -8 -3 46 105
use AOI22X1  AOI22X1_235
timestamp 1745462530
transform 1 0 2928 0 1 1970
box -8 -3 46 105
use AOI22X1  AOI22X1_236
timestamp 1745462530
transform 1 0 808 0 1 2170
box -8 -3 46 105
use AOI22X1  AOI22X1_237
timestamp 1745462530
transform 1 0 904 0 -1 1970
box -8 -3 46 105
use AOI22X1  AOI22X1_238
timestamp 1745462530
transform 1 0 1432 0 -1 2970
box -8 -3 46 105
use AOI22X1  AOI22X1_239
timestamp 1745462530
transform 1 0 1176 0 1 2370
box -8 -3 46 105
use AOI22X1  AOI22X1_240
timestamp 1745462530
transform 1 0 1216 0 1 970
box -8 -3 46 105
use AOI22X1  AOI22X1_241
timestamp 1745462530
transform 1 0 1248 0 -1 1370
box -8 -3 46 105
use AOI22X1  AOI22X1_242
timestamp 1745462530
transform 1 0 880 0 -1 970
box -8 -3 46 105
use AOI22X1  AOI22X1_243
timestamp 1745462530
transform 1 0 976 0 1 1170
box -8 -3 46 105
use AOI22X1  AOI22X1_244
timestamp 1745462530
transform 1 0 3624 0 1 770
box -8 -3 46 105
use AOI22X1  AOI22X1_245
timestamp 1745462530
transform 1 0 3600 0 1 970
box -8 -3 46 105
use AOI22X1  AOI22X1_246
timestamp 1745462530
transform 1 0 2824 0 1 770
box -8 -3 46 105
use AOI22X1  AOI22X1_247
timestamp 1745462530
transform 1 0 2776 0 1 1170
box -8 -3 46 105
use AOI22X1  AOI22X1_248
timestamp 1745462530
transform 1 0 3568 0 1 2570
box -8 -3 46 105
use AOI22X1  AOI22X1_249
timestamp 1745462530
transform 1 0 3544 0 1 2770
box -8 -3 46 105
use AOI22X1  AOI22X1_250
timestamp 1745462530
transform 1 0 3536 0 -1 2170
box -8 -3 46 105
use AOI22X1  AOI22X1_251
timestamp 1745462530
transform 1 0 2992 0 1 1970
box -8 -3 46 105
use AOI22X1  AOI22X1_252
timestamp 1745462530
transform 1 0 704 0 1 2170
box -8 -3 46 105
use AOI22X1  AOI22X1_253
timestamp 1745462530
transform 1 0 768 0 -1 1970
box -8 -3 46 105
use AOI22X1  AOI22X1_254
timestamp 1745462530
transform 1 0 1488 0 -1 2970
box -8 -3 46 105
use AOI22X1  AOI22X1_255
timestamp 1745462530
transform 1 0 1528 0 1 2370
box -8 -3 46 105
use AOI22X1  AOI22X1_256
timestamp 1745462530
transform 1 0 1216 0 -1 970
box -8 -3 46 105
use AOI22X1  AOI22X1_257
timestamp 1745462530
transform 1 0 1280 0 1 1170
box -8 -3 46 105
use AOI22X1  AOI22X1_258
timestamp 1745462530
transform 1 0 784 0 1 770
box -8 -3 46 105
use AOI22X1  AOI22X1_259
timestamp 1745462530
transform 1 0 800 0 1 1170
box -8 -3 46 105
use AOI22X1  AOI22X1_260
timestamp 1745462530
transform 1 0 2160 0 -1 2970
box -8 -3 46 105
use AOI22X1  AOI22X1_261
timestamp 1745462530
transform 1 0 2160 0 1 2970
box -8 -3 46 105
use AOI22X1  AOI22X1_262
timestamp 1745462530
transform 1 0 2112 0 1 2970
box -8 -3 46 105
use AOI22X1  AOI22X1_263
timestamp 1745462530
transform 1 0 2032 0 -1 2970
box -8 -3 46 105
use AOI22X1  AOI22X1_264
timestamp 1745462530
transform 1 0 2056 0 1 2970
box -8 -3 46 105
use AOI22X1  AOI22X1_265
timestamp 1745462530
transform 1 0 2096 0 -1 2970
box -8 -3 46 105
use AOI22X1  AOI22X1_266
timestamp 1745462530
transform 1 0 232 0 1 3170
box -8 -3 46 105
use AOI22X1  AOI22X1_267
timestamp 1745462530
transform 1 0 232 0 -1 3170
box -8 -3 46 105
use AOI22X1  AOI22X1_268
timestamp 1745462530
transform 1 0 344 0 1 3170
box -8 -3 46 105
use AOI22X1  AOI22X1_269
timestamp 1745462530
transform 1 0 440 0 1 3170
box -8 -3 46 105
use AOI22X1  AOI22X1_270
timestamp 1745462530
transform 1 0 544 0 1 3170
box -8 -3 46 105
use AOI22X1  AOI22X1_271
timestamp 1745462530
transform 1 0 1544 0 1 3370
box -8 -3 46 105
use AOI22X1  AOI22X1_272
timestamp 1745462530
transform 1 0 168 0 1 3970
box -8 -3 46 105
use BUFX2  BUFX2_0
timestamp 1745462530
transform 1 0 888 0 -1 3170
box -5 -3 28 105
use BUFX2  BUFX2_1
timestamp 1745462530
transform 1 0 912 0 -1 3170
box -5 -3 28 105
use BUFX2  BUFX2_2
timestamp 1745462530
transform 1 0 1840 0 -1 3170
box -5 -3 28 105
use BUFX2  BUFX2_3
timestamp 1745462530
transform 1 0 2032 0 1 1570
box -5 -3 28 105
use BUFX2  BUFX2_4
timestamp 1745462530
transform 1 0 2008 0 -1 1770
box -5 -3 28 105
use BUFX2  BUFX2_5
timestamp 1745462530
transform 1 0 2104 0 1 1570
box -5 -3 28 105
use BUFX2  BUFX2_6
timestamp 1745462530
transform 1 0 2144 0 -1 3770
box -5 -3 28 105
use BUFX2  BUFX2_7
timestamp 1745462530
transform 1 0 2120 0 -1 3770
box -5 -3 28 105
use BUFX2  BUFX2_8
timestamp 1745462530
transform 1 0 2016 0 -1 3170
box -5 -3 28 105
use BUFX2  BUFX2_9
timestamp 1745462530
transform 1 0 2376 0 -1 3170
box -5 -3 28 105
use BUFX2  BUFX2_10
timestamp 1745462530
transform 1 0 1616 0 -1 3970
box -5 -3 28 105
use BUFX2  BUFX2_11
timestamp 1745462530
transform 1 0 3928 0 -1 3970
box -5 -3 28 105
use BUFX2  BUFX2_12
timestamp 1745462530
transform 1 0 3928 0 -1 3170
box -5 -3 28 105
use BUFX2  BUFX2_13
timestamp 1745462530
transform 1 0 2136 0 1 1370
box -5 -3 28 105
use BUFX2  BUFX2_14
timestamp 1745462530
transform 1 0 2128 0 1 1570
box -5 -3 28 105
use BUFX2  BUFX2_15
timestamp 1745462530
transform 1 0 1960 0 1 1570
box -5 -3 28 105
use BUFX2  BUFX2_16
timestamp 1745462530
transform 1 0 2056 0 1 1570
box -5 -3 28 105
use BUFX2  BUFX2_17
timestamp 1745462530
transform 1 0 1984 0 -1 1770
box -5 -3 28 105
use BUFX2  BUFX2_18
timestamp 1745462530
transform 1 0 1984 0 1 1570
box -5 -3 28 105
use BUFX2  BUFX2_19
timestamp 1745462530
transform 1 0 2208 0 -1 1570
box -5 -3 28 105
use BUFX2  BUFX2_20
timestamp 1745462530
transform 1 0 2112 0 -1 1770
box -5 -3 28 105
use BUFX2  BUFX2_21
timestamp 1745462530
transform 1 0 2144 0 -1 1570
box -5 -3 28 105
use BUFX2  BUFX2_22
timestamp 1745462530
transform 1 0 1360 0 1 2170
box -5 -3 28 105
use BUFX2  BUFX2_23
timestamp 1745462530
transform 1 0 2616 0 -1 1570
box -5 -3 28 105
use BUFX2  BUFX2_24
timestamp 1745462530
transform 1 0 1304 0 -1 1570
box -5 -3 28 105
use BUFX2  BUFX2_25
timestamp 1745462530
transform 1 0 1376 0 -1 2170
box -5 -3 28 105
use BUFX2  BUFX2_26
timestamp 1745462530
transform 1 0 2576 0 -1 2170
box -5 -3 28 105
use BUFX2  BUFX2_27
timestamp 1745462530
transform 1 0 2064 0 1 1770
box -5 -3 28 105
use BUFX2  BUFX2_28
timestamp 1745462530
transform 1 0 2216 0 -1 1770
box -5 -3 28 105
use BUFX2  BUFX2_29
timestamp 1745462530
transform 1 0 2088 0 1 1770
box -5 -3 28 105
use BUFX2  BUFX2_30
timestamp 1745462530
transform 1 0 1744 0 -1 2170
box -5 -3 28 105
use BUFX2  BUFX2_31
timestamp 1745462530
transform 1 0 2264 0 1 3170
box -5 -3 28 105
use BUFX2  BUFX2_32
timestamp 1745462530
transform 1 0 2040 0 -1 3170
box -5 -3 28 105
use BUFX2  BUFX2_33
timestamp 1745462530
transform 1 0 2480 0 -1 2770
box -5 -3 28 105
use BUFX2  BUFX2_34
timestamp 1745462530
transform 1 0 2568 0 1 2570
box -5 -3 28 105
use BUFX2  BUFX2_35
timestamp 1745462530
transform 1 0 2544 0 1 2570
box -5 -3 28 105
use BUFX2  BUFX2_36
timestamp 1745462530
transform 1 0 2632 0 1 2570
box -5 -3 28 105
use BUFX2  BUFX2_37
timestamp 1745462530
transform 1 0 2608 0 1 2570
box -5 -3 28 105
use BUFX2  BUFX2_38
timestamp 1745462530
transform 1 0 2440 0 1 2370
box -5 -3 28 105
use BUFX2  BUFX2_39
timestamp 1745462530
transform 1 0 2504 0 1 2370
box -5 -3 28 105
use BUFX2  BUFX2_40
timestamp 1745462530
transform 1 0 2408 0 1 2370
box -5 -3 28 105
use BUFX2  BUFX2_41
timestamp 1745462530
transform 1 0 2472 0 1 2370
box -5 -3 28 105
use BUFX2  BUFX2_42
timestamp 1745462530
transform 1 0 2464 0 -1 2370
box -5 -3 28 105
use BUFX2  BUFX2_43
timestamp 1745462530
transform 1 0 2488 0 -1 2370
box -5 -3 28 105
use BUFX2  BUFX2_44
timestamp 1745462530
transform 1 0 2520 0 -1 2370
box -5 -3 28 105
use BUFX2  BUFX2_45
timestamp 1745462530
transform 1 0 2544 0 -1 2370
box -5 -3 28 105
use BUFX2  BUFX2_46
timestamp 1745462530
transform 1 0 2456 0 -1 2770
box -5 -3 28 105
use BUFX2  BUFX2_47
timestamp 1745462530
transform 1 0 2512 0 1 2570
box -5 -3 28 105
use BUFX2  BUFX2_48
timestamp 1745462530
transform 1 0 2432 0 -1 2770
box -5 -3 28 105
use BUFX2  BUFX2_49
timestamp 1745462530
transform 1 0 976 0 -1 3170
box -5 -3 28 105
use BUFX2  BUFX2_50
timestamp 1745462530
transform 1 0 1000 0 -1 3170
box -5 -3 28 105
use BUFX2  BUFX2_51
timestamp 1745462530
transform 1 0 944 0 -1 3170
box -5 -3 28 105
use BUFX2  BUFX2_52
timestamp 1745462530
transform 1 0 2136 0 1 3770
box -5 -3 28 105
use BUFX2  BUFX2_53
timestamp 1745462530
transform 1 0 2224 0 -1 1970
box -5 -3 28 105
use BUFX2  BUFX2_54
timestamp 1745462530
transform 1 0 1608 0 1 3970
box -5 -3 28 105
use BUFX2  BUFX2_55
timestamp 1745462530
transform 1 0 2240 0 1 3770
box -5 -3 28 105
use BUFX2  BUFX2_56
timestamp 1745462530
transform 1 0 2184 0 -1 3970
box -5 -3 28 105
use BUFX2  BUFX2_57
timestamp 1745462530
transform 1 0 2272 0 -1 3970
box -5 -3 28 105
use BUFX2  BUFX2_58
timestamp 1745462530
transform 1 0 2128 0 -1 3970
box -5 -3 28 105
use BUFX2  BUFX2_59
timestamp 1745462530
transform 1 0 2152 0 -1 3970
box -5 -3 28 105
use BUFX2  BUFX2_60
timestamp 1745462530
transform 1 0 2568 0 -1 2570
box -5 -3 28 105
use BUFX2  BUFX2_61
timestamp 1745462530
transform 1 0 2352 0 -1 2170
box -5 -3 28 105
use BUFX2  BUFX2_62
timestamp 1745462530
transform 1 0 2536 0 -1 2570
box -5 -3 28 105
use BUFX2  BUFX2_63
timestamp 1745462530
transform 1 0 2328 0 1 1970
box -5 -3 28 105
use BUFX2  BUFX2_64
timestamp 1745462530
transform 1 0 2592 0 1 2370
box -5 -3 28 105
use BUFX2  BUFX2_65
timestamp 1745462530
transform 1 0 2320 0 -1 2170
box -5 -3 28 105
use BUFX2  BUFX2_66
timestamp 1745462530
transform 1 0 2608 0 -1 2570
box -5 -3 28 105
use BUFX2  BUFX2_67
timestamp 1745462530
transform 1 0 2304 0 1 1970
box -5 -3 28 105
use BUFX2  BUFX2_68
timestamp 1745462530
transform 1 0 2456 0 1 1970
box -5 -3 28 105
use BUFX2  BUFX2_69
timestamp 1745462530
transform 1 0 2488 0 -1 2170
box -5 -3 28 105
use BUFX2  BUFX2_70
timestamp 1745462530
transform 1 0 2464 0 -1 2170
box -5 -3 28 105
use BUFX2  BUFX2_71
timestamp 1745462530
transform 1 0 2480 0 1 1970
box -5 -3 28 105
use BUFX2  BUFX2_72
timestamp 1745462530
transform 1 0 2392 0 1 1970
box -5 -3 28 105
use BUFX2  BUFX2_73
timestamp 1745462530
transform 1 0 2408 0 -1 2170
box -5 -3 28 105
use BUFX2  BUFX2_74
timestamp 1745462530
transform 1 0 2376 0 -1 2170
box -5 -3 28 105
use BUFX2  BUFX2_75
timestamp 1745462530
transform 1 0 2416 0 1 1970
box -5 -3 28 105
use BUFX2  BUFX2_76
timestamp 1745462530
transform 1 0 1344 0 -1 3970
box -5 -3 28 105
use BUFX2  BUFX2_77
timestamp 1745462530
transform 1 0 1320 0 -1 3970
box -5 -3 28 105
use BUFX2  BUFX2_78
timestamp 1745462530
transform 1 0 3864 0 -1 3970
box -5 -3 28 105
use BUFX2  BUFX2_79
timestamp 1745462530
transform 1 0 3888 0 -1 3970
box -5 -3 28 105
use BUFX2  BUFX2_80
timestamp 1745462530
transform 1 0 3952 0 -1 3970
box -5 -3 28 105
use BUFX2  BUFX2_81
timestamp 1745462530
transform 1 0 4000 0 -1 3170
box -5 -3 28 105
use BUFX2  BUFX2_82
timestamp 1745462530
transform 1 0 4024 0 -1 3170
box -5 -3 28 105
use BUFX2  BUFX2_83
timestamp 1745462530
transform 1 0 3952 0 -1 3170
box -5 -3 28 105
use BUFX2  BUFX2_84
timestamp 1745462530
transform 1 0 2136 0 -1 1370
box -5 -3 28 105
use BUFX2  BUFX2_85
timestamp 1745462530
transform 1 0 1816 0 -1 1370
box -5 -3 28 105
use BUFX2  BUFX2_86
timestamp 1745462530
transform 1 0 1792 0 -1 1570
box -5 -3 28 105
use BUFX2  BUFX2_87
timestamp 1745462530
transform 1 0 2184 0 1 1970
box -5 -3 28 105
use BUFX2  BUFX2_88
timestamp 1745462530
transform 1 0 2264 0 1 1970
box -5 -3 28 105
use BUFX2  BUFX2_89
timestamp 1745462530
transform 1 0 2176 0 1 1570
box -5 -3 28 105
use BUFX2  BUFX2_90
timestamp 1745462530
transform 1 0 1328 0 1 1370
box -5 -3 28 105
use BUFX2  BUFX2_91
timestamp 1745462530
transform 1 0 1328 0 -1 1570
box -5 -3 28 105
use BUFX2  BUFX2_92
timestamp 1745462530
transform 1 0 1440 0 1 1570
box -5 -3 28 105
use BUFX2  BUFX2_93
timestamp 1745462530
transform 1 0 2200 0 1 1570
box -5 -3 28 105
use BUFX2  BUFX2_94
timestamp 1745462530
transform 1 0 2120 0 -1 1570
box -5 -3 28 105
use BUFX2  BUFX2_95
timestamp 1745462530
transform 1 0 1576 0 1 1370
box -5 -3 28 105
use BUFX2  BUFX2_96
timestamp 1745462530
transform 1 0 1960 0 1 1770
box -5 -3 28 105
use BUFX2  BUFX2_97
timestamp 1745462530
transform 1 0 2288 0 1 1770
box -5 -3 28 105
use BUFX2  BUFX2_98
timestamp 1745462530
transform 1 0 2248 0 1 1770
box -5 -3 28 105
use BUFX2  BUFX2_99
timestamp 1745462530
transform 1 0 1968 0 -1 1570
box -5 -3 28 105
use BUFX2  BUFX2_100
timestamp 1745462530
transform 1 0 1944 0 -1 1570
box -5 -3 28 105
use BUFX2  BUFX2_101
timestamp 1745462530
transform 1 0 1952 0 -1 1770
box -5 -3 28 105
use BUFX2  BUFX2_102
timestamp 1745462530
transform 1 0 2552 0 -1 1570
box -5 -3 28 105
use BUFX2  BUFX2_103
timestamp 1745462530
transform 1 0 2584 0 -1 1570
box -5 -3 28 105
use BUFX2  BUFX2_104
timestamp 1745462530
transform 1 0 2216 0 1 1370
box -5 -3 28 105
use BUFX2  BUFX2_105
timestamp 1745462530
transform 1 0 1616 0 -1 1770
box -5 -3 28 105
use BUFX2  BUFX2_106
timestamp 1745462530
transform 1 0 2088 0 -1 1970
box -5 -3 28 105
use BUFX2  BUFX2_107
timestamp 1745462530
transform 1 0 2248 0 -1 1970
box -5 -3 28 105
use BUFX2  BUFX2_108
timestamp 1745462530
transform 1 0 2184 0 -1 1570
box -5 -3 28 105
use BUFX2  BUFX2_109
timestamp 1745462530
transform 1 0 2176 0 1 1370
box -5 -3 28 105
use BUFX2  BUFX2_110
timestamp 1745462530
transform 1 0 904 0 -1 1570
box -5 -3 28 105
use BUFX2  BUFX2_111
timestamp 1745462530
transform 1 0 2664 0 1 2570
box -5 -3 28 105
use BUFX2  BUFX2_112
timestamp 1745462530
transform 1 0 2448 0 1 2170
box -5 -3 28 105
use BUFX2  BUFX2_113
timestamp 1745462530
transform 1 0 1840 0 -1 2170
box -5 -3 28 105
use BUFX2  BUFX2_114
timestamp 1745462530
transform 1 0 2160 0 -1 1770
box -5 -3 28 105
use BUFX2  BUFX2_115
timestamp 1745462530
transform 1 0 1648 0 -1 1770
box -5 -3 28 105
use BUFX2  BUFX2_116
timestamp 1745462530
transform 1 0 2208 0 1 1970
box -5 -3 28 105
use BUFX2  BUFX2_117
timestamp 1745462530
transform 1 0 1504 0 1 1970
box -5 -3 28 105
use BUFX2  BUFX2_118
timestamp 1745462530
transform 1 0 2568 0 1 1570
box -5 -3 28 105
use BUFX2  BUFX2_119
timestamp 1745462530
transform 1 0 1624 0 1 1570
box -5 -3 28 105
use BUFX2  BUFX2_120
timestamp 1745462530
transform 1 0 2136 0 -1 1770
box -5 -3 28 105
use BUFX2  BUFX2_121
timestamp 1745462530
transform 1 0 1840 0 1 1570
box -5 -3 28 105
use BUFX2  BUFX2_122
timestamp 1745462530
transform 1 0 2360 0 1 1970
box -5 -3 28 105
use BUFX2  BUFX2_123
timestamp 1745462530
transform 1 0 1144 0 -1 2170
box -5 -3 28 105
use BUFX2  BUFX2_124
timestamp 1745462530
transform 1 0 2320 0 1 2170
box -5 -3 28 105
use BUFX2  BUFX2_125
timestamp 1745462530
transform 1 0 1592 0 -1 1370
box -5 -3 28 105
use BUFX2  BUFX2_126
timestamp 1745462530
transform 1 0 1496 0 -1 1970
box -5 -3 28 105
use BUFX2  BUFX2_127
timestamp 1745462530
transform 1 0 2984 0 -1 2770
box -5 -3 28 105
use BUFX2  BUFX2_128
timestamp 1745462530
transform 1 0 2688 0 1 2570
box -5 -3 28 105
use BUFX2  BUFX2_129
timestamp 1745462530
transform 1 0 2944 0 1 2570
box -5 -3 28 105
use BUFX2  BUFX2_130
timestamp 1745462530
transform 1 0 2160 0 -1 1370
box -5 -3 28 105
use BUFX2  BUFX2_131
timestamp 1745462530
transform 1 0 2200 0 -1 3170
box -5 -3 28 105
use BUFX2  BUFX2_132
timestamp 1745462530
transform 1 0 2104 0 -1 3170
box -5 -3 28 105
use BUFX2  BUFX2_133
timestamp 1745462530
transform 1 0 1848 0 1 2170
box -5 -3 28 105
use BUFX2  BUFX2_134
timestamp 1745462530
transform 1 0 1528 0 1 1970
box -5 -3 28 105
use BUFX2  BUFX2_135
timestamp 1745462530
transform 1 0 1288 0 1 1570
box -5 -3 28 105
use BUFX2  BUFX2_136
timestamp 1745462530
transform 1 0 1680 0 -1 1770
box -5 -3 28 105
use BUFX2  BUFX2_137
timestamp 1745462530
transform 1 0 1856 0 -1 1770
box -5 -3 28 105
use BUFX2  BUFX2_138
timestamp 1745462530
transform 1 0 1160 0 1 2170
box -5 -3 28 105
use BUFX2  BUFX2_139
timestamp 1745462530
transform 1 0 3800 0 1 2170
box -5 -3 28 105
use BUFX2  BUFX2_140
timestamp 1745462530
transform 1 0 3800 0 -1 1970
box -5 -3 28 105
use BUFX2  BUFX2_141
timestamp 1745462530
transform 1 0 2552 0 1 1370
box -5 -3 28 105
use BUFX2  BUFX2_142
timestamp 1745462530
transform 1 0 1760 0 -1 1570
box -5 -3 28 105
use BUFX2  BUFX2_143
timestamp 1745462530
transform 1 0 1768 0 1 1970
box -5 -3 28 105
use BUFX2  BUFX2_144
timestamp 1745462530
transform 1 0 2552 0 1 1970
box -5 -3 28 105
use BUFX2  BUFX2_145
timestamp 1745462530
transform 1 0 2576 0 1 1970
box -5 -3 28 105
use BUFX2  BUFX2_146
timestamp 1745462530
transform 1 0 2208 0 1 1770
box -5 -3 28 105
use BUFX2  BUFX2_147
timestamp 1745462530
transform 1 0 1304 0 1 1370
box -5 -3 28 105
use BUFX2  BUFX2_148
timestamp 1745462530
transform 1 0 1296 0 -1 1770
box -5 -3 28 105
use BUFX2  BUFX2_149
timestamp 1745462530
transform 1 0 2864 0 -1 1570
box -5 -3 28 105
use BUFX2  BUFX2_150
timestamp 1745462530
transform 1 0 2888 0 -1 1570
box -5 -3 28 105
use BUFX2  BUFX2_151
timestamp 1745462530
transform 1 0 2576 0 1 1370
box -5 -3 28 105
use BUFX2  BUFX2_152
timestamp 1745462530
transform 1 0 1272 0 -1 1570
box -5 -3 28 105
use BUFX2  BUFX2_153
timestamp 1745462530
transform 1 0 1216 0 1 1570
box -5 -3 28 105
use BUFX2  BUFX2_154
timestamp 1745462530
transform 1 0 2720 0 -1 1770
box -5 -3 28 105
use BUFX2  BUFX2_155
timestamp 1745462530
transform 1 0 2704 0 1 1570
box -5 -3 28 105
use BUFX2  BUFX2_156
timestamp 1745462530
transform 1 0 2312 0 1 1570
box -5 -3 28 105
use BUFX2  BUFX2_157
timestamp 1745462530
transform 1 0 1672 0 -1 1570
box -5 -3 28 105
use BUFX2  BUFX2_158
timestamp 1745462530
transform 1 0 1704 0 -1 1770
box -5 -3 28 105
use BUFX2  BUFX2_159
timestamp 1745462530
transform 1 0 2696 0 -1 1770
box -5 -3 28 105
use BUFX2  BUFX2_160
timestamp 1745462530
transform 1 0 2728 0 1 1570
box -5 -3 28 105
use BUFX2  BUFX2_161
timestamp 1745462530
transform 1 0 2184 0 -1 1370
box -5 -3 28 105
use BUFX2  BUFX2_162
timestamp 1745462530
transform 1 0 1784 0 1 1370
box -5 -3 28 105
use BUFX2  BUFX2_163
timestamp 1745462530
transform 1 0 1784 0 -1 1770
box -5 -3 28 105
use BUFX2  BUFX2_164
timestamp 1745462530
transform 1 0 2840 0 1 2170
box -5 -3 28 105
use BUFX2  BUFX2_165
timestamp 1745462530
transform 1 0 3264 0 1 1970
box -5 -3 28 105
use BUFX2  BUFX2_166
timestamp 1745462530
transform 1 0 2416 0 1 1770
box -5 -3 28 105
use BUFX2  BUFX2_167
timestamp 1745462530
transform 1 0 1112 0 -1 1370
box -5 -3 28 105
use BUFX2  BUFX2_168
timestamp 1745462530
transform 1 0 1104 0 1 1570
box -5 -3 28 105
use BUFX2  BUFX2_169
timestamp 1745462530
transform 1 0 2128 0 -1 3170
box -5 -3 28 105
use BUFX2  BUFX2_170
timestamp 1745462530
transform 1 0 2184 0 1 3570
box -5 -3 28 105
use BUFX2  BUFX2_171
timestamp 1745462530
transform 1 0 2208 0 1 3570
box -5 -3 28 105
use BUFX2  BUFX2_172
timestamp 1745462530
transform 1 0 2192 0 -1 3570
box -5 -3 28 105
use BUFX2  BUFX2_173
timestamp 1745462530
transform 1 0 2048 0 1 3170
box -5 -3 28 105
use BUFX2  BUFX2_174
timestamp 1745462530
transform 1 0 2064 0 -1 3170
box -5 -3 28 105
use DFFNEGX1  DFFNEGX1_0
timestamp 1745462530
transform 1 0 416 0 -1 3770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_1
timestamp 1745462530
transform 1 0 368 0 1 3370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_2
timestamp 1745462530
transform 1 0 136 0 -1 3370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_3
timestamp 1745462530
transform 1 0 392 0 1 3570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_4
timestamp 1745462530
transform 1 0 280 0 -1 3770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_5
timestamp 1745462530
transform 1 0 144 0 -1 3770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_6
timestamp 1745462530
transform 1 0 80 0 1 3370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_7
timestamp 1745462530
transform 1 0 80 0 1 3570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_8
timestamp 1745462530
transform 1 0 504 0 1 3570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_9
timestamp 1745462530
transform 1 0 728 0 -1 3770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_10
timestamp 1745462530
transform 1 0 840 0 -1 3770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_11
timestamp 1745462530
transform 1 0 448 0 -1 3570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_12
timestamp 1745462530
transform 1 0 624 0 1 3570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_13
timestamp 1745462530
transform 1 0 568 0 -1 3570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_14
timestamp 1745462530
transform 1 0 488 0 1 3370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_15
timestamp 1745462530
transform 1 0 592 0 1 3370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_16
timestamp 1745462530
transform 1 0 488 0 -1 3370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_17
timestamp 1745462530
transform 1 0 1168 0 -1 3170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_18
timestamp 1745462530
transform 1 0 1160 0 -1 3370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_19
timestamp 1745462530
transform 1 0 1160 0 1 3570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_20
timestamp 1745462530
transform 1 0 80 0 1 3170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_21
timestamp 1745462530
transform 1 0 680 0 -1 3170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_22
timestamp 1745462530
transform 1 0 600 0 -1 3370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_23
timestamp 1745462530
transform 1 0 368 0 -1 3370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_24
timestamp 1745462530
transform 1 0 256 0 -1 3370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_25
timestamp 1745462530
transform 1 0 88 0 -1 3170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_26
timestamp 1745462530
transform 1 0 2088 0 -1 2770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_27
timestamp 1745462530
transform 1 0 2256 0 1 2970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_28
timestamp 1745462530
transform 1 0 2352 0 1 2770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_29
timestamp 1745462530
transform 1 0 2272 0 -1 2970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_30
timestamp 1745462530
transform 1 0 2184 0 1 2770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_31
timestamp 1745462530
transform 1 0 1984 0 -1 2770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_32
timestamp 1745462530
transform 1 0 720 0 -1 3370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_33
timestamp 1745462530
transform 1 0 1032 0 -1 3170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_34
timestamp 1745462530
transform 1 0 704 0 1 3370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_35
timestamp 1745462530
transform 1 0 1024 0 -1 3770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_36
timestamp 1745462530
transform 1 0 888 0 1 3570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_37
timestamp 1745462530
transform 1 0 752 0 1 3570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_38
timestamp 1745462530
transform 1 0 680 0 -1 3570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_39
timestamp 1745462530
transform 1 0 840 0 -1 3370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_40
timestamp 1745462530
transform 1 0 1392 0 1 3170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_41
timestamp 1745462530
transform 1 0 1280 0 1 3370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_42
timestamp 1745462530
transform 1 0 1168 0 1 3370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_43
timestamp 1745462530
transform 1 0 1456 0 -1 3170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_44
timestamp 1745462530
transform 1 0 1400 0 1 2970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_45
timestamp 1745462530
transform 1 0 1264 0 -1 3570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_46
timestamp 1745462530
transform 1 0 1136 0 1 3170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_47
timestamp 1745462530
transform 1 0 1152 0 -1 3770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_48
timestamp 1745462530
transform 1 0 968 0 1 2970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_49
timestamp 1745462530
transform 1 0 1040 0 1 2770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_50
timestamp 1745462530
transform 1 0 1008 0 -1 2370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_51
timestamp 1745462530
transform 1 0 1072 0 -1 2770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_52
timestamp 1745462530
transform 1 0 968 0 -1 2170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_53
timestamp 1745462530
transform 1 0 1040 0 -1 2570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_54
timestamp 1745462530
transform 1 0 1096 0 1 1970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_55
timestamp 1745462530
transform 1 0 856 0 1 2970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_56
timestamp 1745462530
transform 1 0 800 0 -1 2570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_57
timestamp 1745462530
transform 1 0 80 0 1 2570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_58
timestamp 1745462530
transform 1 0 80 0 1 2170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_59
timestamp 1745462530
transform 1 0 80 0 -1 2170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_60
timestamp 1745462530
transform 1 0 80 0 -1 1770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_61
timestamp 1745462530
transform 1 0 784 0 1 1570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_62
timestamp 1745462530
transform 1 0 80 0 1 1370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_63
timestamp 1745462530
transform 1 0 80 0 1 970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_64
timestamp 1745462530
transform 1 0 88 0 -1 570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_65
timestamp 1745462530
transform 1 0 80 0 1 570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_66
timestamp 1745462530
transform 1 0 640 0 1 570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_67
timestamp 1745462530
transform 1 0 848 0 1 570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_68
timestamp 1745462530
transform 1 0 80 0 -1 1370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_69
timestamp 1745462530
transform 1 0 1008 0 -1 1370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_70
timestamp 1745462530
transform 1 0 968 0 -1 370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_71
timestamp 1745462530
transform 1 0 1000 0 1 370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_72
timestamp 1745462530
transform 1 0 1184 0 -1 370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_73
timestamp 1745462530
transform 1 0 1176 0 1 770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_74
timestamp 1745462530
transform 1 0 1232 0 1 370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_75
timestamp 1745462530
transform 1 0 1272 0 1 970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_76
timestamp 1745462530
transform 1 0 1304 0 -1 1370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_77
timestamp 1745462530
transform 1 0 1368 0 1 1370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_78
timestamp 1745462530
transform 1 0 2088 0 -1 370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_79
timestamp 1745462530
transform 1 0 2072 0 -1 770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_80
timestamp 1745462530
transform 1 0 2080 0 1 170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_81
timestamp 1745462530
transform 1 0 2096 0 -1 570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_82
timestamp 1745462530
transform 1 0 2584 0 1 370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_83
timestamp 1745462530
transform 1 0 2600 0 -1 970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_84
timestamp 1745462530
transform 1 0 2320 0 1 1170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_85
timestamp 1745462530
transform 1 0 2328 0 -1 1570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_86
timestamp 1745462530
transform 1 0 3216 0 1 370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_87
timestamp 1745462530
transform 1 0 3400 0 1 370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_88
timestamp 1745462530
transform 1 0 3984 0 -1 570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_89
timestamp 1745462530
transform 1 0 3456 0 -1 770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_90
timestamp 1745462530
transform 1 0 3944 0 1 570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_91
timestamp 1745462530
transform 1 0 3848 0 -1 770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_92
timestamp 1745462530
transform 1 0 3424 0 -1 970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_93
timestamp 1745462530
transform 1 0 3472 0 -1 1170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_94
timestamp 1745462530
transform 1 0 3936 0 1 1370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_95
timestamp 1745462530
transform 1 0 3352 0 1 1770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_96
timestamp 1745462530
transform 1 0 4064 0 1 1770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_97
timestamp 1745462530
transform 1 0 3600 0 -1 2170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_98
timestamp 1745462530
transform 1 0 4088 0 -1 2170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_99
timestamp 1745462530
transform 1 0 3424 0 1 2170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_100
timestamp 1745462530
transform 1 0 2664 0 1 2170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_101
timestamp 1745462530
transform 1 0 2480 0 1 2170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_102
timestamp 1745462530
transform 1 0 3440 0 1 2770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_103
timestamp 1745462530
transform 1 0 3240 0 1 2970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_104
timestamp 1745462530
transform 1 0 3360 0 -1 2970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_105
timestamp 1745462530
transform 1 0 3352 0 1 2970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_106
timestamp 1745462530
transform 1 0 3376 0 -1 2570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_107
timestamp 1745462530
transform 1 0 3408 0 -1 2370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_108
timestamp 1745462530
transform 1 0 2832 0 1 2770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_109
timestamp 1745462530
transform 1 0 2728 0 1 2570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_110
timestamp 1745462530
transform 1 0 2648 0 -1 2970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_111
timestamp 1745462530
transform 1 0 1000 0 -1 2970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_112
timestamp 1745462530
transform 1 0 1808 0 -1 2970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_113
timestamp 1745462530
transform 1 0 1904 0 -1 2170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_114
timestamp 1745462530
transform 1 0 1864 0 -1 2770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_115
timestamp 1745462530
transform 1 0 1968 0 1 1970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_116
timestamp 1745462530
transform 1 0 1704 0 1 2570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_117
timestamp 1745462530
transform 1 0 1872 0 -1 1970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_118
timestamp 1745462530
transform 1 0 744 0 1 2970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_119
timestamp 1745462530
transform 1 0 640 0 1 2970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_120
timestamp 1745462530
transform 1 0 432 0 -1 2970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_121
timestamp 1745462530
transform 1 0 344 0 -1 2170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_122
timestamp 1745462530
transform 1 0 240 0 1 1970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_123
timestamp 1745462530
transform 1 0 296 0 -1 1770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_124
timestamp 1745462530
transform 1 0 752 0 -1 1770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_125
timestamp 1745462530
transform 1 0 200 0 1 1370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_126
timestamp 1745462530
transform 1 0 80 0 1 770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_127
timestamp 1745462530
transform 1 0 88 0 1 170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_128
timestamp 1745462530
transform 1 0 88 0 1 370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_129
timestamp 1745462530
transform 1 0 760 0 1 370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_130
timestamp 1745462530
transform 1 0 880 0 1 370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_131
timestamp 1745462530
transform 1 0 104 0 1 1170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_132
timestamp 1745462530
transform 1 0 792 0 -1 1570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_133
timestamp 1745462530
transform 1 0 1560 0 1 170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_134
timestamp 1745462530
transform 1 0 1976 0 1 370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_135
timestamp 1745462530
transform 1 0 1968 0 1 170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_136
timestamp 1745462530
transform 1 0 1960 0 -1 770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_137
timestamp 1745462530
transform 1 0 1976 0 -1 370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_138
timestamp 1745462530
transform 1 0 2048 0 -1 970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_139
timestamp 1745462530
transform 1 0 2144 0 -1 1170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_140
timestamp 1745462530
transform 1 0 2064 0 1 1170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_141
timestamp 1745462530
transform 1 0 2344 0 1 170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_142
timestamp 1745462530
transform 1 0 2328 0 -1 770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_143
timestamp 1745462530
transform 1 0 2456 0 1 170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_144
timestamp 1745462530
transform 1 0 2344 0 1 370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_145
timestamp 1745462530
transform 1 0 2448 0 1 370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_146
timestamp 1745462530
transform 1 0 2144 0 1 770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_147
timestamp 1745462530
transform 1 0 2560 0 1 970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_148
timestamp 1745462530
transform 1 0 2552 0 1 1170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_149
timestamp 1745462530
transform 1 0 3424 0 -1 370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_150
timestamp 1745462530
transform 1 0 3680 0 -1 570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_151
timestamp 1745462530
transform 1 0 4272 0 1 370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_152
timestamp 1745462530
transform 1 0 3832 0 1 570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_153
timestamp 1745462530
transform 1 0 4280 0 -1 570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_154
timestamp 1745462530
transform 1 0 4120 0 -1 770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_155
timestamp 1745462530
transform 1 0 3744 0 -1 970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_156
timestamp 1745462530
transform 1 0 3696 0 -1 1170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_157
timestamp 1745462530
transform 1 0 4176 0 1 1170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_158
timestamp 1745462530
transform 1 0 3744 0 -1 1370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_159
timestamp 1745462530
transform 1 0 4272 0 1 1370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_160
timestamp 1745462530
transform 1 0 3864 0 1 1570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_161
timestamp 1745462530
transform 1 0 3976 0 1 1570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_162
timestamp 1745462530
transform 1 0 3936 0 -1 1770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_163
timestamp 1745462530
transform 1 0 3048 0 1 1770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_164
timestamp 1745462530
transform 1 0 2528 0 1 1770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_165
timestamp 1745462530
transform 1 0 3864 0 1 2570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_166
timestamp 1745462530
transform 1 0 3640 0 -1 3170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_167
timestamp 1745462530
transform 1 0 3896 0 1 2770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_168
timestamp 1745462530
transform 1 0 3784 0 -1 2970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_169
timestamp 1745462530
transform 1 0 3880 0 -1 2570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_170
timestamp 1745462530
transform 1 0 3968 0 -1 2370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_171
timestamp 1745462530
transform 1 0 3808 0 -1 3170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_172
timestamp 1745462530
transform 1 0 3048 0 1 2370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_173
timestamp 1745462530
transform 1 0 2384 0 -1 2970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_174
timestamp 1745462530
transform 1 0 1000 0 1 2570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_175
timestamp 1745462530
transform 1 0 1696 0 -1 2970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_176
timestamp 1745462530
transform 1 0 1640 0 -1 2170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_177
timestamp 1745462530
transform 1 0 1712 0 -1 2770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_178
timestamp 1745462530
transform 1 0 1664 0 1 1970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_179
timestamp 1745462530
transform 1 0 1592 0 -1 2570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_180
timestamp 1745462530
transform 1 0 1536 0 1 1770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_181
timestamp 1745462530
transform 1 0 296 0 -1 2770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_182
timestamp 1745462530
transform 1 0 392 0 1 2570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_183
timestamp 1745462530
transform 1 0 200 0 1 2570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_184
timestamp 1745462530
transform 1 0 416 0 -1 2370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_185
timestamp 1745462530
transform 1 0 392 0 1 2170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_186
timestamp 1745462530
transform 1 0 424 0 1 1570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_187
timestamp 1745462530
transform 1 0 536 0 -1 1570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_188
timestamp 1745462530
transform 1 0 320 0 1 1370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_189
timestamp 1745462530
transform 1 0 256 0 1 770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_190
timestamp 1745462530
transform 1 0 160 0 -1 170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_191
timestamp 1745462530
transform 1 0 256 0 -1 370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_192
timestamp 1745462530
transform 1 0 416 0 -1 170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_193
timestamp 1745462530
transform 1 0 800 0 -1 170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_194
timestamp 1745462530
transform 1 0 248 0 -1 1170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_195
timestamp 1745462530
transform 1 0 656 0 -1 1570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_196
timestamp 1745462530
transform 1 0 1664 0 -1 170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_197
timestamp 1745462530
transform 1 0 1776 0 -1 370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_198
timestamp 1745462530
transform 1 0 1776 0 -1 170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_199
timestamp 1745462530
transform 1 0 1808 0 1 770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_200
timestamp 1745462530
transform 1 0 1968 0 -1 170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_201
timestamp 1745462530
transform 1 0 1888 0 1 970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_202
timestamp 1745462530
transform 1 0 1880 0 -1 1170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_203
timestamp 1745462530
transform 1 0 1856 0 -1 1370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_204
timestamp 1745462530
transform 1 0 2080 0 -1 170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_205
timestamp 1745462530
transform 1 0 2056 0 1 570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_206
timestamp 1745462530
transform 1 0 2216 0 -1 170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_207
timestamp 1745462530
transform 1 0 2088 0 1 370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_208
timestamp 1745462530
transform 1 0 2344 0 -1 170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_209
timestamp 1745462530
transform 1 0 2160 0 -1 970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_210
timestamp 1745462530
transform 1 0 2176 0 1 1170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_211
timestamp 1745462530
transform 1 0 2216 0 -1 1370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_212
timestamp 1745462530
transform 1 0 3448 0 -1 170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_213
timestamp 1745462530
transform 1 0 3792 0 -1 170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_214
timestamp 1745462530
transform 1 0 4264 0 -1 170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_215
timestamp 1745462530
transform 1 0 4040 0 -1 370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_216
timestamp 1745462530
transform 1 0 4272 0 1 170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_217
timestamp 1745462530
transform 1 0 4280 0 -1 970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_218
timestamp 1745462530
transform 1 0 4280 0 1 1170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_219
timestamp 1745462530
transform 1 0 3984 0 1 1170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_220
timestamp 1745462530
transform 1 0 4272 0 -1 1370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_221
timestamp 1745462530
transform 1 0 3616 0 -1 1370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_222
timestamp 1745462530
transform 1 0 4280 0 -1 1570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_223
timestamp 1745462530
transform 1 0 3592 0 -1 1770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_224
timestamp 1745462530
transform 1 0 4280 0 -1 1770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_225
timestamp 1745462530
transform 1 0 3280 0 -1 1970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_226
timestamp 1745462530
transform 1 0 2840 0 -1 1970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_227
timestamp 1745462530
transform 1 0 2544 0 -1 1970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_228
timestamp 1745462530
transform 1 0 4240 0 1 2570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_229
timestamp 1745462530
transform 1 0 3952 0 -1 2970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_230
timestamp 1745462530
transform 1 0 4280 0 1 2770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_231
timestamp 1745462530
transform 1 0 4280 0 -1 2970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_232
timestamp 1745462530
transform 1 0 4264 0 1 2370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_233
timestamp 1745462530
transform 1 0 4152 0 1 2170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_234
timestamp 1745462530
transform 1 0 4104 0 -1 2970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_235
timestamp 1745462530
transform 1 0 2776 0 -1 2370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_236
timestamp 1745462530
transform 1 0 2496 0 -1 2970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_237
timestamp 1745462530
transform 1 0 1112 0 -1 2970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_238
timestamp 1745462530
transform 1 0 1328 0 -1 2970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_239
timestamp 1745462530
transform 1 0 1272 0 -1 2170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_240
timestamp 1745462530
transform 1 0 1216 0 -1 2970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_241
timestamp 1745462530
transform 1 0 1296 0 1 1970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_242
timestamp 1745462530
transform 1 0 1200 0 1 2570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_243
timestamp 1745462530
transform 1 0 1224 0 1 1770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_244
timestamp 1745462530
transform 1 0 320 0 -1 2970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_245
timestamp 1745462530
transform 1 0 552 0 -1 2970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_246
timestamp 1745462530
transform 1 0 176 0 -1 2970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_247
timestamp 1745462530
transform 1 0 408 0 -1 2570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_248
timestamp 1745462530
transform 1 0 464 0 1 1970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_249
timestamp 1745462530
transform 1 0 336 0 -1 1970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_250
timestamp 1745462530
transform 1 0 792 0 1 1770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_251
timestamp 1745462530
transform 1 0 432 0 1 1370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_252
timestamp 1745462530
transform 1 0 456 0 1 970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_253
timestamp 1745462530
transform 1 0 296 0 -1 170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_254
timestamp 1745462530
transform 1 0 376 0 -1 370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_255
timestamp 1745462530
transform 1 0 680 0 -1 170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_256
timestamp 1745462530
transform 1 0 912 0 -1 170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_257
timestamp 1745462530
transform 1 0 440 0 -1 1170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_258
timestamp 1745462530
transform 1 0 560 0 1 1370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_259
timestamp 1745462530
transform 1 0 1024 0 -1 170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_260
timestamp 1745462530
transform 1 0 1488 0 -1 570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_261
timestamp 1745462530
transform 1 0 1368 0 -1 170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_262
timestamp 1745462530
transform 1 0 1280 0 1 770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_263
timestamp 1745462530
transform 1 0 1560 0 -1 170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_264
timestamp 1745462530
transform 1 0 1512 0 1 770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_265
timestamp 1745462530
transform 1 0 1544 0 -1 1170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_266
timestamp 1745462530
transform 1 0 1568 0 -1 1570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_267
timestamp 1745462530
transform 1 0 2840 0 -1 370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_268
timestamp 1745462530
transform 1 0 3136 0 -1 770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_269
timestamp 1745462530
transform 1 0 2712 0 -1 370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_270
timestamp 1745462530
transform 1 0 3064 0 -1 570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_271
timestamp 1745462530
transform 1 0 3024 0 -1 370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_272
timestamp 1745462530
transform 1 0 2896 0 1 770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_273
timestamp 1745462530
transform 1 0 2880 0 -1 1170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_274
timestamp 1745462530
transform 1 0 2912 0 1 1370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_275
timestamp 1745462530
transform 1 0 3128 0 -1 370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_276
timestamp 1745462530
transform 1 0 3104 0 1 370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_277
timestamp 1745462530
transform 1 0 4104 0 -1 570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_278
timestamp 1745462530
transform 1 0 3336 0 -1 770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_279
timestamp 1745462530
transform 1 0 4192 0 1 570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_280
timestamp 1745462530
transform 1 0 3976 0 -1 770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_281
timestamp 1745462530
transform 1 0 3248 0 -1 970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_282
timestamp 1745462530
transform 1 0 3224 0 1 1170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_283
timestamp 1745462530
transform 1 0 4064 0 -1 1370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_284
timestamp 1745462530
transform 1 0 3496 0 -1 1370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_285
timestamp 1745462530
transform 1 0 4104 0 -1 1570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_286
timestamp 1745462530
transform 1 0 3440 0 1 1570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_287
timestamp 1745462530
transform 1 0 4200 0 1 1570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_288
timestamp 1745462530
transform 1 0 3248 0 1 1570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_289
timestamp 1745462530
transform 1 0 2776 0 1 1570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_290
timestamp 1745462530
transform 1 0 2736 0 -1 1970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_291
timestamp 1745462530
transform 1 0 3152 0 -1 2770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_292
timestamp 1745462530
transform 1 0 2872 0 -1 2970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_293
timestamp 1745462530
transform 1 0 3056 0 1 2770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_294
timestamp 1745462530
transform 1 0 3072 0 1 2970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_295
timestamp 1745462530
transform 1 0 3256 0 -1 2570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_296
timestamp 1745462530
transform 1 0 3120 0 -1 2370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_297
timestamp 1745462530
transform 1 0 3048 0 -1 2970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_298
timestamp 1745462530
transform 1 0 2672 0 -1 2370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_299
timestamp 1745462530
transform 1 0 2672 0 -1 2770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_300
timestamp 1745462530
transform 1 0 1536 0 -1 2970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_301
timestamp 1745462530
transform 1 0 1536 0 -1 2170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_302
timestamp 1745462530
transform 1 0 1512 0 -1 2770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_303
timestamp 1745462530
transform 1 0 1368 0 -1 1970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_304
timestamp 1745462530
transform 1 0 1368 0 -1 2770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_305
timestamp 1745462530
transform 1 0 1328 0 -1 1770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_306
timestamp 1745462530
transform 1 0 72 0 -1 2770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_307
timestamp 1745462530
transform 1 0 464 0 -1 2770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_308
timestamp 1745462530
transform 1 0 80 0 1 2770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_309
timestamp 1745462530
transform 1 0 968 0 -1 2770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_310
timestamp 1745462530
transform 1 0 80 0 1 2370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_311
timestamp 1745462530
transform 1 0 72 0 1 1970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_312
timestamp 1745462530
transform 1 0 80 0 -1 1970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_313
timestamp 1745462530
transform 1 0 472 0 1 1770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_314
timestamp 1745462530
transform 1 0 80 0 -1 1570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_315
timestamp 1745462530
transform 1 0 256 0 -1 1370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_316
timestamp 1745462530
transform 1 0 448 0 1 170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_317
timestamp 1745462530
transform 1 0 496 0 -1 370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_318
timestamp 1745462530
transform 1 0 584 0 1 170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_319
timestamp 1745462530
transform 1 0 712 0 1 170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_320
timestamp 1745462530
transform 1 0 360 0 -1 1370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_321
timestamp 1745462530
transform 1 0 736 0 -1 1370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_322
timestamp 1745462530
transform 1 0 968 0 1 170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_323
timestamp 1745462530
transform 1 0 952 0 1 570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_324
timestamp 1745462530
transform 1 0 1240 0 1 170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_325
timestamp 1745462530
transform 1 0 1104 0 -1 770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_326
timestamp 1745462530
transform 1 0 1168 0 -1 170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_327
timestamp 1745462530
transform 1 0 1272 0 -1 970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_328
timestamp 1745462530
transform 1 0 1280 0 -1 1170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_329
timestamp 1745462530
transform 1 0 2008 0 -1 1570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_330
timestamp 1745462530
transform 1 0 2680 0 -1 170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_331
timestamp 1745462530
transform 1 0 2808 0 -1 770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_332
timestamp 1745462530
transform 1 0 2544 0 -1 170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_333
timestamp 1745462530
transform 1 0 2712 0 1 370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_334
timestamp 1745462530
transform 1 0 3000 0 -1 170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_335
timestamp 1745462530
transform 1 0 2672 0 1 770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_336
timestamp 1745462530
transform 1 0 2656 0 1 1170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_337
timestamp 1745462530
transform 1 0 2664 0 -1 1570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_338
timestamp 1745462530
transform 1 0 3224 0 -1 170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_339
timestamp 1745462530
transform 1 0 3560 0 -1 170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_340
timestamp 1745462530
transform 1 0 3672 0 -1 170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_341
timestamp 1745462530
transform 1 0 3592 0 1 170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_342
timestamp 1745462530
transform 1 0 4272 0 -1 770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_343
timestamp 1745462530
transform 1 0 4272 0 1 770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_344
timestamp 1745462530
transform 1 0 4080 0 -1 970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_345
timestamp 1745462530
transform 1 0 3584 0 -1 1170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_346
timestamp 1745462530
transform 1 0 4272 0 1 1770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_347
timestamp 1745462530
transform 1 0 3536 0 1 1770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_348
timestamp 1745462530
transform 1 0 4280 0 -1 1970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_349
timestamp 1745462530
transform 1 0 3704 0 -1 2170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_350
timestamp 1745462530
transform 1 0 4280 0 -1 2170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_351
timestamp 1745462530
transform 1 0 3632 0 1 2170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_352
timestamp 1745462530
transform 1 0 2808 0 1 1970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_353
timestamp 1745462530
transform 1 0 2608 0 1 1970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_354
timestamp 1745462530
transform 1 0 3624 0 1 2570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_355
timestamp 1745462530
transform 1 0 3560 0 1 2970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_356
timestamp 1745462530
transform 1 0 3672 0 1 2770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_357
timestamp 1745462530
transform 1 0 3592 0 -1 2970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_358
timestamp 1745462530
transform 1 0 3704 0 1 2370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_359
timestamp 1745462530
transform 1 0 3656 0 -1 2370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_360
timestamp 1745462530
transform 1 0 3456 0 1 2970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_361
timestamp 1745462530
transform 1 0 2952 0 -1 2570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_362
timestamp 1745462530
transform 1 0 2512 0 -1 2770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_363
timestamp 1745462530
transform 1 0 1904 0 1 2970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_364
timestamp 1745462530
transform 1 0 1928 0 1 2770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_365
timestamp 1745462530
transform 1 0 2040 0 1 2170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_366
timestamp 1745462530
transform 1 0 2000 0 1 2570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_367
timestamp 1745462530
transform 1 0 2072 0 1 1970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_368
timestamp 1745462530
transform 1 0 1712 0 1 2370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_369
timestamp 1745462530
transform 1 0 1720 0 1 1770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_370
timestamp 1745462530
transform 1 0 248 0 -1 2570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_371
timestamp 1745462530
transform 1 0 496 0 1 2370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_372
timestamp 1745462530
transform 1 0 80 0 -1 2570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_373
timestamp 1745462530
transform 1 0 896 0 -1 2370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_374
timestamp 1745462530
transform 1 0 272 0 1 2370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_375
timestamp 1745462530
transform 1 0 200 0 1 2170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_376
timestamp 1745462530
transform 1 0 208 0 -1 1970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_377
timestamp 1745462530
transform 1 0 520 0 -1 1970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_378
timestamp 1745462530
transform 1 0 192 0 1 1570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_379
timestamp 1745462530
transform 1 0 88 0 -1 970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_380
timestamp 1745462530
transform 1 0 136 0 -1 770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_381
timestamp 1745462530
transform 1 0 560 0 -1 570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_382
timestamp 1745462530
transform 1 0 560 0 1 370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_383
timestamp 1745462530
transform 1 0 720 0 -1 570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_384
timestamp 1745462530
transform 1 0 536 0 -1 1370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_385
timestamp 1745462530
transform 1 0 680 0 1 1170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_386
timestamp 1745462530
transform 1 0 1344 0 1 370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_387
timestamp 1745462530
transform 1 0 1736 0 -1 570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_388
timestamp 1745462530
transform 1 0 1512 0 1 370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_389
timestamp 1745462530
transform 1 0 1664 0 1 770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_390
timestamp 1745462530
transform 1 0 1704 0 1 370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_391
timestamp 1745462530
transform 1 0 1736 0 -1 970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_392
timestamp 1745462530
transform 1 0 1696 0 1 1170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_393
timestamp 1745462530
transform 1 0 1704 0 -1 1370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_394
timestamp 1745462530
transform 1 0 2896 0 -1 170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_395
timestamp 1745462530
transform 1 0 3088 0 1 570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_396
timestamp 1745462530
transform 1 0 2784 0 -1 170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_397
timestamp 1745462530
transform 1 0 2992 0 1 370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_398
timestamp 1745462530
transform 1 0 3112 0 -1 170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_399
timestamp 1745462530
transform 1 0 2944 0 -1 970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_400
timestamp 1745462530
transform 1 0 2984 0 1 1170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_401
timestamp 1745462530
transform 1 0 2880 0 -1 1370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_402
timestamp 1745462530
transform 1 0 3336 0 -1 170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_403
timestamp 1745462530
transform 1 0 3904 0 -1 170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_404
timestamp 1745462530
transform 1 0 4128 0 -1 170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_405
timestamp 1745462530
transform 1 0 4024 0 -1 170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_406
timestamp 1745462530
transform 1 0 4152 0 -1 370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_407
timestamp 1745462530
transform 1 0 4272 0 -1 1170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_408
timestamp 1745462530
transform 1 0 4176 0 -1 1170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_409
timestamp 1745462530
transform 1 0 4080 0 1 1170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_410
timestamp 1745462530
transform 1 0 4152 0 -1 1770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_411
timestamp 1745462530
transform 1 0 3952 0 1 1770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_412
timestamp 1745462530
transform 1 0 4272 0 1 2170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_413
timestamp 1745462530
transform 1 0 4000 0 1 1970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_414
timestamp 1745462530
transform 1 0 4184 0 -1 2170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_415
timestamp 1745462530
transform 1 0 3944 0 1 2170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_416
timestamp 1745462530
transform 1 0 3184 0 1 2170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_417
timestamp 1745462530
transform 1 0 2992 0 1 2170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_418
timestamp 1745462530
transform 1 0 4232 0 -1 2770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_419
timestamp 1745462530
transform 1 0 3984 0 1 2970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_420
timestamp 1745462530
transform 1 0 4176 0 1 2770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_421
timestamp 1745462530
transform 1 0 4240 0 1 2970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_422
timestamp 1745462530
transform 1 0 4272 0 -1 2570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_423
timestamp 1745462530
transform 1 0 4280 0 -1 2370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_424
timestamp 1745462530
transform 1 0 4072 0 -1 3170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_425
timestamp 1745462530
transform 1 0 2880 0 -1 2770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_426
timestamp 1745462530
transform 1 0 2760 0 -1 2970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_427
timestamp 1745462530
transform 1 0 3008 0 1 3770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_428
timestamp 1745462530
transform 1 0 1336 0 1 3770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_429
timestamp 1745462530
transform 1 0 2776 0 1 3770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_430
timestamp 1745462530
transform 1 0 1448 0 1 3770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_431
timestamp 1745462530
transform 1 0 3896 0 -1 3770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_432
timestamp 1745462530
transform 1 0 4104 0 -1 3370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_433
timestamp 1745462530
transform 1 0 4272 0 1 3170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_434
timestamp 1745462530
transform 1 0 4272 0 -1 3170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_435
timestamp 1745462530
transform 1 0 1488 0 1 3970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_436
timestamp 1745462530
transform 1 0 1608 0 -1 4170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_437
timestamp 1745462530
transform 1 0 1376 0 -1 3970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_438
timestamp 1745462530
transform 1 0 1504 0 -1 3970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_439
timestamp 1745462530
transform 1 0 3912 0 -1 3370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_440
timestamp 1745462530
transform 1 0 4088 0 1 3170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_441
timestamp 1745462530
transform 1 0 4280 0 1 3370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_442
timestamp 1745462530
transform 1 0 4280 0 -1 3370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_443
timestamp 1745462530
transform 1 0 1736 0 -1 4170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_444
timestamp 1745462530
transform 1 0 1816 0 1 3970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_445
timestamp 1745462530
transform 1 0 1920 0 -1 4170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_446
timestamp 1745462530
transform 1 0 1904 0 1 3570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_447
timestamp 1745462530
transform 1 0 4032 0 1 3370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_448
timestamp 1745462530
transform 1 0 4272 0 -1 3570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_449
timestamp 1745462530
transform 1 0 4104 0 1 3570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_450
timestamp 1745462530
transform 1 0 4152 0 -1 3570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_451
timestamp 1745462530
transform 1 0 2904 0 1 3770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_452
timestamp 1745462530
transform 1 0 2568 0 -1 3970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_453
timestamp 1745462530
transform 1 0 1968 0 1 3970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_454
timestamp 1745462530
transform 1 0 1896 0 1 3770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_455
timestamp 1745462530
transform 1 0 3920 0 1 3570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_456
timestamp 1745462530
transform 1 0 4280 0 1 3570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_457
timestamp 1745462530
transform 1 0 4272 0 -1 3970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_458
timestamp 1745462530
transform 1 0 4280 0 1 3770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_459
timestamp 1745462530
transform 1 0 2856 0 1 3970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_460
timestamp 1745462530
transform 1 0 2544 0 -1 4170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_461
timestamp 1745462530
transform 1 0 2200 0 1 4170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_462
timestamp 1745462530
transform 1 0 2432 0 1 4170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_463
timestamp 1745462530
transform 1 0 3720 0 1 4170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_464
timestamp 1745462530
transform 1 0 3752 0 -1 3970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_465
timestamp 1745462530
transform 1 0 3912 0 1 4170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_466
timestamp 1745462530
transform 1 0 3832 0 1 3970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_467
timestamp 1745462530
transform 1 0 2896 0 -1 4170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_468
timestamp 1745462530
transform 1 0 2712 0 1 4170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_469
timestamp 1745462530
transform 1 0 2024 0 1 4170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_470
timestamp 1745462530
transform 1 0 2336 0 1 4170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_471
timestamp 1745462530
transform 1 0 3184 0 1 4170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_472
timestamp 1745462530
transform 1 0 3624 0 1 3970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_473
timestamp 1745462530
transform 1 0 3376 0 1 4170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_474
timestamp 1745462530
transform 1 0 3528 0 1 4170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_475
timestamp 1745462530
transform 1 0 3088 0 1 4170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_476
timestamp 1745462530
transform 1 0 2800 0 -1 4170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_477
timestamp 1745462530
transform 1 0 2240 0 1 3970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_478
timestamp 1745462530
transform 1 0 2448 0 1 3970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_479
timestamp 1745462530
transform 1 0 3280 0 1 4170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_480
timestamp 1745462530
transform 1 0 3712 0 1 3770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_481
timestamp 1745462530
transform 1 0 3624 0 1 4170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_482
timestamp 1745462530
transform 1 0 3824 0 1 3770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_483
timestamp 1745462530
transform 1 0 3072 0 -1 4170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_484
timestamp 1745462530
transform 1 0 2736 0 1 3970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_485
timestamp 1745462530
transform 1 0 2056 0 -1 4170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_486
timestamp 1745462530
transform 1 0 2448 0 -1 3970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_487
timestamp 1745462530
transform 1 0 3112 0 1 3970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_488
timestamp 1745462530
transform 1 0 3240 0 1 3770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_489
timestamp 1745462530
transform 1 0 3232 0 1 3970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_490
timestamp 1745462530
transform 1 0 3344 0 1 3970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_491
timestamp 1745462530
transform 1 0 984 0 1 3770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_492
timestamp 1745462530
transform 1 0 856 0 1 3770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_493
timestamp 1745462530
transform 1 0 232 0 1 4170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_494
timestamp 1745462530
transform 1 0 352 0 -1 4170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_495
timestamp 1745462530
transform 1 0 344 0 1 4170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_496
timestamp 1745462530
transform 1 0 224 0 -1 4170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_497
timestamp 1745462530
transform 1 0 336 0 -1 3970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_498
timestamp 1745462530
transform 1 0 192 0 -1 3970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_499
timestamp 1745462530
transform 1 0 368 0 1 3770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_500
timestamp 1745462530
transform 1 0 248 0 1 3770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_501
timestamp 1745462530
transform 1 0 544 0 -1 3770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_502
timestamp 1745462530
transform 1 0 512 0 1 3770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_503
timestamp 1745462530
transform 1 0 632 0 -1 3970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_504
timestamp 1745462530
transform 1 0 944 0 1 3970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_505
timestamp 1745462530
transform 1 0 816 0 1 4170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_506
timestamp 1745462530
transform 1 0 912 0 1 4170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_507
timestamp 1745462530
transform 1 0 488 0 -1 4170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_508
timestamp 1745462530
transform 1 0 456 0 1 4170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_509
timestamp 1745462530
transform 1 0 640 0 1 3770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_510
timestamp 1745462530
transform 1 0 808 0 -1 3970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_511
timestamp 1745462530
transform 1 0 736 0 1 3970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_512
timestamp 1745462530
transform 1 0 720 0 1 4170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_513
timestamp 1745462530
transform 1 0 928 0 -1 3970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_514
timestamp 1745462530
transform 1 0 1096 0 -1 3970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_515
timestamp 1745462530
transform 1 0 1008 0 1 4170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_516
timestamp 1745462530
transform 1 0 1104 0 1 4170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_517
timestamp 1745462530
transform 1 0 1208 0 -1 3970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_518
timestamp 1745462530
transform 1 0 1200 0 1 4170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_519
timestamp 1745462530
transform 1 0 1248 0 -1 4170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_520
timestamp 1745462530
transform 1 0 1296 0 1 4170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_521
timestamp 1745462530
transform 1 0 1392 0 1 4170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_522
timestamp 1745462530
transform 1 0 4168 0 1 4170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_523
timestamp 1745462530
transform 1 0 4272 0 1 3970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_524
timestamp 1745462530
transform 1 0 4272 0 1 4170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_525
timestamp 1745462530
transform 1 0 4280 0 -1 4170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_526
timestamp 1745462530
transform 1 0 1544 0 1 4170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_527
timestamp 1745462530
transform 1 0 1640 0 1 4170
box -8 -3 104 105
use FILL  FILL_0
timestamp 1745462530
transform 1 0 4368 0 1 4170
box -8 -3 16 105
use FILL  FILL_1
timestamp 1745462530
transform 1 0 4264 0 1 4170
box -8 -3 16 105
use FILL  FILL_2
timestamp 1745462530
transform 1 0 4160 0 1 4170
box -8 -3 16 105
use FILL  FILL_3
timestamp 1745462530
transform 1 0 712 0 1 4170
box -8 -3 16 105
use FILL  FILL_4
timestamp 1745462530
transform 1 0 704 0 1 4170
box -8 -3 16 105
use FILL  FILL_5
timestamp 1745462530
transform 1 0 648 0 1 4170
box -8 -3 16 105
use FILL  FILL_6
timestamp 1745462530
transform 1 0 552 0 1 4170
box -8 -3 16 105
use FILL  FILL_7
timestamp 1745462530
transform 1 0 448 0 1 4170
box -8 -3 16 105
use FILL  FILL_8
timestamp 1745462530
transform 1 0 440 0 1 4170
box -8 -3 16 105
use FILL  FILL_9
timestamp 1745462530
transform 1 0 336 0 1 4170
box -8 -3 16 105
use FILL  FILL_10
timestamp 1745462530
transform 1 0 328 0 1 4170
box -8 -3 16 105
use FILL  FILL_11
timestamp 1745462530
transform 1 0 224 0 1 4170
box -8 -3 16 105
use FILL  FILL_12
timestamp 1745462530
transform 1 0 216 0 1 4170
box -8 -3 16 105
use FILL  FILL_13
timestamp 1745462530
transform 1 0 160 0 1 4170
box -8 -3 16 105
use FILL  FILL_14
timestamp 1745462530
transform 1 0 112 0 1 4170
box -8 -3 16 105
use FILL  FILL_15
timestamp 1745462530
transform 1 0 72 0 1 4170
box -8 -3 16 105
use FILL  FILL_16
timestamp 1745462530
transform 1 0 4272 0 -1 4170
box -8 -3 16 105
use FILL  FILL_17
timestamp 1745462530
transform 1 0 4208 0 -1 4170
box -8 -3 16 105
use FILL  FILL_18
timestamp 1745462530
transform 1 0 4168 0 -1 4170
box -8 -3 16 105
use FILL  FILL_19
timestamp 1745462530
transform 1 0 4104 0 -1 4170
box -8 -3 16 105
use FILL  FILL_20
timestamp 1745462530
transform 1 0 3976 0 -1 4170
box -8 -3 16 105
use FILL  FILL_21
timestamp 1745462530
transform 1 0 3912 0 -1 4170
box -8 -3 16 105
use FILL  FILL_22
timestamp 1745462530
transform 1 0 3904 0 -1 4170
box -8 -3 16 105
use FILL  FILL_23
timestamp 1745462530
transform 1 0 3760 0 -1 4170
box -8 -3 16 105
use FILL  FILL_24
timestamp 1745462530
transform 1 0 3680 0 -1 4170
box -8 -3 16 105
use FILL  FILL_25
timestamp 1745462530
transform 1 0 3576 0 -1 4170
box -8 -3 16 105
use FILL  FILL_26
timestamp 1745462530
transform 1 0 3416 0 -1 4170
box -8 -3 16 105
use FILL  FILL_27
timestamp 1745462530
transform 1 0 3280 0 -1 4170
box -8 -3 16 105
use FILL  FILL_28
timestamp 1745462530
transform 1 0 3064 0 -1 4170
box -8 -3 16 105
use FILL  FILL_29
timestamp 1745462530
transform 1 0 2792 0 -1 4170
box -8 -3 16 105
use FILL  FILL_30
timestamp 1745462530
transform 1 0 2696 0 -1 4170
box -8 -3 16 105
use FILL  FILL_31
timestamp 1745462530
transform 1 0 2536 0 -1 4170
box -8 -3 16 105
use FILL  FILL_32
timestamp 1745462530
transform 1 0 2456 0 -1 4170
box -8 -3 16 105
use FILL  FILL_33
timestamp 1745462530
transform 1 0 2392 0 -1 4170
box -8 -3 16 105
use FILL  FILL_34
timestamp 1745462530
transform 1 0 1600 0 -1 4170
box -8 -3 16 105
use FILL  FILL_35
timestamp 1745462530
transform 1 0 1520 0 -1 4170
box -8 -3 16 105
use FILL  FILL_36
timestamp 1745462530
transform 1 0 1392 0 -1 4170
box -8 -3 16 105
use FILL  FILL_37
timestamp 1745462530
transform 1 0 1192 0 -1 4170
box -8 -3 16 105
use FILL  FILL_38
timestamp 1745462530
transform 1 0 1136 0 -1 4170
box -8 -3 16 105
use FILL  FILL_39
timestamp 1745462530
transform 1 0 1104 0 -1 4170
box -8 -3 16 105
use FILL  FILL_40
timestamp 1745462530
transform 1 0 1024 0 -1 4170
box -8 -3 16 105
use FILL  FILL_41
timestamp 1745462530
transform 1 0 960 0 -1 4170
box -8 -3 16 105
use FILL  FILL_42
timestamp 1745462530
transform 1 0 824 0 -1 4170
box -8 -3 16 105
use FILL  FILL_43
timestamp 1745462530
transform 1 0 744 0 -1 4170
box -8 -3 16 105
use FILL  FILL_44
timestamp 1745462530
transform 1 0 680 0 -1 4170
box -8 -3 16 105
use FILL  FILL_45
timestamp 1745462530
transform 1 0 600 0 -1 4170
box -8 -3 16 105
use FILL  FILL_46
timestamp 1745462530
transform 1 0 216 0 -1 4170
box -8 -3 16 105
use FILL  FILL_47
timestamp 1745462530
transform 1 0 4368 0 1 3970
box -8 -3 16 105
use FILL  FILL_48
timestamp 1745462530
transform 1 0 4264 0 1 3970
box -8 -3 16 105
use FILL  FILL_49
timestamp 1745462530
transform 1 0 4256 0 1 3970
box -8 -3 16 105
use FILL  FILL_50
timestamp 1745462530
transform 1 0 4192 0 1 3970
box -8 -3 16 105
use FILL  FILL_51
timestamp 1745462530
transform 1 0 4152 0 1 3970
box -8 -3 16 105
use FILL  FILL_52
timestamp 1745462530
transform 1 0 4144 0 1 3970
box -8 -3 16 105
use FILL  FILL_53
timestamp 1745462530
transform 1 0 4088 0 1 3970
box -8 -3 16 105
use FILL  FILL_54
timestamp 1745462530
transform 1 0 4080 0 1 3970
box -8 -3 16 105
use FILL  FILL_55
timestamp 1745462530
transform 1 0 4040 0 1 3970
box -8 -3 16 105
use FILL  FILL_56
timestamp 1745462530
transform 1 0 4000 0 1 3970
box -8 -3 16 105
use FILL  FILL_57
timestamp 1745462530
transform 1 0 3992 0 1 3970
box -8 -3 16 105
use FILL  FILL_58
timestamp 1745462530
transform 1 0 3984 0 1 3970
box -8 -3 16 105
use FILL  FILL_59
timestamp 1745462530
transform 1 0 3944 0 1 3970
box -8 -3 16 105
use FILL  FILL_60
timestamp 1745462530
transform 1 0 3936 0 1 3970
box -8 -3 16 105
use FILL  FILL_61
timestamp 1745462530
transform 1 0 3928 0 1 3970
box -8 -3 16 105
use FILL  FILL_62
timestamp 1745462530
transform 1 0 3824 0 1 3970
box -8 -3 16 105
use FILL  FILL_63
timestamp 1745462530
transform 1 0 3816 0 1 3970
box -8 -3 16 105
use FILL  FILL_64
timestamp 1745462530
transform 1 0 3792 0 1 3970
box -8 -3 16 105
use FILL  FILL_65
timestamp 1745462530
transform 1 0 3728 0 1 3970
box -8 -3 16 105
use FILL  FILL_66
timestamp 1745462530
transform 1 0 3720 0 1 3970
box -8 -3 16 105
use FILL  FILL_67
timestamp 1745462530
transform 1 0 3616 0 1 3970
box -8 -3 16 105
use FILL  FILL_68
timestamp 1745462530
transform 1 0 3608 0 1 3970
box -8 -3 16 105
use FILL  FILL_69
timestamp 1745462530
transform 1 0 3600 0 1 3970
box -8 -3 16 105
use FILL  FILL_70
timestamp 1745462530
transform 1 0 3536 0 1 3970
box -8 -3 16 105
use FILL  FILL_71
timestamp 1745462530
transform 1 0 3488 0 1 3970
box -8 -3 16 105
use FILL  FILL_72
timestamp 1745462530
transform 1 0 3448 0 1 3970
box -8 -3 16 105
use FILL  FILL_73
timestamp 1745462530
transform 1 0 3440 0 1 3970
box -8 -3 16 105
use FILL  FILL_74
timestamp 1745462530
transform 1 0 3336 0 1 3970
box -8 -3 16 105
use FILL  FILL_75
timestamp 1745462530
transform 1 0 3328 0 1 3970
box -8 -3 16 105
use FILL  FILL_76
timestamp 1745462530
transform 1 0 3224 0 1 3970
box -8 -3 16 105
use FILL  FILL_77
timestamp 1745462530
transform 1 0 3216 0 1 3970
box -8 -3 16 105
use FILL  FILL_78
timestamp 1745462530
transform 1 0 3208 0 1 3970
box -8 -3 16 105
use FILL  FILL_79
timestamp 1745462530
transform 1 0 3104 0 1 3970
box -8 -3 16 105
use FILL  FILL_80
timestamp 1745462530
transform 1 0 3096 0 1 3970
box -8 -3 16 105
use FILL  FILL_81
timestamp 1745462530
transform 1 0 3032 0 1 3970
box -8 -3 16 105
use FILL  FILL_82
timestamp 1745462530
transform 1 0 3024 0 1 3970
box -8 -3 16 105
use FILL  FILL_83
timestamp 1745462530
transform 1 0 3016 0 1 3970
box -8 -3 16 105
use FILL  FILL_84
timestamp 1745462530
transform 1 0 2952 0 1 3970
box -8 -3 16 105
use FILL  FILL_85
timestamp 1745462530
transform 1 0 2848 0 1 3970
box -8 -3 16 105
use FILL  FILL_86
timestamp 1745462530
transform 1 0 2840 0 1 3970
box -8 -3 16 105
use FILL  FILL_87
timestamp 1745462530
transform 1 0 2832 0 1 3970
box -8 -3 16 105
use FILL  FILL_88
timestamp 1745462530
transform 1 0 2728 0 1 3970
box -8 -3 16 105
use FILL  FILL_89
timestamp 1745462530
transform 1 0 2704 0 1 3970
box -8 -3 16 105
use FILL  FILL_90
timestamp 1745462530
transform 1 0 2656 0 1 3970
box -8 -3 16 105
use FILL  FILL_91
timestamp 1745462530
transform 1 0 2648 0 1 3970
box -8 -3 16 105
use FILL  FILL_92
timestamp 1745462530
transform 1 0 2624 0 1 3970
box -8 -3 16 105
use FILL  FILL_93
timestamp 1745462530
transform 1 0 2576 0 1 3970
box -8 -3 16 105
use FILL  FILL_94
timestamp 1745462530
transform 1 0 2552 0 1 3970
box -8 -3 16 105
use FILL  FILL_95
timestamp 1745462530
transform 1 0 2544 0 1 3970
box -8 -3 16 105
use FILL  FILL_96
timestamp 1745462530
transform 1 0 2440 0 1 3970
box -8 -3 16 105
use FILL  FILL_97
timestamp 1745462530
transform 1 0 2432 0 1 3970
box -8 -3 16 105
use FILL  FILL_98
timestamp 1745462530
transform 1 0 2424 0 1 3970
box -8 -3 16 105
use FILL  FILL_99
timestamp 1745462530
transform 1 0 2344 0 1 3970
box -8 -3 16 105
use FILL  FILL_100
timestamp 1745462530
transform 1 0 2336 0 1 3970
box -8 -3 16 105
use FILL  FILL_101
timestamp 1745462530
transform 1 0 2232 0 1 3970
box -8 -3 16 105
use FILL  FILL_102
timestamp 1745462530
transform 1 0 2224 0 1 3970
box -8 -3 16 105
use FILL  FILL_103
timestamp 1745462530
transform 1 0 2216 0 1 3970
box -8 -3 16 105
use FILL  FILL_104
timestamp 1745462530
transform 1 0 2192 0 1 3970
box -8 -3 16 105
use FILL  FILL_105
timestamp 1745462530
transform 1 0 2144 0 1 3970
box -8 -3 16 105
use FILL  FILL_106
timestamp 1745462530
transform 1 0 2136 0 1 3970
box -8 -3 16 105
use FILL  FILL_107
timestamp 1745462530
transform 1 0 2128 0 1 3970
box -8 -3 16 105
use FILL  FILL_108
timestamp 1745462530
transform 1 0 2080 0 1 3970
box -8 -3 16 105
use FILL  FILL_109
timestamp 1745462530
transform 1 0 2072 0 1 3970
box -8 -3 16 105
use FILL  FILL_110
timestamp 1745462530
transform 1 0 2064 0 1 3970
box -8 -3 16 105
use FILL  FILL_111
timestamp 1745462530
transform 1 0 1960 0 1 3970
box -8 -3 16 105
use FILL  FILL_112
timestamp 1745462530
transform 1 0 1952 0 1 3970
box -8 -3 16 105
use FILL  FILL_113
timestamp 1745462530
transform 1 0 1928 0 1 3970
box -8 -3 16 105
use FILL  FILL_114
timestamp 1745462530
transform 1 0 1920 0 1 3970
box -8 -3 16 105
use FILL  FILL_115
timestamp 1745462530
transform 1 0 1912 0 1 3970
box -8 -3 16 105
use FILL  FILL_116
timestamp 1745462530
transform 1 0 1808 0 1 3970
box -8 -3 16 105
use FILL  FILL_117
timestamp 1745462530
transform 1 0 1800 0 1 3970
box -8 -3 16 105
use FILL  FILL_118
timestamp 1745462530
transform 1 0 1792 0 1 3970
box -8 -3 16 105
use FILL  FILL_119
timestamp 1745462530
transform 1 0 1784 0 1 3970
box -8 -3 16 105
use FILL  FILL_120
timestamp 1745462530
transform 1 0 1728 0 1 3970
box -8 -3 16 105
use FILL  FILL_121
timestamp 1745462530
transform 1 0 1720 0 1 3970
box -8 -3 16 105
use FILL  FILL_122
timestamp 1745462530
transform 1 0 1672 0 1 3970
box -8 -3 16 105
use FILL  FILL_123
timestamp 1745462530
transform 1 0 1664 0 1 3970
box -8 -3 16 105
use FILL  FILL_124
timestamp 1745462530
transform 1 0 1656 0 1 3970
box -8 -3 16 105
use FILL  FILL_125
timestamp 1745462530
transform 1 0 1648 0 1 3970
box -8 -3 16 105
use FILL  FILL_126
timestamp 1745462530
transform 1 0 1600 0 1 3970
box -8 -3 16 105
use FILL  FILL_127
timestamp 1745462530
transform 1 0 1592 0 1 3970
box -8 -3 16 105
use FILL  FILL_128
timestamp 1745462530
transform 1 0 1584 0 1 3970
box -8 -3 16 105
use FILL  FILL_129
timestamp 1745462530
transform 1 0 1480 0 1 3970
box -8 -3 16 105
use FILL  FILL_130
timestamp 1745462530
transform 1 0 1472 0 1 3970
box -8 -3 16 105
use FILL  FILL_131
timestamp 1745462530
transform 1 0 1464 0 1 3970
box -8 -3 16 105
use FILL  FILL_132
timestamp 1745462530
transform 1 0 1456 0 1 3970
box -8 -3 16 105
use FILL  FILL_133
timestamp 1745462530
transform 1 0 1448 0 1 3970
box -8 -3 16 105
use FILL  FILL_134
timestamp 1745462530
transform 1 0 1440 0 1 3970
box -8 -3 16 105
use FILL  FILL_135
timestamp 1745462530
transform 1 0 1432 0 1 3970
box -8 -3 16 105
use FILL  FILL_136
timestamp 1745462530
transform 1 0 1424 0 1 3970
box -8 -3 16 105
use FILL  FILL_137
timestamp 1745462530
transform 1 0 1416 0 1 3970
box -8 -3 16 105
use FILL  FILL_138
timestamp 1745462530
transform 1 0 1408 0 1 3970
box -8 -3 16 105
use FILL  FILL_139
timestamp 1745462530
transform 1 0 1400 0 1 3970
box -8 -3 16 105
use FILL  FILL_140
timestamp 1745462530
transform 1 0 1392 0 1 3970
box -8 -3 16 105
use FILL  FILL_141
timestamp 1745462530
transform 1 0 1384 0 1 3970
box -8 -3 16 105
use FILL  FILL_142
timestamp 1745462530
transform 1 0 1360 0 1 3970
box -8 -3 16 105
use FILL  FILL_143
timestamp 1745462530
transform 1 0 1336 0 1 3970
box -8 -3 16 105
use FILL  FILL_144
timestamp 1745462530
transform 1 0 1328 0 1 3970
box -8 -3 16 105
use FILL  FILL_145
timestamp 1745462530
transform 1 0 1320 0 1 3970
box -8 -3 16 105
use FILL  FILL_146
timestamp 1745462530
transform 1 0 1312 0 1 3970
box -8 -3 16 105
use FILL  FILL_147
timestamp 1745462530
transform 1 0 1280 0 1 3970
box -8 -3 16 105
use FILL  FILL_148
timestamp 1745462530
transform 1 0 1240 0 1 3970
box -8 -3 16 105
use FILL  FILL_149
timestamp 1745462530
transform 1 0 1232 0 1 3970
box -8 -3 16 105
use FILL  FILL_150
timestamp 1745462530
transform 1 0 1192 0 1 3970
box -8 -3 16 105
use FILL  FILL_151
timestamp 1745462530
transform 1 0 1184 0 1 3970
box -8 -3 16 105
use FILL  FILL_152
timestamp 1745462530
transform 1 0 1152 0 1 3970
box -8 -3 16 105
use FILL  FILL_153
timestamp 1745462530
transform 1 0 1120 0 1 3970
box -8 -3 16 105
use FILL  FILL_154
timestamp 1745462530
transform 1 0 1112 0 1 3970
box -8 -3 16 105
use FILL  FILL_155
timestamp 1745462530
transform 1 0 1104 0 1 3970
box -8 -3 16 105
use FILL  FILL_156
timestamp 1745462530
transform 1 0 1048 0 1 3970
box -8 -3 16 105
use FILL  FILL_157
timestamp 1745462530
transform 1 0 1040 0 1 3970
box -8 -3 16 105
use FILL  FILL_158
timestamp 1745462530
transform 1 0 936 0 1 3970
box -8 -3 16 105
use FILL  FILL_159
timestamp 1745462530
transform 1 0 928 0 1 3970
box -8 -3 16 105
use FILL  FILL_160
timestamp 1745462530
transform 1 0 920 0 1 3970
box -8 -3 16 105
use FILL  FILL_161
timestamp 1745462530
transform 1 0 872 0 1 3970
box -8 -3 16 105
use FILL  FILL_162
timestamp 1745462530
transform 1 0 840 0 1 3970
box -8 -3 16 105
use FILL  FILL_163
timestamp 1745462530
transform 1 0 832 0 1 3970
box -8 -3 16 105
use FILL  FILL_164
timestamp 1745462530
transform 1 0 728 0 1 3970
box -8 -3 16 105
use FILL  FILL_165
timestamp 1745462530
transform 1 0 720 0 1 3970
box -8 -3 16 105
use FILL  FILL_166
timestamp 1745462530
transform 1 0 680 0 1 3970
box -8 -3 16 105
use FILL  FILL_167
timestamp 1745462530
transform 1 0 624 0 1 3970
box -8 -3 16 105
use FILL  FILL_168
timestamp 1745462530
transform 1 0 616 0 1 3970
box -8 -3 16 105
use FILL  FILL_169
timestamp 1745462530
transform 1 0 608 0 1 3970
box -8 -3 16 105
use FILL  FILL_170
timestamp 1745462530
transform 1 0 552 0 1 3970
box -8 -3 16 105
use FILL  FILL_171
timestamp 1745462530
transform 1 0 472 0 1 3970
box -8 -3 16 105
use FILL  FILL_172
timestamp 1745462530
transform 1 0 416 0 1 3970
box -8 -3 16 105
use FILL  FILL_173
timestamp 1745462530
transform 1 0 376 0 1 3970
box -8 -3 16 105
use FILL  FILL_174
timestamp 1745462530
transform 1 0 368 0 1 3970
box -8 -3 16 105
use FILL  FILL_175
timestamp 1745462530
transform 1 0 296 0 1 3970
box -8 -3 16 105
use FILL  FILL_176
timestamp 1745462530
transform 1 0 256 0 1 3970
box -8 -3 16 105
use FILL  FILL_177
timestamp 1745462530
transform 1 0 248 0 1 3970
box -8 -3 16 105
use FILL  FILL_178
timestamp 1745462530
transform 1 0 208 0 1 3970
box -8 -3 16 105
use FILL  FILL_179
timestamp 1745462530
transform 1 0 160 0 1 3970
box -8 -3 16 105
use FILL  FILL_180
timestamp 1745462530
transform 1 0 128 0 1 3970
box -8 -3 16 105
use FILL  FILL_181
timestamp 1745462530
transform 1 0 72 0 1 3970
box -8 -3 16 105
use FILL  FILL_182
timestamp 1745462530
transform 1 0 4368 0 -1 3970
box -8 -3 16 105
use FILL  FILL_183
timestamp 1745462530
transform 1 0 4264 0 -1 3970
box -8 -3 16 105
use FILL  FILL_184
timestamp 1745462530
transform 1 0 4256 0 -1 3970
box -8 -3 16 105
use FILL  FILL_185
timestamp 1745462530
transform 1 0 4192 0 -1 3970
box -8 -3 16 105
use FILL  FILL_186
timestamp 1745462530
transform 1 0 4152 0 -1 3970
box -8 -3 16 105
use FILL  FILL_187
timestamp 1745462530
transform 1 0 4120 0 -1 3970
box -8 -3 16 105
use FILL  FILL_188
timestamp 1745462530
transform 1 0 4064 0 -1 3970
box -8 -3 16 105
use FILL  FILL_189
timestamp 1745462530
transform 1 0 4024 0 -1 3970
box -8 -3 16 105
use FILL  FILL_190
timestamp 1745462530
transform 1 0 3984 0 -1 3970
box -8 -3 16 105
use FILL  FILL_191
timestamp 1745462530
transform 1 0 3976 0 -1 3970
box -8 -3 16 105
use FILL  FILL_192
timestamp 1745462530
transform 1 0 3920 0 -1 3970
box -8 -3 16 105
use FILL  FILL_193
timestamp 1745462530
transform 1 0 3912 0 -1 3970
box -8 -3 16 105
use FILL  FILL_194
timestamp 1745462530
transform 1 0 3856 0 -1 3970
box -8 -3 16 105
use FILL  FILL_195
timestamp 1745462530
transform 1 0 3848 0 -1 3970
box -8 -3 16 105
use FILL  FILL_196
timestamp 1745462530
transform 1 0 3744 0 -1 3970
box -8 -3 16 105
use FILL  FILL_197
timestamp 1745462530
transform 1 0 3720 0 -1 3970
box -8 -3 16 105
use FILL  FILL_198
timestamp 1745462530
transform 1 0 3656 0 -1 3970
box -8 -3 16 105
use FILL  FILL_199
timestamp 1745462530
transform 1 0 3648 0 -1 3970
box -8 -3 16 105
use FILL  FILL_200
timestamp 1745462530
transform 1 0 3584 0 -1 3970
box -8 -3 16 105
use FILL  FILL_201
timestamp 1745462530
transform 1 0 3536 0 -1 3970
box -8 -3 16 105
use FILL  FILL_202
timestamp 1745462530
transform 1 0 3496 0 -1 3970
box -8 -3 16 105
use FILL  FILL_203
timestamp 1745462530
transform 1 0 3432 0 -1 3970
box -8 -3 16 105
use FILL  FILL_204
timestamp 1745462530
transform 1 0 3424 0 -1 3970
box -8 -3 16 105
use FILL  FILL_205
timestamp 1745462530
transform 1 0 3416 0 -1 3970
box -8 -3 16 105
use FILL  FILL_206
timestamp 1745462530
transform 1 0 3352 0 -1 3970
box -8 -3 16 105
use FILL  FILL_207
timestamp 1745462530
transform 1 0 3344 0 -1 3970
box -8 -3 16 105
use FILL  FILL_208
timestamp 1745462530
transform 1 0 3280 0 -1 3970
box -8 -3 16 105
use FILL  FILL_209
timestamp 1745462530
transform 1 0 3216 0 -1 3970
box -8 -3 16 105
use FILL  FILL_210
timestamp 1745462530
transform 1 0 3208 0 -1 3970
box -8 -3 16 105
use FILL  FILL_211
timestamp 1745462530
transform 1 0 3144 0 -1 3970
box -8 -3 16 105
use FILL  FILL_212
timestamp 1745462530
transform 1 0 3136 0 -1 3970
box -8 -3 16 105
use FILL  FILL_213
timestamp 1745462530
transform 1 0 3072 0 -1 3970
box -8 -3 16 105
use FILL  FILL_214
timestamp 1745462530
transform 1 0 2984 0 -1 3970
box -8 -3 16 105
use FILL  FILL_215
timestamp 1745462530
transform 1 0 2976 0 -1 3970
box -8 -3 16 105
use FILL  FILL_216
timestamp 1745462530
transform 1 0 2968 0 -1 3970
box -8 -3 16 105
use FILL  FILL_217
timestamp 1745462530
transform 1 0 2888 0 -1 3970
box -8 -3 16 105
use FILL  FILL_218
timestamp 1745462530
transform 1 0 2824 0 -1 3970
box -8 -3 16 105
use FILL  FILL_219
timestamp 1745462530
transform 1 0 2800 0 -1 3970
box -8 -3 16 105
use FILL  FILL_220
timestamp 1745462530
transform 1 0 2752 0 -1 3970
box -8 -3 16 105
use FILL  FILL_221
timestamp 1745462530
transform 1 0 2664 0 -1 3970
box -8 -3 16 105
use FILL  FILL_222
timestamp 1745462530
transform 1 0 2544 0 -1 3970
box -8 -3 16 105
use FILL  FILL_223
timestamp 1745462530
transform 1 0 2440 0 -1 3970
box -8 -3 16 105
use FILL  FILL_224
timestamp 1745462530
transform 1 0 2432 0 -1 3970
box -8 -3 16 105
use FILL  FILL_225
timestamp 1745462530
transform 1 0 2264 0 -1 3970
box -8 -3 16 105
use FILL  FILL_226
timestamp 1745462530
transform 1 0 2176 0 -1 3970
box -8 -3 16 105
use FILL  FILL_227
timestamp 1745462530
transform 1 0 2120 0 -1 3970
box -8 -3 16 105
use FILL  FILL_228
timestamp 1745462530
transform 1 0 1984 0 -1 3970
box -8 -3 16 105
use FILL  FILL_229
timestamp 1745462530
transform 1 0 1976 0 -1 3970
box -8 -3 16 105
use FILL  FILL_230
timestamp 1745462530
transform 1 0 1912 0 -1 3970
box -8 -3 16 105
use FILL  FILL_231
timestamp 1745462530
transform 1 0 1832 0 -1 3970
box -8 -3 16 105
use FILL  FILL_232
timestamp 1745462530
transform 1 0 1768 0 -1 3970
box -8 -3 16 105
use FILL  FILL_233
timestamp 1745462530
transform 1 0 1760 0 -1 3970
box -8 -3 16 105
use FILL  FILL_234
timestamp 1745462530
transform 1 0 1696 0 -1 3970
box -8 -3 16 105
use FILL  FILL_235
timestamp 1745462530
transform 1 0 1496 0 -1 3970
box -8 -3 16 105
use FILL  FILL_236
timestamp 1745462530
transform 1 0 1472 0 -1 3970
box -8 -3 16 105
use FILL  FILL_237
timestamp 1745462530
transform 1 0 1368 0 -1 3970
box -8 -3 16 105
use FILL  FILL_238
timestamp 1745462530
transform 1 0 1312 0 -1 3970
box -8 -3 16 105
use FILL  FILL_239
timestamp 1745462530
transform 1 0 1304 0 -1 3970
box -8 -3 16 105
use FILL  FILL_240
timestamp 1745462530
transform 1 0 1200 0 -1 3970
box -8 -3 16 105
use FILL  FILL_241
timestamp 1745462530
transform 1 0 1192 0 -1 3970
box -8 -3 16 105
use FILL  FILL_242
timestamp 1745462530
transform 1 0 1088 0 -1 3970
box -8 -3 16 105
use FILL  FILL_243
timestamp 1745462530
transform 1 0 1080 0 -1 3970
box -8 -3 16 105
use FILL  FILL_244
timestamp 1745462530
transform 1 0 1032 0 -1 3970
box -8 -3 16 105
use FILL  FILL_245
timestamp 1745462530
transform 1 0 1024 0 -1 3970
box -8 -3 16 105
use FILL  FILL_246
timestamp 1745462530
transform 1 0 920 0 -1 3970
box -8 -3 16 105
use FILL  FILL_247
timestamp 1745462530
transform 1 0 912 0 -1 3970
box -8 -3 16 105
use FILL  FILL_248
timestamp 1745462530
transform 1 0 904 0 -1 3970
box -8 -3 16 105
use FILL  FILL_249
timestamp 1745462530
transform 1 0 800 0 -1 3970
box -8 -3 16 105
use FILL  FILL_250
timestamp 1745462530
transform 1 0 792 0 -1 3970
box -8 -3 16 105
use FILL  FILL_251
timestamp 1745462530
transform 1 0 736 0 -1 3970
box -8 -3 16 105
use FILL  FILL_252
timestamp 1745462530
transform 1 0 728 0 -1 3970
box -8 -3 16 105
use FILL  FILL_253
timestamp 1745462530
transform 1 0 624 0 -1 3970
box -8 -3 16 105
use FILL  FILL_254
timestamp 1745462530
transform 1 0 616 0 -1 3970
box -8 -3 16 105
use FILL  FILL_255
timestamp 1745462530
transform 1 0 576 0 -1 3970
box -8 -3 16 105
use FILL  FILL_256
timestamp 1745462530
transform 1 0 568 0 -1 3970
box -8 -3 16 105
use FILL  FILL_257
timestamp 1745462530
transform 1 0 536 0 -1 3970
box -8 -3 16 105
use FILL  FILL_258
timestamp 1745462530
transform 1 0 496 0 -1 3970
box -8 -3 16 105
use FILL  FILL_259
timestamp 1745462530
transform 1 0 488 0 -1 3970
box -8 -3 16 105
use FILL  FILL_260
timestamp 1745462530
transform 1 0 456 0 -1 3970
box -8 -3 16 105
use FILL  FILL_261
timestamp 1745462530
transform 1 0 448 0 -1 3970
box -8 -3 16 105
use FILL  FILL_262
timestamp 1745462530
transform 1 0 440 0 -1 3970
box -8 -3 16 105
use FILL  FILL_263
timestamp 1745462530
transform 1 0 432 0 -1 3970
box -8 -3 16 105
use FILL  FILL_264
timestamp 1745462530
transform 1 0 328 0 -1 3970
box -8 -3 16 105
use FILL  FILL_265
timestamp 1745462530
transform 1 0 320 0 -1 3970
box -8 -3 16 105
use FILL  FILL_266
timestamp 1745462530
transform 1 0 296 0 -1 3970
box -8 -3 16 105
use FILL  FILL_267
timestamp 1745462530
transform 1 0 288 0 -1 3970
box -8 -3 16 105
use FILL  FILL_268
timestamp 1745462530
transform 1 0 184 0 -1 3970
box -8 -3 16 105
use FILL  FILL_269
timestamp 1745462530
transform 1 0 176 0 -1 3970
box -8 -3 16 105
use FILL  FILL_270
timestamp 1745462530
transform 1 0 144 0 -1 3970
box -8 -3 16 105
use FILL  FILL_271
timestamp 1745462530
transform 1 0 136 0 -1 3970
box -8 -3 16 105
use FILL  FILL_272
timestamp 1745462530
transform 1 0 112 0 -1 3970
box -8 -3 16 105
use FILL  FILL_273
timestamp 1745462530
transform 1 0 72 0 -1 3970
box -8 -3 16 105
use FILL  FILL_274
timestamp 1745462530
transform 1 0 4272 0 1 3770
box -8 -3 16 105
use FILL  FILL_275
timestamp 1745462530
transform 1 0 4264 0 1 3770
box -8 -3 16 105
use FILL  FILL_276
timestamp 1745462530
transform 1 0 4144 0 1 3770
box -8 -3 16 105
use FILL  FILL_277
timestamp 1745462530
transform 1 0 4136 0 1 3770
box -8 -3 16 105
use FILL  FILL_278
timestamp 1745462530
transform 1 0 4064 0 1 3770
box -8 -3 16 105
use FILL  FILL_279
timestamp 1745462530
transform 1 0 4016 0 1 3770
box -8 -3 16 105
use FILL  FILL_280
timestamp 1745462530
transform 1 0 4008 0 1 3770
box -8 -3 16 105
use FILL  FILL_281
timestamp 1745462530
transform 1 0 3960 0 1 3770
box -8 -3 16 105
use FILL  FILL_282
timestamp 1745462530
transform 1 0 3928 0 1 3770
box -8 -3 16 105
use FILL  FILL_283
timestamp 1745462530
transform 1 0 3920 0 1 3770
box -8 -3 16 105
use FILL  FILL_284
timestamp 1745462530
transform 1 0 3816 0 1 3770
box -8 -3 16 105
use FILL  FILL_285
timestamp 1745462530
transform 1 0 3808 0 1 3770
box -8 -3 16 105
use FILL  FILL_286
timestamp 1745462530
transform 1 0 3704 0 1 3770
box -8 -3 16 105
use FILL  FILL_287
timestamp 1745462530
transform 1 0 3664 0 1 3770
box -8 -3 16 105
use FILL  FILL_288
timestamp 1745462530
transform 1 0 3600 0 1 3770
box -8 -3 16 105
use FILL  FILL_289
timestamp 1745462530
transform 1 0 3560 0 1 3770
box -8 -3 16 105
use FILL  FILL_290
timestamp 1745462530
transform 1 0 3512 0 1 3770
box -8 -3 16 105
use FILL  FILL_291
timestamp 1745462530
transform 1 0 3464 0 1 3770
box -8 -3 16 105
use FILL  FILL_292
timestamp 1745462530
transform 1 0 3408 0 1 3770
box -8 -3 16 105
use FILL  FILL_293
timestamp 1745462530
transform 1 0 3400 0 1 3770
box -8 -3 16 105
use FILL  FILL_294
timestamp 1745462530
transform 1 0 3336 0 1 3770
box -8 -3 16 105
use FILL  FILL_295
timestamp 1745462530
transform 1 0 3232 0 1 3770
box -8 -3 16 105
use FILL  FILL_296
timestamp 1745462530
transform 1 0 3176 0 1 3770
box -8 -3 16 105
use FILL  FILL_297
timestamp 1745462530
transform 1 0 3168 0 1 3770
box -8 -3 16 105
use FILL  FILL_298
timestamp 1745462530
transform 1 0 3104 0 1 3770
box -8 -3 16 105
use FILL  FILL_299
timestamp 1745462530
transform 1 0 3000 0 1 3770
box -8 -3 16 105
use FILL  FILL_300
timestamp 1745462530
transform 1 0 2896 0 1 3770
box -8 -3 16 105
use FILL  FILL_301
timestamp 1745462530
transform 1 0 2872 0 1 3770
box -8 -3 16 105
use FILL  FILL_302
timestamp 1745462530
transform 1 0 2768 0 1 3770
box -8 -3 16 105
use FILL  FILL_303
timestamp 1745462530
transform 1 0 2696 0 1 3770
box -8 -3 16 105
use FILL  FILL_304
timestamp 1745462530
transform 1 0 2656 0 1 3770
box -8 -3 16 105
use FILL  FILL_305
timestamp 1745462530
transform 1 0 2608 0 1 3770
box -8 -3 16 105
use FILL  FILL_306
timestamp 1745462530
transform 1 0 2576 0 1 3770
box -8 -3 16 105
use FILL  FILL_307
timestamp 1745462530
transform 1 0 2528 0 1 3770
box -8 -3 16 105
use FILL  FILL_308
timestamp 1745462530
transform 1 0 2464 0 1 3770
box -8 -3 16 105
use FILL  FILL_309
timestamp 1745462530
transform 1 0 2456 0 1 3770
box -8 -3 16 105
use FILL  FILL_310
timestamp 1745462530
transform 1 0 2424 0 1 3770
box -8 -3 16 105
use FILL  FILL_311
timestamp 1745462530
transform 1 0 2392 0 1 3770
box -8 -3 16 105
use FILL  FILL_312
timestamp 1745462530
transform 1 0 2384 0 1 3770
box -8 -3 16 105
use FILL  FILL_313
timestamp 1745462530
transform 1 0 2344 0 1 3770
box -8 -3 16 105
use FILL  FILL_314
timestamp 1745462530
transform 1 0 2304 0 1 3770
box -8 -3 16 105
use FILL  FILL_315
timestamp 1745462530
transform 1 0 2296 0 1 3770
box -8 -3 16 105
use FILL  FILL_316
timestamp 1745462530
transform 1 0 2232 0 1 3770
box -8 -3 16 105
use FILL  FILL_317
timestamp 1745462530
transform 1 0 2224 0 1 3770
box -8 -3 16 105
use FILL  FILL_318
timestamp 1745462530
transform 1 0 2184 0 1 3770
box -8 -3 16 105
use FILL  FILL_319
timestamp 1745462530
transform 1 0 2160 0 1 3770
box -8 -3 16 105
use FILL  FILL_320
timestamp 1745462530
transform 1 0 2128 0 1 3770
box -8 -3 16 105
use FILL  FILL_321
timestamp 1745462530
transform 1 0 2088 0 1 3770
box -8 -3 16 105
use FILL  FILL_322
timestamp 1745462530
transform 1 0 2056 0 1 3770
box -8 -3 16 105
use FILL  FILL_323
timestamp 1745462530
transform 1 0 1992 0 1 3770
box -8 -3 16 105
use FILL  FILL_324
timestamp 1745462530
transform 1 0 1888 0 1 3770
box -8 -3 16 105
use FILL  FILL_325
timestamp 1745462530
transform 1 0 1880 0 1 3770
box -8 -3 16 105
use FILL  FILL_326
timestamp 1745462530
transform 1 0 1816 0 1 3770
box -8 -3 16 105
use FILL  FILL_327
timestamp 1745462530
transform 1 0 1768 0 1 3770
box -8 -3 16 105
use FILL  FILL_328
timestamp 1745462530
transform 1 0 1760 0 1 3770
box -8 -3 16 105
use FILL  FILL_329
timestamp 1745462530
transform 1 0 1712 0 1 3770
box -8 -3 16 105
use FILL  FILL_330
timestamp 1745462530
transform 1 0 1648 0 1 3770
box -8 -3 16 105
use FILL  FILL_331
timestamp 1745462530
transform 1 0 1640 0 1 3770
box -8 -3 16 105
use FILL  FILL_332
timestamp 1745462530
transform 1 0 1576 0 1 3770
box -8 -3 16 105
use FILL  FILL_333
timestamp 1745462530
transform 1 0 1552 0 1 3770
box -8 -3 16 105
use FILL  FILL_334
timestamp 1745462530
transform 1 0 1544 0 1 3770
box -8 -3 16 105
use FILL  FILL_335
timestamp 1745462530
transform 1 0 1440 0 1 3770
box -8 -3 16 105
use FILL  FILL_336
timestamp 1745462530
transform 1 0 1432 0 1 3770
box -8 -3 16 105
use FILL  FILL_337
timestamp 1745462530
transform 1 0 1328 0 1 3770
box -8 -3 16 105
use FILL  FILL_338
timestamp 1745462530
transform 1 0 1320 0 1 3770
box -8 -3 16 105
use FILL  FILL_339
timestamp 1745462530
transform 1 0 1264 0 1 3770
box -8 -3 16 105
use FILL  FILL_340
timestamp 1745462530
transform 1 0 1256 0 1 3770
box -8 -3 16 105
use FILL  FILL_341
timestamp 1745462530
transform 1 0 1248 0 1 3770
box -8 -3 16 105
use FILL  FILL_342
timestamp 1745462530
transform 1 0 1200 0 1 3770
box -8 -3 16 105
use FILL  FILL_343
timestamp 1745462530
transform 1 0 1168 0 1 3770
box -8 -3 16 105
use FILL  FILL_344
timestamp 1745462530
transform 1 0 1160 0 1 3770
box -8 -3 16 105
use FILL  FILL_345
timestamp 1745462530
transform 1 0 1096 0 1 3770
box -8 -3 16 105
use FILL  FILL_346
timestamp 1745462530
transform 1 0 1088 0 1 3770
box -8 -3 16 105
use FILL  FILL_347
timestamp 1745462530
transform 1 0 1080 0 1 3770
box -8 -3 16 105
use FILL  FILL_348
timestamp 1745462530
transform 1 0 976 0 1 3770
box -8 -3 16 105
use FILL  FILL_349
timestamp 1745462530
transform 1 0 968 0 1 3770
box -8 -3 16 105
use FILL  FILL_350
timestamp 1745462530
transform 1 0 960 0 1 3770
box -8 -3 16 105
use FILL  FILL_351
timestamp 1745462530
transform 1 0 952 0 1 3770
box -8 -3 16 105
use FILL  FILL_352
timestamp 1745462530
transform 1 0 848 0 1 3770
box -8 -3 16 105
use FILL  FILL_353
timestamp 1745462530
transform 1 0 840 0 1 3770
box -8 -3 16 105
use FILL  FILL_354
timestamp 1745462530
transform 1 0 832 0 1 3770
box -8 -3 16 105
use FILL  FILL_355
timestamp 1745462530
transform 1 0 824 0 1 3770
box -8 -3 16 105
use FILL  FILL_356
timestamp 1745462530
transform 1 0 816 0 1 3770
box -8 -3 16 105
use FILL  FILL_357
timestamp 1745462530
transform 1 0 808 0 1 3770
box -8 -3 16 105
use FILL  FILL_358
timestamp 1745462530
transform 1 0 752 0 1 3770
box -8 -3 16 105
use FILL  FILL_359
timestamp 1745462530
transform 1 0 744 0 1 3770
box -8 -3 16 105
use FILL  FILL_360
timestamp 1745462530
transform 1 0 736 0 1 3770
box -8 -3 16 105
use FILL  FILL_361
timestamp 1745462530
transform 1 0 632 0 1 3770
box -8 -3 16 105
use FILL  FILL_362
timestamp 1745462530
transform 1 0 624 0 1 3770
box -8 -3 16 105
use FILL  FILL_363
timestamp 1745462530
transform 1 0 616 0 1 3770
box -8 -3 16 105
use FILL  FILL_364
timestamp 1745462530
transform 1 0 608 0 1 3770
box -8 -3 16 105
use FILL  FILL_365
timestamp 1745462530
transform 1 0 504 0 1 3770
box -8 -3 16 105
use FILL  FILL_366
timestamp 1745462530
transform 1 0 496 0 1 3770
box -8 -3 16 105
use FILL  FILL_367
timestamp 1745462530
transform 1 0 472 0 1 3770
box -8 -3 16 105
use FILL  FILL_368
timestamp 1745462530
transform 1 0 464 0 1 3770
box -8 -3 16 105
use FILL  FILL_369
timestamp 1745462530
transform 1 0 360 0 1 3770
box -8 -3 16 105
use FILL  FILL_370
timestamp 1745462530
transform 1 0 352 0 1 3770
box -8 -3 16 105
use FILL  FILL_371
timestamp 1745462530
transform 1 0 344 0 1 3770
box -8 -3 16 105
use FILL  FILL_372
timestamp 1745462530
transform 1 0 240 0 1 3770
box -8 -3 16 105
use FILL  FILL_373
timestamp 1745462530
transform 1 0 232 0 1 3770
box -8 -3 16 105
use FILL  FILL_374
timestamp 1745462530
transform 1 0 224 0 1 3770
box -8 -3 16 105
use FILL  FILL_375
timestamp 1745462530
transform 1 0 184 0 1 3770
box -8 -3 16 105
use FILL  FILL_376
timestamp 1745462530
transform 1 0 144 0 1 3770
box -8 -3 16 105
use FILL  FILL_377
timestamp 1745462530
transform 1 0 136 0 1 3770
box -8 -3 16 105
use FILL  FILL_378
timestamp 1745462530
transform 1 0 96 0 1 3770
box -8 -3 16 105
use FILL  FILL_379
timestamp 1745462530
transform 1 0 72 0 1 3770
box -8 -3 16 105
use FILL  FILL_380
timestamp 1745462530
transform 1 0 4352 0 -1 3770
box -8 -3 16 105
use FILL  FILL_381
timestamp 1745462530
transform 1 0 4344 0 -1 3770
box -8 -3 16 105
use FILL  FILL_382
timestamp 1745462530
transform 1 0 4336 0 -1 3770
box -8 -3 16 105
use FILL  FILL_383
timestamp 1745462530
transform 1 0 4272 0 -1 3770
box -8 -3 16 105
use FILL  FILL_384
timestamp 1745462530
transform 1 0 4264 0 -1 3770
box -8 -3 16 105
use FILL  FILL_385
timestamp 1745462530
transform 1 0 4216 0 -1 3770
box -8 -3 16 105
use FILL  FILL_386
timestamp 1745462530
transform 1 0 4184 0 -1 3770
box -8 -3 16 105
use FILL  FILL_387
timestamp 1745462530
transform 1 0 4136 0 -1 3770
box -8 -3 16 105
use FILL  FILL_388
timestamp 1745462530
transform 1 0 4088 0 -1 3770
box -8 -3 16 105
use FILL  FILL_389
timestamp 1745462530
transform 1 0 4080 0 -1 3770
box -8 -3 16 105
use FILL  FILL_390
timestamp 1745462530
transform 1 0 4032 0 -1 3770
box -8 -3 16 105
use FILL  FILL_391
timestamp 1745462530
transform 1 0 4000 0 -1 3770
box -8 -3 16 105
use FILL  FILL_392
timestamp 1745462530
transform 1 0 3992 0 -1 3770
box -8 -3 16 105
use FILL  FILL_393
timestamp 1745462530
transform 1 0 3888 0 -1 3770
box -8 -3 16 105
use FILL  FILL_394
timestamp 1745462530
transform 1 0 3864 0 -1 3770
box -8 -3 16 105
use FILL  FILL_395
timestamp 1745462530
transform 1 0 3856 0 -1 3770
box -8 -3 16 105
use FILL  FILL_396
timestamp 1745462530
transform 1 0 3792 0 -1 3770
box -8 -3 16 105
use FILL  FILL_397
timestamp 1745462530
transform 1 0 3784 0 -1 3770
box -8 -3 16 105
use FILL  FILL_398
timestamp 1745462530
transform 1 0 3720 0 -1 3770
box -8 -3 16 105
use FILL  FILL_399
timestamp 1745462530
transform 1 0 3712 0 -1 3770
box -8 -3 16 105
use FILL  FILL_400
timestamp 1745462530
transform 1 0 3648 0 -1 3770
box -8 -3 16 105
use FILL  FILL_401
timestamp 1745462530
transform 1 0 3640 0 -1 3770
box -8 -3 16 105
use FILL  FILL_402
timestamp 1745462530
transform 1 0 3544 0 -1 3770
box -8 -3 16 105
use FILL  FILL_403
timestamp 1745462530
transform 1 0 3496 0 -1 3770
box -8 -3 16 105
use FILL  FILL_404
timestamp 1745462530
transform 1 0 3448 0 -1 3770
box -8 -3 16 105
use FILL  FILL_405
timestamp 1745462530
transform 1 0 3440 0 -1 3770
box -8 -3 16 105
use FILL  FILL_406
timestamp 1745462530
transform 1 0 3376 0 -1 3770
box -8 -3 16 105
use FILL  FILL_407
timestamp 1745462530
transform 1 0 3312 0 -1 3770
box -8 -3 16 105
use FILL  FILL_408
timestamp 1745462530
transform 1 0 3256 0 -1 3770
box -8 -3 16 105
use FILL  FILL_409
timestamp 1745462530
transform 1 0 3184 0 -1 3770
box -8 -3 16 105
use FILL  FILL_410
timestamp 1745462530
transform 1 0 3112 0 -1 3770
box -8 -3 16 105
use FILL  FILL_411
timestamp 1745462530
transform 1 0 3048 0 -1 3770
box -8 -3 16 105
use FILL  FILL_412
timestamp 1745462530
transform 1 0 3040 0 -1 3770
box -8 -3 16 105
use FILL  FILL_413
timestamp 1745462530
transform 1 0 2976 0 -1 3770
box -8 -3 16 105
use FILL  FILL_414
timestamp 1745462530
transform 1 0 2912 0 -1 3770
box -8 -3 16 105
use FILL  FILL_415
timestamp 1745462530
transform 1 0 2904 0 -1 3770
box -8 -3 16 105
use FILL  FILL_416
timestamp 1745462530
transform 1 0 2840 0 -1 3770
box -8 -3 16 105
use FILL  FILL_417
timestamp 1745462530
transform 1 0 2832 0 -1 3770
box -8 -3 16 105
use FILL  FILL_418
timestamp 1745462530
transform 1 0 2768 0 -1 3770
box -8 -3 16 105
use FILL  FILL_419
timestamp 1745462530
transform 1 0 2728 0 -1 3770
box -8 -3 16 105
use FILL  FILL_420
timestamp 1745462530
transform 1 0 2696 0 -1 3770
box -8 -3 16 105
use FILL  FILL_421
timestamp 1745462530
transform 1 0 2688 0 -1 3770
box -8 -3 16 105
use FILL  FILL_422
timestamp 1745462530
transform 1 0 2648 0 -1 3770
box -8 -3 16 105
use FILL  FILL_423
timestamp 1745462530
transform 1 0 2608 0 -1 3770
box -8 -3 16 105
use FILL  FILL_424
timestamp 1745462530
transform 1 0 2568 0 -1 3770
box -8 -3 16 105
use FILL  FILL_425
timestamp 1745462530
transform 1 0 2528 0 -1 3770
box -8 -3 16 105
use FILL  FILL_426
timestamp 1745462530
transform 1 0 2496 0 -1 3770
box -8 -3 16 105
use FILL  FILL_427
timestamp 1745462530
transform 1 0 2488 0 -1 3770
box -8 -3 16 105
use FILL  FILL_428
timestamp 1745462530
transform 1 0 2448 0 -1 3770
box -8 -3 16 105
use FILL  FILL_429
timestamp 1745462530
transform 1 0 2440 0 -1 3770
box -8 -3 16 105
use FILL  FILL_430
timestamp 1745462530
transform 1 0 2400 0 -1 3770
box -8 -3 16 105
use FILL  FILL_431
timestamp 1745462530
transform 1 0 2392 0 -1 3770
box -8 -3 16 105
use FILL  FILL_432
timestamp 1745462530
transform 1 0 2384 0 -1 3770
box -8 -3 16 105
use FILL  FILL_433
timestamp 1745462530
transform 1 0 2344 0 -1 3770
box -8 -3 16 105
use FILL  FILL_434
timestamp 1745462530
transform 1 0 2312 0 -1 3770
box -8 -3 16 105
use FILL  FILL_435
timestamp 1745462530
transform 1 0 2304 0 -1 3770
box -8 -3 16 105
use FILL  FILL_436
timestamp 1745462530
transform 1 0 2264 0 -1 3770
box -8 -3 16 105
use FILL  FILL_437
timestamp 1745462530
transform 1 0 2256 0 -1 3770
box -8 -3 16 105
use FILL  FILL_438
timestamp 1745462530
transform 1 0 2248 0 -1 3770
box -8 -3 16 105
use FILL  FILL_439
timestamp 1745462530
transform 1 0 2208 0 -1 3770
box -8 -3 16 105
use FILL  FILL_440
timestamp 1745462530
transform 1 0 2176 0 -1 3770
box -8 -3 16 105
use FILL  FILL_441
timestamp 1745462530
transform 1 0 2168 0 -1 3770
box -8 -3 16 105
use FILL  FILL_442
timestamp 1745462530
transform 1 0 2112 0 -1 3770
box -8 -3 16 105
use FILL  FILL_443
timestamp 1745462530
transform 1 0 2040 0 -1 3770
box -8 -3 16 105
use FILL  FILL_444
timestamp 1745462530
transform 1 0 2016 0 -1 3770
box -8 -3 16 105
use FILL  FILL_445
timestamp 1745462530
transform 1 0 1952 0 -1 3770
box -8 -3 16 105
use FILL  FILL_446
timestamp 1745462530
transform 1 0 1944 0 -1 3770
box -8 -3 16 105
use FILL  FILL_447
timestamp 1745462530
transform 1 0 1872 0 -1 3770
box -8 -3 16 105
use FILL  FILL_448
timestamp 1745462530
transform 1 0 1864 0 -1 3770
box -8 -3 16 105
use FILL  FILL_449
timestamp 1745462530
transform 1 0 1856 0 -1 3770
box -8 -3 16 105
use FILL  FILL_450
timestamp 1745462530
transform 1 0 1808 0 -1 3770
box -8 -3 16 105
use FILL  FILL_451
timestamp 1745462530
transform 1 0 1760 0 -1 3770
box -8 -3 16 105
use FILL  FILL_452
timestamp 1745462530
transform 1 0 1752 0 -1 3770
box -8 -3 16 105
use FILL  FILL_453
timestamp 1745462530
transform 1 0 1688 0 -1 3770
box -8 -3 16 105
use FILL  FILL_454
timestamp 1745462530
transform 1 0 1648 0 -1 3770
box -8 -3 16 105
use FILL  FILL_455
timestamp 1745462530
transform 1 0 1616 0 -1 3770
box -8 -3 16 105
use FILL  FILL_456
timestamp 1745462530
transform 1 0 1608 0 -1 3770
box -8 -3 16 105
use FILL  FILL_457
timestamp 1745462530
transform 1 0 1544 0 -1 3770
box -8 -3 16 105
use FILL  FILL_458
timestamp 1745462530
transform 1 0 1536 0 -1 3770
box -8 -3 16 105
use FILL  FILL_459
timestamp 1745462530
transform 1 0 1512 0 -1 3770
box -8 -3 16 105
use FILL  FILL_460
timestamp 1745462530
transform 1 0 1464 0 -1 3770
box -8 -3 16 105
use FILL  FILL_461
timestamp 1745462530
transform 1 0 1456 0 -1 3770
box -8 -3 16 105
use FILL  FILL_462
timestamp 1745462530
transform 1 0 1384 0 -1 3770
box -8 -3 16 105
use FILL  FILL_463
timestamp 1745462530
transform 1 0 1376 0 -1 3770
box -8 -3 16 105
use FILL  FILL_464
timestamp 1745462530
transform 1 0 1320 0 -1 3770
box -8 -3 16 105
use FILL  FILL_465
timestamp 1745462530
transform 1 0 1312 0 -1 3770
box -8 -3 16 105
use FILL  FILL_466
timestamp 1745462530
transform 1 0 1304 0 -1 3770
box -8 -3 16 105
use FILL  FILL_467
timestamp 1745462530
transform 1 0 1248 0 -1 3770
box -8 -3 16 105
use FILL  FILL_468
timestamp 1745462530
transform 1 0 1144 0 -1 3770
box -8 -3 16 105
use FILL  FILL_469
timestamp 1745462530
transform 1 0 1120 0 -1 3770
box -8 -3 16 105
use FILL  FILL_470
timestamp 1745462530
transform 1 0 1016 0 -1 3770
box -8 -3 16 105
use FILL  FILL_471
timestamp 1745462530
transform 1 0 1008 0 -1 3770
box -8 -3 16 105
use FILL  FILL_472
timestamp 1745462530
transform 1 0 1000 0 -1 3770
box -8 -3 16 105
use FILL  FILL_473
timestamp 1745462530
transform 1 0 944 0 -1 3770
box -8 -3 16 105
use FILL  FILL_474
timestamp 1745462530
transform 1 0 936 0 -1 3770
box -8 -3 16 105
use FILL  FILL_475
timestamp 1745462530
transform 1 0 832 0 -1 3770
box -8 -3 16 105
use FILL  FILL_476
timestamp 1745462530
transform 1 0 824 0 -1 3770
box -8 -3 16 105
use FILL  FILL_477
timestamp 1745462530
transform 1 0 720 0 -1 3770
box -8 -3 16 105
use FILL  FILL_478
timestamp 1745462530
transform 1 0 712 0 -1 3770
box -8 -3 16 105
use FILL  FILL_479
timestamp 1745462530
transform 1 0 656 0 -1 3770
box -8 -3 16 105
use FILL  FILL_480
timestamp 1745462530
transform 1 0 648 0 -1 3770
box -8 -3 16 105
use FILL  FILL_481
timestamp 1745462530
transform 1 0 640 0 -1 3770
box -8 -3 16 105
use FILL  FILL_482
timestamp 1745462530
transform 1 0 536 0 -1 3770
box -8 -3 16 105
use FILL  FILL_483
timestamp 1745462530
transform 1 0 528 0 -1 3770
box -8 -3 16 105
use FILL  FILL_484
timestamp 1745462530
transform 1 0 520 0 -1 3770
box -8 -3 16 105
use FILL  FILL_485
timestamp 1745462530
transform 1 0 512 0 -1 3770
box -8 -3 16 105
use FILL  FILL_486
timestamp 1745462530
transform 1 0 408 0 -1 3770
box -8 -3 16 105
use FILL  FILL_487
timestamp 1745462530
transform 1 0 400 0 -1 3770
box -8 -3 16 105
use FILL  FILL_488
timestamp 1745462530
transform 1 0 392 0 -1 3770
box -8 -3 16 105
use FILL  FILL_489
timestamp 1745462530
transform 1 0 384 0 -1 3770
box -8 -3 16 105
use FILL  FILL_490
timestamp 1745462530
transform 1 0 376 0 -1 3770
box -8 -3 16 105
use FILL  FILL_491
timestamp 1745462530
transform 1 0 272 0 -1 3770
box -8 -3 16 105
use FILL  FILL_492
timestamp 1745462530
transform 1 0 264 0 -1 3770
box -8 -3 16 105
use FILL  FILL_493
timestamp 1745462530
transform 1 0 256 0 -1 3770
box -8 -3 16 105
use FILL  FILL_494
timestamp 1745462530
transform 1 0 248 0 -1 3770
box -8 -3 16 105
use FILL  FILL_495
timestamp 1745462530
transform 1 0 240 0 -1 3770
box -8 -3 16 105
use FILL  FILL_496
timestamp 1745462530
transform 1 0 136 0 -1 3770
box -8 -3 16 105
use FILL  FILL_497
timestamp 1745462530
transform 1 0 128 0 -1 3770
box -8 -3 16 105
use FILL  FILL_498
timestamp 1745462530
transform 1 0 120 0 -1 3770
box -8 -3 16 105
use FILL  FILL_499
timestamp 1745462530
transform 1 0 112 0 -1 3770
box -8 -3 16 105
use FILL  FILL_500
timestamp 1745462530
transform 1 0 104 0 -1 3770
box -8 -3 16 105
use FILL  FILL_501
timestamp 1745462530
transform 1 0 96 0 -1 3770
box -8 -3 16 105
use FILL  FILL_502
timestamp 1745462530
transform 1 0 88 0 -1 3770
box -8 -3 16 105
use FILL  FILL_503
timestamp 1745462530
transform 1 0 80 0 -1 3770
box -8 -3 16 105
use FILL  FILL_504
timestamp 1745462530
transform 1 0 72 0 -1 3770
box -8 -3 16 105
use FILL  FILL_505
timestamp 1745462530
transform 1 0 4200 0 1 3570
box -8 -3 16 105
use FILL  FILL_506
timestamp 1745462530
transform 1 0 4080 0 1 3570
box -8 -3 16 105
use FILL  FILL_507
timestamp 1745462530
transform 1 0 4016 0 1 3570
box -8 -3 16 105
use FILL  FILL_508
timestamp 1745462530
transform 1 0 3896 0 1 3570
box -8 -3 16 105
use FILL  FILL_509
timestamp 1745462530
transform 1 0 3840 0 1 3570
box -8 -3 16 105
use FILL  FILL_510
timestamp 1745462530
transform 1 0 3832 0 1 3570
box -8 -3 16 105
use FILL  FILL_511
timestamp 1745462530
transform 1 0 3760 0 1 3570
box -8 -3 16 105
use FILL  FILL_512
timestamp 1745462530
transform 1 0 3752 0 1 3570
box -8 -3 16 105
use FILL  FILL_513
timestamp 1745462530
transform 1 0 3688 0 1 3570
box -8 -3 16 105
use FILL  FILL_514
timestamp 1745462530
transform 1 0 3648 0 1 3570
box -8 -3 16 105
use FILL  FILL_515
timestamp 1745462530
transform 1 0 3544 0 1 3570
box -8 -3 16 105
use FILL  FILL_516
timestamp 1745462530
transform 1 0 3480 0 1 3570
box -8 -3 16 105
use FILL  FILL_517
timestamp 1745462530
transform 1 0 3384 0 1 3570
box -8 -3 16 105
use FILL  FILL_518
timestamp 1745462530
transform 1 0 3376 0 1 3570
box -8 -3 16 105
use FILL  FILL_519
timestamp 1745462530
transform 1 0 3240 0 1 3570
box -8 -3 16 105
use FILL  FILL_520
timestamp 1745462530
transform 1 0 3232 0 1 3570
box -8 -3 16 105
use FILL  FILL_521
timestamp 1745462530
transform 1 0 3112 0 1 3570
box -8 -3 16 105
use FILL  FILL_522
timestamp 1745462530
transform 1 0 3104 0 1 3570
box -8 -3 16 105
use FILL  FILL_523
timestamp 1745462530
transform 1 0 3040 0 1 3570
box -8 -3 16 105
use FILL  FILL_524
timestamp 1745462530
transform 1 0 3032 0 1 3570
box -8 -3 16 105
use FILL  FILL_525
timestamp 1745462530
transform 1 0 2960 0 1 3570
box -8 -3 16 105
use FILL  FILL_526
timestamp 1745462530
transform 1 0 2952 0 1 3570
box -8 -3 16 105
use FILL  FILL_527
timestamp 1745462530
transform 1 0 2888 0 1 3570
box -8 -3 16 105
use FILL  FILL_528
timestamp 1745462530
transform 1 0 2880 0 1 3570
box -8 -3 16 105
use FILL  FILL_529
timestamp 1745462530
transform 1 0 2816 0 1 3570
box -8 -3 16 105
use FILL  FILL_530
timestamp 1745462530
transform 1 0 2808 0 1 3570
box -8 -3 16 105
use FILL  FILL_531
timestamp 1745462530
transform 1 0 2800 0 1 3570
box -8 -3 16 105
use FILL  FILL_532
timestamp 1745462530
transform 1 0 2736 0 1 3570
box -8 -3 16 105
use FILL  FILL_533
timestamp 1745462530
transform 1 0 2696 0 1 3570
box -8 -3 16 105
use FILL  FILL_534
timestamp 1745462530
transform 1 0 2664 0 1 3570
box -8 -3 16 105
use FILL  FILL_535
timestamp 1745462530
transform 1 0 2624 0 1 3570
box -8 -3 16 105
use FILL  FILL_536
timestamp 1745462530
transform 1 0 2616 0 1 3570
box -8 -3 16 105
use FILL  FILL_537
timestamp 1745462530
transform 1 0 2576 0 1 3570
box -8 -3 16 105
use FILL  FILL_538
timestamp 1745462530
transform 1 0 2536 0 1 3570
box -8 -3 16 105
use FILL  FILL_539
timestamp 1745462530
transform 1 0 2496 0 1 3570
box -8 -3 16 105
use FILL  FILL_540
timestamp 1745462530
transform 1 0 2448 0 1 3570
box -8 -3 16 105
use FILL  FILL_541
timestamp 1745462530
transform 1 0 2440 0 1 3570
box -8 -3 16 105
use FILL  FILL_542
timestamp 1745462530
transform 1 0 2400 0 1 3570
box -8 -3 16 105
use FILL  FILL_543
timestamp 1745462530
transform 1 0 2368 0 1 3570
box -8 -3 16 105
use FILL  FILL_544
timestamp 1745462530
transform 1 0 2360 0 1 3570
box -8 -3 16 105
use FILL  FILL_545
timestamp 1745462530
transform 1 0 2320 0 1 3570
box -8 -3 16 105
use FILL  FILL_546
timestamp 1745462530
transform 1 0 2312 0 1 3570
box -8 -3 16 105
use FILL  FILL_547
timestamp 1745462530
transform 1 0 2280 0 1 3570
box -8 -3 16 105
use FILL  FILL_548
timestamp 1745462530
transform 1 0 2240 0 1 3570
box -8 -3 16 105
use FILL  FILL_549
timestamp 1745462530
transform 1 0 2232 0 1 3570
box -8 -3 16 105
use FILL  FILL_550
timestamp 1745462530
transform 1 0 2176 0 1 3570
box -8 -3 16 105
use FILL  FILL_551
timestamp 1745462530
transform 1 0 2168 0 1 3570
box -8 -3 16 105
use FILL  FILL_552
timestamp 1745462530
transform 1 0 2128 0 1 3570
box -8 -3 16 105
use FILL  FILL_553
timestamp 1745462530
transform 1 0 2120 0 1 3570
box -8 -3 16 105
use FILL  FILL_554
timestamp 1745462530
transform 1 0 2072 0 1 3570
box -8 -3 16 105
use FILL  FILL_555
timestamp 1745462530
transform 1 0 2064 0 1 3570
box -8 -3 16 105
use FILL  FILL_556
timestamp 1745462530
transform 1 0 2000 0 1 3570
box -8 -3 16 105
use FILL  FILL_557
timestamp 1745462530
transform 1 0 1896 0 1 3570
box -8 -3 16 105
use FILL  FILL_558
timestamp 1745462530
transform 1 0 1856 0 1 3570
box -8 -3 16 105
use FILL  FILL_559
timestamp 1745462530
transform 1 0 1848 0 1 3570
box -8 -3 16 105
use FILL  FILL_560
timestamp 1745462530
transform 1 0 1808 0 1 3570
box -8 -3 16 105
use FILL  FILL_561
timestamp 1745462530
transform 1 0 1800 0 1 3570
box -8 -3 16 105
use FILL  FILL_562
timestamp 1745462530
transform 1 0 1760 0 1 3570
box -8 -3 16 105
use FILL  FILL_563
timestamp 1745462530
transform 1 0 1720 0 1 3570
box -8 -3 16 105
use FILL  FILL_564
timestamp 1745462530
transform 1 0 1680 0 1 3570
box -8 -3 16 105
use FILL  FILL_565
timestamp 1745462530
transform 1 0 1648 0 1 3570
box -8 -3 16 105
use FILL  FILL_566
timestamp 1745462530
transform 1 0 1616 0 1 3570
box -8 -3 16 105
use FILL  FILL_567
timestamp 1745462530
transform 1 0 1576 0 1 3570
box -8 -3 16 105
use FILL  FILL_568
timestamp 1745462530
transform 1 0 1536 0 1 3570
box -8 -3 16 105
use FILL  FILL_569
timestamp 1745462530
transform 1 0 1488 0 1 3570
box -8 -3 16 105
use FILL  FILL_570
timestamp 1745462530
transform 1 0 1448 0 1 3570
box -8 -3 16 105
use FILL  FILL_571
timestamp 1745462530
transform 1 0 1408 0 1 3570
box -8 -3 16 105
use FILL  FILL_572
timestamp 1745462530
transform 1 0 1368 0 1 3570
box -8 -3 16 105
use FILL  FILL_573
timestamp 1745462530
transform 1 0 1360 0 1 3570
box -8 -3 16 105
use FILL  FILL_574
timestamp 1745462530
transform 1 0 1312 0 1 3570
box -8 -3 16 105
use FILL  FILL_575
timestamp 1745462530
transform 1 0 1264 0 1 3570
box -8 -3 16 105
use FILL  FILL_576
timestamp 1745462530
transform 1 0 1256 0 1 3570
box -8 -3 16 105
use FILL  FILL_577
timestamp 1745462530
transform 1 0 1152 0 1 3570
box -8 -3 16 105
use FILL  FILL_578
timestamp 1745462530
transform 1 0 1144 0 1 3570
box -8 -3 16 105
use FILL  FILL_579
timestamp 1745462530
transform 1 0 1064 0 1 3570
box -8 -3 16 105
use FILL  FILL_580
timestamp 1745462530
transform 1 0 1056 0 1 3570
box -8 -3 16 105
use FILL  FILL_581
timestamp 1745462530
transform 1 0 1048 0 1 3570
box -8 -3 16 105
use FILL  FILL_582
timestamp 1745462530
transform 1 0 1040 0 1 3570
box -8 -3 16 105
use FILL  FILL_583
timestamp 1745462530
transform 1 0 984 0 1 3570
box -8 -3 16 105
use FILL  FILL_584
timestamp 1745462530
transform 1 0 880 0 1 3570
box -8 -3 16 105
use FILL  FILL_585
timestamp 1745462530
transform 1 0 872 0 1 3570
box -8 -3 16 105
use FILL  FILL_586
timestamp 1745462530
transform 1 0 848 0 1 3570
box -8 -3 16 105
use FILL  FILL_587
timestamp 1745462530
transform 1 0 744 0 1 3570
box -8 -3 16 105
use FILL  FILL_588
timestamp 1745462530
transform 1 0 736 0 1 3570
box -8 -3 16 105
use FILL  FILL_589
timestamp 1745462530
transform 1 0 728 0 1 3570
box -8 -3 16 105
use FILL  FILL_590
timestamp 1745462530
transform 1 0 720 0 1 3570
box -8 -3 16 105
use FILL  FILL_591
timestamp 1745462530
transform 1 0 616 0 1 3570
box -8 -3 16 105
use FILL  FILL_592
timestamp 1745462530
transform 1 0 608 0 1 3570
box -8 -3 16 105
use FILL  FILL_593
timestamp 1745462530
transform 1 0 600 0 1 3570
box -8 -3 16 105
use FILL  FILL_594
timestamp 1745462530
transform 1 0 496 0 1 3570
box -8 -3 16 105
use FILL  FILL_595
timestamp 1745462530
transform 1 0 488 0 1 3570
box -8 -3 16 105
use FILL  FILL_596
timestamp 1745462530
transform 1 0 384 0 1 3570
box -8 -3 16 105
use FILL  FILL_597
timestamp 1745462530
transform 1 0 376 0 1 3570
box -8 -3 16 105
use FILL  FILL_598
timestamp 1745462530
transform 1 0 368 0 1 3570
box -8 -3 16 105
use FILL  FILL_599
timestamp 1745462530
transform 1 0 312 0 1 3570
box -8 -3 16 105
use FILL  FILL_600
timestamp 1745462530
transform 1 0 240 0 1 3570
box -8 -3 16 105
use FILL  FILL_601
timestamp 1745462530
transform 1 0 232 0 1 3570
box -8 -3 16 105
use FILL  FILL_602
timestamp 1745462530
transform 1 0 176 0 1 3570
box -8 -3 16 105
use FILL  FILL_603
timestamp 1745462530
transform 1 0 72 0 1 3570
box -8 -3 16 105
use FILL  FILL_604
timestamp 1745462530
transform 1 0 4368 0 -1 3570
box -8 -3 16 105
use FILL  FILL_605
timestamp 1745462530
transform 1 0 4264 0 -1 3570
box -8 -3 16 105
use FILL  FILL_606
timestamp 1745462530
transform 1 0 4256 0 -1 3570
box -8 -3 16 105
use FILL  FILL_607
timestamp 1745462530
transform 1 0 4248 0 -1 3570
box -8 -3 16 105
use FILL  FILL_608
timestamp 1745462530
transform 1 0 4144 0 -1 3570
box -8 -3 16 105
use FILL  FILL_609
timestamp 1745462530
transform 1 0 4104 0 -1 3570
box -8 -3 16 105
use FILL  FILL_610
timestamp 1745462530
transform 1 0 4056 0 -1 3570
box -8 -3 16 105
use FILL  FILL_611
timestamp 1745462530
transform 1 0 4048 0 -1 3570
box -8 -3 16 105
use FILL  FILL_612
timestamp 1745462530
transform 1 0 4040 0 -1 3570
box -8 -3 16 105
use FILL  FILL_613
timestamp 1745462530
transform 1 0 4016 0 -1 3570
box -8 -3 16 105
use FILL  FILL_614
timestamp 1745462530
transform 1 0 4008 0 -1 3570
box -8 -3 16 105
use FILL  FILL_615
timestamp 1745462530
transform 1 0 4000 0 -1 3570
box -8 -3 16 105
use FILL  FILL_616
timestamp 1745462530
transform 1 0 3992 0 -1 3570
box -8 -3 16 105
use FILL  FILL_617
timestamp 1745462530
transform 1 0 3928 0 -1 3570
box -8 -3 16 105
use FILL  FILL_618
timestamp 1745462530
transform 1 0 3920 0 -1 3570
box -8 -3 16 105
use FILL  FILL_619
timestamp 1745462530
transform 1 0 3912 0 -1 3570
box -8 -3 16 105
use FILL  FILL_620
timestamp 1745462530
transform 1 0 3848 0 -1 3570
box -8 -3 16 105
use FILL  FILL_621
timestamp 1745462530
transform 1 0 3840 0 -1 3570
box -8 -3 16 105
use FILL  FILL_622
timestamp 1745462530
transform 1 0 3776 0 -1 3570
box -8 -3 16 105
use FILL  FILL_623
timestamp 1745462530
transform 1 0 3768 0 -1 3570
box -8 -3 16 105
use FILL  FILL_624
timestamp 1745462530
transform 1 0 3704 0 -1 3570
box -8 -3 16 105
use FILL  FILL_625
timestamp 1745462530
transform 1 0 3664 0 -1 3570
box -8 -3 16 105
use FILL  FILL_626
timestamp 1745462530
transform 1 0 3624 0 -1 3570
box -8 -3 16 105
use FILL  FILL_627
timestamp 1745462530
transform 1 0 3584 0 -1 3570
box -8 -3 16 105
use FILL  FILL_628
timestamp 1745462530
transform 1 0 3536 0 -1 3570
box -8 -3 16 105
use FILL  FILL_629
timestamp 1745462530
transform 1 0 3448 0 -1 3570
box -8 -3 16 105
use FILL  FILL_630
timestamp 1745462530
transform 1 0 3368 0 -1 3570
box -8 -3 16 105
use FILL  FILL_631
timestamp 1745462530
transform 1 0 3248 0 -1 3570
box -8 -3 16 105
use FILL  FILL_632
timestamp 1745462530
transform 1 0 3168 0 -1 3570
box -8 -3 16 105
use FILL  FILL_633
timestamp 1745462530
transform 1 0 3088 0 -1 3570
box -8 -3 16 105
use FILL  FILL_634
timestamp 1745462530
transform 1 0 3040 0 -1 3570
box -8 -3 16 105
use FILL  FILL_635
timestamp 1745462530
transform 1 0 2920 0 -1 3570
box -8 -3 16 105
use FILL  FILL_636
timestamp 1745462530
transform 1 0 2912 0 -1 3570
box -8 -3 16 105
use FILL  FILL_637
timestamp 1745462530
transform 1 0 2864 0 -1 3570
box -8 -3 16 105
use FILL  FILL_638
timestamp 1745462530
transform 1 0 2824 0 -1 3570
box -8 -3 16 105
use FILL  FILL_639
timestamp 1745462530
transform 1 0 2776 0 -1 3570
box -8 -3 16 105
use FILL  FILL_640
timestamp 1745462530
transform 1 0 2736 0 -1 3570
box -8 -3 16 105
use FILL  FILL_641
timestamp 1745462530
transform 1 0 2728 0 -1 3570
box -8 -3 16 105
use FILL  FILL_642
timestamp 1745462530
transform 1 0 2680 0 -1 3570
box -8 -3 16 105
use FILL  FILL_643
timestamp 1745462530
transform 1 0 2640 0 -1 3570
box -8 -3 16 105
use FILL  FILL_644
timestamp 1745462530
transform 1 0 2592 0 -1 3570
box -8 -3 16 105
use FILL  FILL_645
timestamp 1745462530
transform 1 0 2584 0 -1 3570
box -8 -3 16 105
use FILL  FILL_646
timestamp 1745462530
transform 1 0 2536 0 -1 3570
box -8 -3 16 105
use FILL  FILL_647
timestamp 1745462530
transform 1 0 2528 0 -1 3570
box -8 -3 16 105
use FILL  FILL_648
timestamp 1745462530
transform 1 0 2480 0 -1 3570
box -8 -3 16 105
use FILL  FILL_649
timestamp 1745462530
transform 1 0 2472 0 -1 3570
box -8 -3 16 105
use FILL  FILL_650
timestamp 1745462530
transform 1 0 2424 0 -1 3570
box -8 -3 16 105
use FILL  FILL_651
timestamp 1745462530
transform 1 0 2376 0 -1 3570
box -8 -3 16 105
use FILL  FILL_652
timestamp 1745462530
transform 1 0 2368 0 -1 3570
box -8 -3 16 105
use FILL  FILL_653
timestamp 1745462530
transform 1 0 2360 0 -1 3570
box -8 -3 16 105
use FILL  FILL_654
timestamp 1745462530
transform 1 0 2320 0 -1 3570
box -8 -3 16 105
use FILL  FILL_655
timestamp 1745462530
transform 1 0 2280 0 -1 3570
box -8 -3 16 105
use FILL  FILL_656
timestamp 1745462530
transform 1 0 2272 0 -1 3570
box -8 -3 16 105
use FILL  FILL_657
timestamp 1745462530
transform 1 0 2264 0 -1 3570
box -8 -3 16 105
use FILL  FILL_658
timestamp 1745462530
transform 1 0 2224 0 -1 3570
box -8 -3 16 105
use FILL  FILL_659
timestamp 1745462530
transform 1 0 2216 0 -1 3570
box -8 -3 16 105
use FILL  FILL_660
timestamp 1745462530
transform 1 0 2168 0 -1 3570
box -8 -3 16 105
use FILL  FILL_661
timestamp 1745462530
transform 1 0 2160 0 -1 3570
box -8 -3 16 105
use FILL  FILL_662
timestamp 1745462530
transform 1 0 2152 0 -1 3570
box -8 -3 16 105
use FILL  FILL_663
timestamp 1745462530
transform 1 0 2112 0 -1 3570
box -8 -3 16 105
use FILL  FILL_664
timestamp 1745462530
transform 1 0 2104 0 -1 3570
box -8 -3 16 105
use FILL  FILL_665
timestamp 1745462530
transform 1 0 2072 0 -1 3570
box -8 -3 16 105
use FILL  FILL_666
timestamp 1745462530
transform 1 0 2040 0 -1 3570
box -8 -3 16 105
use FILL  FILL_667
timestamp 1745462530
transform 1 0 2032 0 -1 3570
box -8 -3 16 105
use FILL  FILL_668
timestamp 1745462530
transform 1 0 2024 0 -1 3570
box -8 -3 16 105
use FILL  FILL_669
timestamp 1745462530
transform 1 0 1984 0 -1 3570
box -8 -3 16 105
use FILL  FILL_670
timestamp 1745462530
transform 1 0 1976 0 -1 3570
box -8 -3 16 105
use FILL  FILL_671
timestamp 1745462530
transform 1 0 1944 0 -1 3570
box -8 -3 16 105
use FILL  FILL_672
timestamp 1745462530
transform 1 0 1936 0 -1 3570
box -8 -3 16 105
use FILL  FILL_673
timestamp 1745462530
transform 1 0 1896 0 -1 3570
box -8 -3 16 105
use FILL  FILL_674
timestamp 1745462530
transform 1 0 1888 0 -1 3570
box -8 -3 16 105
use FILL  FILL_675
timestamp 1745462530
transform 1 0 1880 0 -1 3570
box -8 -3 16 105
use FILL  FILL_676
timestamp 1745462530
transform 1 0 1840 0 -1 3570
box -8 -3 16 105
use FILL  FILL_677
timestamp 1745462530
transform 1 0 1808 0 -1 3570
box -8 -3 16 105
use FILL  FILL_678
timestamp 1745462530
transform 1 0 1800 0 -1 3570
box -8 -3 16 105
use FILL  FILL_679
timestamp 1745462530
transform 1 0 1736 0 -1 3570
box -8 -3 16 105
use FILL  FILL_680
timestamp 1745462530
transform 1 0 1728 0 -1 3570
box -8 -3 16 105
use FILL  FILL_681
timestamp 1745462530
transform 1 0 1664 0 -1 3570
box -8 -3 16 105
use FILL  FILL_682
timestamp 1745462530
transform 1 0 1656 0 -1 3570
box -8 -3 16 105
use FILL  FILL_683
timestamp 1745462530
transform 1 0 1648 0 -1 3570
box -8 -3 16 105
use FILL  FILL_684
timestamp 1745462530
transform 1 0 1592 0 -1 3570
box -8 -3 16 105
use FILL  FILL_685
timestamp 1745462530
transform 1 0 1560 0 -1 3570
box -8 -3 16 105
use FILL  FILL_686
timestamp 1745462530
transform 1 0 1512 0 -1 3570
box -8 -3 16 105
use FILL  FILL_687
timestamp 1745462530
transform 1 0 1488 0 -1 3570
box -8 -3 16 105
use FILL  FILL_688
timestamp 1745462530
transform 1 0 1440 0 -1 3570
box -8 -3 16 105
use FILL  FILL_689
timestamp 1745462530
transform 1 0 1432 0 -1 3570
box -8 -3 16 105
use FILL  FILL_690
timestamp 1745462530
transform 1 0 1360 0 -1 3570
box -8 -3 16 105
use FILL  FILL_691
timestamp 1745462530
transform 1 0 1256 0 -1 3570
box -8 -3 16 105
use FILL  FILL_692
timestamp 1745462530
transform 1 0 1248 0 -1 3570
box -8 -3 16 105
use FILL  FILL_693
timestamp 1745462530
transform 1 0 1184 0 -1 3570
box -8 -3 16 105
use FILL  FILL_694
timestamp 1745462530
transform 1 0 1176 0 -1 3570
box -8 -3 16 105
use FILL  FILL_695
timestamp 1745462530
transform 1 0 1112 0 -1 3570
box -8 -3 16 105
use FILL  FILL_696
timestamp 1745462530
transform 1 0 1080 0 -1 3570
box -8 -3 16 105
use FILL  FILL_697
timestamp 1745462530
transform 1 0 1024 0 -1 3570
box -8 -3 16 105
use FILL  FILL_698
timestamp 1745462530
transform 1 0 960 0 -1 3570
box -8 -3 16 105
use FILL  FILL_699
timestamp 1745462530
transform 1 0 920 0 -1 3570
box -8 -3 16 105
use FILL  FILL_700
timestamp 1745462530
transform 1 0 880 0 -1 3570
box -8 -3 16 105
use FILL  FILL_701
timestamp 1745462530
transform 1 0 840 0 -1 3570
box -8 -3 16 105
use FILL  FILL_702
timestamp 1745462530
transform 1 0 784 0 -1 3570
box -8 -3 16 105
use FILL  FILL_703
timestamp 1745462530
transform 1 0 776 0 -1 3570
box -8 -3 16 105
use FILL  FILL_704
timestamp 1745462530
transform 1 0 672 0 -1 3570
box -8 -3 16 105
use FILL  FILL_705
timestamp 1745462530
transform 1 0 664 0 -1 3570
box -8 -3 16 105
use FILL  FILL_706
timestamp 1745462530
transform 1 0 560 0 -1 3570
box -8 -3 16 105
use FILL  FILL_707
timestamp 1745462530
transform 1 0 552 0 -1 3570
box -8 -3 16 105
use FILL  FILL_708
timestamp 1745462530
transform 1 0 544 0 -1 3570
box -8 -3 16 105
use FILL  FILL_709
timestamp 1745462530
transform 1 0 440 0 -1 3570
box -8 -3 16 105
use FILL  FILL_710
timestamp 1745462530
transform 1 0 432 0 -1 3570
box -8 -3 16 105
use FILL  FILL_711
timestamp 1745462530
transform 1 0 376 0 -1 3570
box -8 -3 16 105
use FILL  FILL_712
timestamp 1745462530
transform 1 0 312 0 -1 3570
box -8 -3 16 105
use FILL  FILL_713
timestamp 1745462530
transform 1 0 304 0 -1 3570
box -8 -3 16 105
use FILL  FILL_714
timestamp 1745462530
transform 1 0 256 0 -1 3570
box -8 -3 16 105
use FILL  FILL_715
timestamp 1745462530
transform 1 0 216 0 -1 3570
box -8 -3 16 105
use FILL  FILL_716
timestamp 1745462530
transform 1 0 208 0 -1 3570
box -8 -3 16 105
use FILL  FILL_717
timestamp 1745462530
transform 1 0 152 0 -1 3570
box -8 -3 16 105
use FILL  FILL_718
timestamp 1745462530
transform 1 0 144 0 -1 3570
box -8 -3 16 105
use FILL  FILL_719
timestamp 1745462530
transform 1 0 96 0 -1 3570
box -8 -3 16 105
use FILL  FILL_720
timestamp 1745462530
transform 1 0 72 0 -1 3570
box -8 -3 16 105
use FILL  FILL_721
timestamp 1745462530
transform 1 0 4272 0 1 3370
box -8 -3 16 105
use FILL  FILL_722
timestamp 1745462530
transform 1 0 4248 0 1 3370
box -8 -3 16 105
use FILL  FILL_723
timestamp 1745462530
transform 1 0 4184 0 1 3370
box -8 -3 16 105
use FILL  FILL_724
timestamp 1745462530
transform 1 0 4024 0 1 3370
box -8 -3 16 105
use FILL  FILL_725
timestamp 1745462530
transform 1 0 4016 0 1 3370
box -8 -3 16 105
use FILL  FILL_726
timestamp 1745462530
transform 1 0 3888 0 1 3370
box -8 -3 16 105
use FILL  FILL_727
timestamp 1745462530
transform 1 0 3880 0 1 3370
box -8 -3 16 105
use FILL  FILL_728
timestamp 1745462530
transform 1 0 3872 0 1 3370
box -8 -3 16 105
use FILL  FILL_729
timestamp 1745462530
transform 1 0 3800 0 1 3370
box -8 -3 16 105
use FILL  FILL_730
timestamp 1745462530
transform 1 0 3792 0 1 3370
box -8 -3 16 105
use FILL  FILL_731
timestamp 1745462530
transform 1 0 3728 0 1 3370
box -8 -3 16 105
use FILL  FILL_732
timestamp 1745462530
transform 1 0 3656 0 1 3370
box -8 -3 16 105
use FILL  FILL_733
timestamp 1745462530
transform 1 0 3464 0 1 3370
box -8 -3 16 105
use FILL  FILL_734
timestamp 1745462530
transform 1 0 3344 0 1 3370
box -8 -3 16 105
use FILL  FILL_735
timestamp 1745462530
transform 1 0 3264 0 1 3370
box -8 -3 16 105
use FILL  FILL_736
timestamp 1745462530
transform 1 0 3184 0 1 3370
box -8 -3 16 105
use FILL  FILL_737
timestamp 1745462530
transform 1 0 3104 0 1 3370
box -8 -3 16 105
use FILL  FILL_738
timestamp 1745462530
transform 1 0 3024 0 1 3370
box -8 -3 16 105
use FILL  FILL_739
timestamp 1745462530
transform 1 0 2960 0 1 3370
box -8 -3 16 105
use FILL  FILL_740
timestamp 1745462530
transform 1 0 2880 0 1 3370
box -8 -3 16 105
use FILL  FILL_741
timestamp 1745462530
transform 1 0 2872 0 1 3370
box -8 -3 16 105
use FILL  FILL_742
timestamp 1745462530
transform 1 0 2808 0 1 3370
box -8 -3 16 105
use FILL  FILL_743
timestamp 1745462530
transform 1 0 2768 0 1 3370
box -8 -3 16 105
use FILL  FILL_744
timestamp 1745462530
transform 1 0 2760 0 1 3370
box -8 -3 16 105
use FILL  FILL_745
timestamp 1745462530
transform 1 0 2712 0 1 3370
box -8 -3 16 105
use FILL  FILL_746
timestamp 1745462530
transform 1 0 2672 0 1 3370
box -8 -3 16 105
use FILL  FILL_747
timestamp 1745462530
transform 1 0 2624 0 1 3370
box -8 -3 16 105
use FILL  FILL_748
timestamp 1745462530
transform 1 0 2576 0 1 3370
box -8 -3 16 105
use FILL  FILL_749
timestamp 1745462530
transform 1 0 2568 0 1 3370
box -8 -3 16 105
use FILL  FILL_750
timestamp 1745462530
transform 1 0 2520 0 1 3370
box -8 -3 16 105
use FILL  FILL_751
timestamp 1745462530
transform 1 0 2472 0 1 3370
box -8 -3 16 105
use FILL  FILL_752
timestamp 1745462530
transform 1 0 2464 0 1 3370
box -8 -3 16 105
use FILL  FILL_753
timestamp 1745462530
transform 1 0 2424 0 1 3370
box -8 -3 16 105
use FILL  FILL_754
timestamp 1745462530
transform 1 0 2384 0 1 3370
box -8 -3 16 105
use FILL  FILL_755
timestamp 1745462530
transform 1 0 2344 0 1 3370
box -8 -3 16 105
use FILL  FILL_756
timestamp 1745462530
transform 1 0 2304 0 1 3370
box -8 -3 16 105
use FILL  FILL_757
timestamp 1745462530
transform 1 0 2296 0 1 3370
box -8 -3 16 105
use FILL  FILL_758
timestamp 1745462530
transform 1 0 2256 0 1 3370
box -8 -3 16 105
use FILL  FILL_759
timestamp 1745462530
transform 1 0 2248 0 1 3370
box -8 -3 16 105
use FILL  FILL_760
timestamp 1745462530
transform 1 0 2208 0 1 3370
box -8 -3 16 105
use FILL  FILL_761
timestamp 1745462530
transform 1 0 2176 0 1 3370
box -8 -3 16 105
use FILL  FILL_762
timestamp 1745462530
transform 1 0 2136 0 1 3370
box -8 -3 16 105
use FILL  FILL_763
timestamp 1745462530
transform 1 0 2128 0 1 3370
box -8 -3 16 105
use FILL  FILL_764
timestamp 1745462530
transform 1 0 2120 0 1 3370
box -8 -3 16 105
use FILL  FILL_765
timestamp 1745462530
transform 1 0 2072 0 1 3370
box -8 -3 16 105
use FILL  FILL_766
timestamp 1745462530
transform 1 0 2064 0 1 3370
box -8 -3 16 105
use FILL  FILL_767
timestamp 1745462530
transform 1 0 2016 0 1 3370
box -8 -3 16 105
use FILL  FILL_768
timestamp 1745462530
transform 1 0 2008 0 1 3370
box -8 -3 16 105
use FILL  FILL_769
timestamp 1745462530
transform 1 0 1968 0 1 3370
box -8 -3 16 105
use FILL  FILL_770
timestamp 1745462530
transform 1 0 1960 0 1 3370
box -8 -3 16 105
use FILL  FILL_771
timestamp 1745462530
transform 1 0 1952 0 1 3370
box -8 -3 16 105
use FILL  FILL_772
timestamp 1745462530
transform 1 0 1920 0 1 3370
box -8 -3 16 105
use FILL  FILL_773
timestamp 1745462530
transform 1 0 1880 0 1 3370
box -8 -3 16 105
use FILL  FILL_774
timestamp 1745462530
transform 1 0 1872 0 1 3370
box -8 -3 16 105
use FILL  FILL_775
timestamp 1745462530
transform 1 0 1864 0 1 3370
box -8 -3 16 105
use FILL  FILL_776
timestamp 1745462530
transform 1 0 1824 0 1 3370
box -8 -3 16 105
use FILL  FILL_777
timestamp 1745462530
transform 1 0 1784 0 1 3370
box -8 -3 16 105
use FILL  FILL_778
timestamp 1745462530
transform 1 0 1760 0 1 3370
box -8 -3 16 105
use FILL  FILL_779
timestamp 1745462530
transform 1 0 1720 0 1 3370
box -8 -3 16 105
use FILL  FILL_780
timestamp 1745462530
transform 1 0 1688 0 1 3370
box -8 -3 16 105
use FILL  FILL_781
timestamp 1745462530
transform 1 0 1648 0 1 3370
box -8 -3 16 105
use FILL  FILL_782
timestamp 1745462530
transform 1 0 1608 0 1 3370
box -8 -3 16 105
use FILL  FILL_783
timestamp 1745462530
transform 1 0 1600 0 1 3370
box -8 -3 16 105
use FILL  FILL_784
timestamp 1745462530
transform 1 0 1536 0 1 3370
box -8 -3 16 105
use FILL  FILL_785
timestamp 1745462530
transform 1 0 1528 0 1 3370
box -8 -3 16 105
use FILL  FILL_786
timestamp 1745462530
transform 1 0 1464 0 1 3370
box -8 -3 16 105
use FILL  FILL_787
timestamp 1745462530
transform 1 0 1456 0 1 3370
box -8 -3 16 105
use FILL  FILL_788
timestamp 1745462530
transform 1 0 1416 0 1 3370
box -8 -3 16 105
use FILL  FILL_789
timestamp 1745462530
transform 1 0 1376 0 1 3370
box -8 -3 16 105
use FILL  FILL_790
timestamp 1745462530
transform 1 0 1272 0 1 3370
box -8 -3 16 105
use FILL  FILL_791
timestamp 1745462530
transform 1 0 1264 0 1 3370
box -8 -3 16 105
use FILL  FILL_792
timestamp 1745462530
transform 1 0 1160 0 1 3370
box -8 -3 16 105
use FILL  FILL_793
timestamp 1745462530
transform 1 0 1096 0 1 3370
box -8 -3 16 105
use FILL  FILL_794
timestamp 1745462530
transform 1 0 1088 0 1 3370
box -8 -3 16 105
use FILL  FILL_795
timestamp 1745462530
transform 1 0 992 0 1 3370
box -8 -3 16 105
use FILL  FILL_796
timestamp 1745462530
transform 1 0 984 0 1 3370
box -8 -3 16 105
use FILL  FILL_797
timestamp 1745462530
transform 1 0 912 0 1 3370
box -8 -3 16 105
use FILL  FILL_798
timestamp 1745462530
transform 1 0 872 0 1 3370
box -8 -3 16 105
use FILL  FILL_799
timestamp 1745462530
transform 1 0 864 0 1 3370
box -8 -3 16 105
use FILL  FILL_800
timestamp 1745462530
transform 1 0 808 0 1 3370
box -8 -3 16 105
use FILL  FILL_801
timestamp 1745462530
transform 1 0 800 0 1 3370
box -8 -3 16 105
use FILL  FILL_802
timestamp 1745462530
transform 1 0 696 0 1 3370
box -8 -3 16 105
use FILL  FILL_803
timestamp 1745462530
transform 1 0 688 0 1 3370
box -8 -3 16 105
use FILL  FILL_804
timestamp 1745462530
transform 1 0 584 0 1 3370
box -8 -3 16 105
use FILL  FILL_805
timestamp 1745462530
transform 1 0 480 0 1 3370
box -8 -3 16 105
use FILL  FILL_806
timestamp 1745462530
transform 1 0 472 0 1 3370
box -8 -3 16 105
use FILL  FILL_807
timestamp 1745462530
transform 1 0 464 0 1 3370
box -8 -3 16 105
use FILL  FILL_808
timestamp 1745462530
transform 1 0 360 0 1 3370
box -8 -3 16 105
use FILL  FILL_809
timestamp 1745462530
transform 1 0 296 0 1 3370
box -8 -3 16 105
use FILL  FILL_810
timestamp 1745462530
transform 1 0 288 0 1 3370
box -8 -3 16 105
use FILL  FILL_811
timestamp 1745462530
transform 1 0 232 0 1 3370
box -8 -3 16 105
use FILL  FILL_812
timestamp 1745462530
transform 1 0 176 0 1 3370
box -8 -3 16 105
use FILL  FILL_813
timestamp 1745462530
transform 1 0 72 0 1 3370
box -8 -3 16 105
use FILL  FILL_814
timestamp 1745462530
transform 1 0 4256 0 -1 3370
box -8 -3 16 105
use FILL  FILL_815
timestamp 1745462530
transform 1 0 4080 0 -1 3370
box -8 -3 16 105
use FILL  FILL_816
timestamp 1745462530
transform 1 0 3904 0 -1 3370
box -8 -3 16 105
use FILL  FILL_817
timestamp 1745462530
transform 1 0 3896 0 -1 3370
box -8 -3 16 105
use FILL  FILL_818
timestamp 1745462530
transform 1 0 3840 0 -1 3370
box -8 -3 16 105
use FILL  FILL_819
timestamp 1745462530
transform 1 0 3800 0 -1 3370
box -8 -3 16 105
use FILL  FILL_820
timestamp 1745462530
transform 1 0 3760 0 -1 3370
box -8 -3 16 105
use FILL  FILL_821
timestamp 1745462530
transform 1 0 3688 0 -1 3370
box -8 -3 16 105
use FILL  FILL_822
timestamp 1745462530
transform 1 0 3680 0 -1 3370
box -8 -3 16 105
use FILL  FILL_823
timestamp 1745462530
transform 1 0 3608 0 -1 3370
box -8 -3 16 105
use FILL  FILL_824
timestamp 1745462530
transform 1 0 3568 0 -1 3370
box -8 -3 16 105
use FILL  FILL_825
timestamp 1745462530
transform 1 0 3528 0 -1 3370
box -8 -3 16 105
use FILL  FILL_826
timestamp 1745462530
transform 1 0 3480 0 -1 3370
box -8 -3 16 105
use FILL  FILL_827
timestamp 1745462530
transform 1 0 3432 0 -1 3370
box -8 -3 16 105
use FILL  FILL_828
timestamp 1745462530
transform 1 0 3384 0 -1 3370
box -8 -3 16 105
use FILL  FILL_829
timestamp 1745462530
transform 1 0 3336 0 -1 3370
box -8 -3 16 105
use FILL  FILL_830
timestamp 1745462530
transform 1 0 3296 0 -1 3370
box -8 -3 16 105
use FILL  FILL_831
timestamp 1745462530
transform 1 0 3256 0 -1 3370
box -8 -3 16 105
use FILL  FILL_832
timestamp 1745462530
transform 1 0 3208 0 -1 3370
box -8 -3 16 105
use FILL  FILL_833
timestamp 1745462530
transform 1 0 3160 0 -1 3370
box -8 -3 16 105
use FILL  FILL_834
timestamp 1745462530
transform 1 0 3120 0 -1 3370
box -8 -3 16 105
use FILL  FILL_835
timestamp 1745462530
transform 1 0 3112 0 -1 3370
box -8 -3 16 105
use FILL  FILL_836
timestamp 1745462530
transform 1 0 3072 0 -1 3370
box -8 -3 16 105
use FILL  FILL_837
timestamp 1745462530
transform 1 0 3064 0 -1 3370
box -8 -3 16 105
use FILL  FILL_838
timestamp 1745462530
transform 1 0 3008 0 -1 3370
box -8 -3 16 105
use FILL  FILL_839
timestamp 1745462530
transform 1 0 3000 0 -1 3370
box -8 -3 16 105
use FILL  FILL_840
timestamp 1745462530
transform 1 0 2920 0 -1 3370
box -8 -3 16 105
use FILL  FILL_841
timestamp 1745462530
transform 1 0 2912 0 -1 3370
box -8 -3 16 105
use FILL  FILL_842
timestamp 1745462530
transform 1 0 2904 0 -1 3370
box -8 -3 16 105
use FILL  FILL_843
timestamp 1745462530
transform 1 0 2856 0 -1 3370
box -8 -3 16 105
use FILL  FILL_844
timestamp 1745462530
transform 1 0 2848 0 -1 3370
box -8 -3 16 105
use FILL  FILL_845
timestamp 1745462530
transform 1 0 2808 0 -1 3370
box -8 -3 16 105
use FILL  FILL_846
timestamp 1745462530
transform 1 0 2800 0 -1 3370
box -8 -3 16 105
use FILL  FILL_847
timestamp 1745462530
transform 1 0 2792 0 -1 3370
box -8 -3 16 105
use FILL  FILL_848
timestamp 1745462530
transform 1 0 2744 0 -1 3370
box -8 -3 16 105
use FILL  FILL_849
timestamp 1745462530
transform 1 0 2736 0 -1 3370
box -8 -3 16 105
use FILL  FILL_850
timestamp 1745462530
transform 1 0 2696 0 -1 3370
box -8 -3 16 105
use FILL  FILL_851
timestamp 1745462530
transform 1 0 2688 0 -1 3370
box -8 -3 16 105
use FILL  FILL_852
timestamp 1745462530
transform 1 0 2656 0 -1 3370
box -8 -3 16 105
use FILL  FILL_853
timestamp 1745462530
transform 1 0 2616 0 -1 3370
box -8 -3 16 105
use FILL  FILL_854
timestamp 1745462530
transform 1 0 2608 0 -1 3370
box -8 -3 16 105
use FILL  FILL_855
timestamp 1745462530
transform 1 0 2600 0 -1 3370
box -8 -3 16 105
use FILL  FILL_856
timestamp 1745462530
transform 1 0 2552 0 -1 3370
box -8 -3 16 105
use FILL  FILL_857
timestamp 1745462530
transform 1 0 2544 0 -1 3370
box -8 -3 16 105
use FILL  FILL_858
timestamp 1745462530
transform 1 0 2536 0 -1 3370
box -8 -3 16 105
use FILL  FILL_859
timestamp 1745462530
transform 1 0 2488 0 -1 3370
box -8 -3 16 105
use FILL  FILL_860
timestamp 1745462530
transform 1 0 2480 0 -1 3370
box -8 -3 16 105
use FILL  FILL_861
timestamp 1745462530
transform 1 0 2472 0 -1 3370
box -8 -3 16 105
use FILL  FILL_862
timestamp 1745462530
transform 1 0 2432 0 -1 3370
box -8 -3 16 105
use FILL  FILL_863
timestamp 1745462530
transform 1 0 2424 0 -1 3370
box -8 -3 16 105
use FILL  FILL_864
timestamp 1745462530
transform 1 0 2416 0 -1 3370
box -8 -3 16 105
use FILL  FILL_865
timestamp 1745462530
transform 1 0 2376 0 -1 3370
box -8 -3 16 105
use FILL  FILL_866
timestamp 1745462530
transform 1 0 2368 0 -1 3370
box -8 -3 16 105
use FILL  FILL_867
timestamp 1745462530
transform 1 0 2360 0 -1 3370
box -8 -3 16 105
use FILL  FILL_868
timestamp 1745462530
transform 1 0 2320 0 -1 3370
box -8 -3 16 105
use FILL  FILL_869
timestamp 1745462530
transform 1 0 2312 0 -1 3370
box -8 -3 16 105
use FILL  FILL_870
timestamp 1745462530
transform 1 0 2304 0 -1 3370
box -8 -3 16 105
use FILL  FILL_871
timestamp 1745462530
transform 1 0 2264 0 -1 3370
box -8 -3 16 105
use FILL  FILL_872
timestamp 1745462530
transform 1 0 2256 0 -1 3370
box -8 -3 16 105
use FILL  FILL_873
timestamp 1745462530
transform 1 0 2216 0 -1 3370
box -8 -3 16 105
use FILL  FILL_874
timestamp 1745462530
transform 1 0 2208 0 -1 3370
box -8 -3 16 105
use FILL  FILL_875
timestamp 1745462530
transform 1 0 2184 0 -1 3370
box -8 -3 16 105
use FILL  FILL_876
timestamp 1745462530
transform 1 0 2176 0 -1 3370
box -8 -3 16 105
use FILL  FILL_877
timestamp 1745462530
transform 1 0 2144 0 -1 3370
box -8 -3 16 105
use FILL  FILL_878
timestamp 1745462530
transform 1 0 2112 0 -1 3370
box -8 -3 16 105
use FILL  FILL_879
timestamp 1745462530
transform 1 0 2104 0 -1 3370
box -8 -3 16 105
use FILL  FILL_880
timestamp 1745462530
transform 1 0 2096 0 -1 3370
box -8 -3 16 105
use FILL  FILL_881
timestamp 1745462530
transform 1 0 2056 0 -1 3370
box -8 -3 16 105
use FILL  FILL_882
timestamp 1745462530
transform 1 0 2048 0 -1 3370
box -8 -3 16 105
use FILL  FILL_883
timestamp 1745462530
transform 1 0 2016 0 -1 3370
box -8 -3 16 105
use FILL  FILL_884
timestamp 1745462530
transform 1 0 2008 0 -1 3370
box -8 -3 16 105
use FILL  FILL_885
timestamp 1745462530
transform 1 0 1968 0 -1 3370
box -8 -3 16 105
use FILL  FILL_886
timestamp 1745462530
transform 1 0 1960 0 -1 3370
box -8 -3 16 105
use FILL  FILL_887
timestamp 1745462530
transform 1 0 1952 0 -1 3370
box -8 -3 16 105
use FILL  FILL_888
timestamp 1745462530
transform 1 0 1920 0 -1 3370
box -8 -3 16 105
use FILL  FILL_889
timestamp 1745462530
transform 1 0 1888 0 -1 3370
box -8 -3 16 105
use FILL  FILL_890
timestamp 1745462530
transform 1 0 1880 0 -1 3370
box -8 -3 16 105
use FILL  FILL_891
timestamp 1745462530
transform 1 0 1840 0 -1 3370
box -8 -3 16 105
use FILL  FILL_892
timestamp 1745462530
transform 1 0 1832 0 -1 3370
box -8 -3 16 105
use FILL  FILL_893
timestamp 1745462530
transform 1 0 1824 0 -1 3370
box -8 -3 16 105
use FILL  FILL_894
timestamp 1745462530
transform 1 0 1784 0 -1 3370
box -8 -3 16 105
use FILL  FILL_895
timestamp 1745462530
transform 1 0 1776 0 -1 3370
box -8 -3 16 105
use FILL  FILL_896
timestamp 1745462530
transform 1 0 1744 0 -1 3370
box -8 -3 16 105
use FILL  FILL_897
timestamp 1745462530
transform 1 0 1736 0 -1 3370
box -8 -3 16 105
use FILL  FILL_898
timestamp 1745462530
transform 1 0 1696 0 -1 3370
box -8 -3 16 105
use FILL  FILL_899
timestamp 1745462530
transform 1 0 1656 0 -1 3370
box -8 -3 16 105
use FILL  FILL_900
timestamp 1745462530
transform 1 0 1616 0 -1 3370
box -8 -3 16 105
use FILL  FILL_901
timestamp 1745462530
transform 1 0 1608 0 -1 3370
box -8 -3 16 105
use FILL  FILL_902
timestamp 1745462530
transform 1 0 1568 0 -1 3370
box -8 -3 16 105
use FILL  FILL_903
timestamp 1745462530
transform 1 0 1528 0 -1 3370
box -8 -3 16 105
use FILL  FILL_904
timestamp 1745462530
transform 1 0 1488 0 -1 3370
box -8 -3 16 105
use FILL  FILL_905
timestamp 1745462530
transform 1 0 1448 0 -1 3370
box -8 -3 16 105
use FILL  FILL_906
timestamp 1745462530
transform 1 0 1440 0 -1 3370
box -8 -3 16 105
use FILL  FILL_907
timestamp 1745462530
transform 1 0 1400 0 -1 3370
box -8 -3 16 105
use FILL  FILL_908
timestamp 1745462530
transform 1 0 1360 0 -1 3370
box -8 -3 16 105
use FILL  FILL_909
timestamp 1745462530
transform 1 0 1352 0 -1 3370
box -8 -3 16 105
use FILL  FILL_910
timestamp 1745462530
transform 1 0 1304 0 -1 3370
box -8 -3 16 105
use FILL  FILL_911
timestamp 1745462530
transform 1 0 1296 0 -1 3370
box -8 -3 16 105
use FILL  FILL_912
timestamp 1745462530
transform 1 0 1256 0 -1 3370
box -8 -3 16 105
use FILL  FILL_913
timestamp 1745462530
transform 1 0 1152 0 -1 3370
box -8 -3 16 105
use FILL  FILL_914
timestamp 1745462530
transform 1 0 1144 0 -1 3370
box -8 -3 16 105
use FILL  FILL_915
timestamp 1745462530
transform 1 0 1136 0 -1 3370
box -8 -3 16 105
use FILL  FILL_916
timestamp 1745462530
transform 1 0 1088 0 -1 3370
box -8 -3 16 105
use FILL  FILL_917
timestamp 1745462530
transform 1 0 1024 0 -1 3370
box -8 -3 16 105
use FILL  FILL_918
timestamp 1745462530
transform 1 0 1016 0 -1 3370
box -8 -3 16 105
use FILL  FILL_919
timestamp 1745462530
transform 1 0 1008 0 -1 3370
box -8 -3 16 105
use FILL  FILL_920
timestamp 1745462530
transform 1 0 944 0 -1 3370
box -8 -3 16 105
use FILL  FILL_921
timestamp 1745462530
transform 1 0 936 0 -1 3370
box -8 -3 16 105
use FILL  FILL_922
timestamp 1745462530
transform 1 0 832 0 -1 3370
box -8 -3 16 105
use FILL  FILL_923
timestamp 1745462530
transform 1 0 824 0 -1 3370
box -8 -3 16 105
use FILL  FILL_924
timestamp 1745462530
transform 1 0 816 0 -1 3370
box -8 -3 16 105
use FILL  FILL_925
timestamp 1745462530
transform 1 0 712 0 -1 3370
box -8 -3 16 105
use FILL  FILL_926
timestamp 1745462530
transform 1 0 704 0 -1 3370
box -8 -3 16 105
use FILL  FILL_927
timestamp 1745462530
transform 1 0 696 0 -1 3370
box -8 -3 16 105
use FILL  FILL_928
timestamp 1745462530
transform 1 0 592 0 -1 3370
box -8 -3 16 105
use FILL  FILL_929
timestamp 1745462530
transform 1 0 584 0 -1 3370
box -8 -3 16 105
use FILL  FILL_930
timestamp 1745462530
transform 1 0 480 0 -1 3370
box -8 -3 16 105
use FILL  FILL_931
timestamp 1745462530
transform 1 0 472 0 -1 3370
box -8 -3 16 105
use FILL  FILL_932
timestamp 1745462530
transform 1 0 464 0 -1 3370
box -8 -3 16 105
use FILL  FILL_933
timestamp 1745462530
transform 1 0 360 0 -1 3370
box -8 -3 16 105
use FILL  FILL_934
timestamp 1745462530
transform 1 0 352 0 -1 3370
box -8 -3 16 105
use FILL  FILL_935
timestamp 1745462530
transform 1 0 248 0 -1 3370
box -8 -3 16 105
use FILL  FILL_936
timestamp 1745462530
transform 1 0 240 0 -1 3370
box -8 -3 16 105
use FILL  FILL_937
timestamp 1745462530
transform 1 0 232 0 -1 3370
box -8 -3 16 105
use FILL  FILL_938
timestamp 1745462530
transform 1 0 128 0 -1 3370
box -8 -3 16 105
use FILL  FILL_939
timestamp 1745462530
transform 1 0 120 0 -1 3370
box -8 -3 16 105
use FILL  FILL_940
timestamp 1745462530
transform 1 0 112 0 -1 3370
box -8 -3 16 105
use FILL  FILL_941
timestamp 1745462530
transform 1 0 104 0 -1 3370
box -8 -3 16 105
use FILL  FILL_942
timestamp 1745462530
transform 1 0 96 0 -1 3370
box -8 -3 16 105
use FILL  FILL_943
timestamp 1745462530
transform 1 0 88 0 -1 3370
box -8 -3 16 105
use FILL  FILL_944
timestamp 1745462530
transform 1 0 80 0 -1 3370
box -8 -3 16 105
use FILL  FILL_945
timestamp 1745462530
transform 1 0 72 0 -1 3370
box -8 -3 16 105
use FILL  FILL_946
timestamp 1745462530
transform 1 0 4368 0 1 3170
box -8 -3 16 105
use FILL  FILL_947
timestamp 1745462530
transform 1 0 4248 0 1 3170
box -8 -3 16 105
use FILL  FILL_948
timestamp 1745462530
transform 1 0 4184 0 1 3170
box -8 -3 16 105
use FILL  FILL_949
timestamp 1745462530
transform 1 0 4064 0 1 3170
box -8 -3 16 105
use FILL  FILL_950
timestamp 1745462530
transform 1 0 4000 0 1 3170
box -8 -3 16 105
use FILL  FILL_951
timestamp 1745462530
transform 1 0 3992 0 1 3170
box -8 -3 16 105
use FILL  FILL_952
timestamp 1745462530
transform 1 0 3984 0 1 3170
box -8 -3 16 105
use FILL  FILL_953
timestamp 1745462530
transform 1 0 3920 0 1 3170
box -8 -3 16 105
use FILL  FILL_954
timestamp 1745462530
transform 1 0 3864 0 1 3170
box -8 -3 16 105
use FILL  FILL_955
timestamp 1745462530
transform 1 0 3856 0 1 3170
box -8 -3 16 105
use FILL  FILL_956
timestamp 1745462530
transform 1 0 3816 0 1 3170
box -8 -3 16 105
use FILL  FILL_957
timestamp 1745462530
transform 1 0 3776 0 1 3170
box -8 -3 16 105
use FILL  FILL_958
timestamp 1745462530
transform 1 0 3736 0 1 3170
box -8 -3 16 105
use FILL  FILL_959
timestamp 1745462530
transform 1 0 3680 0 1 3170
box -8 -3 16 105
use FILL  FILL_960
timestamp 1745462530
transform 1 0 3672 0 1 3170
box -8 -3 16 105
use FILL  FILL_961
timestamp 1745462530
transform 1 0 3632 0 1 3170
box -8 -3 16 105
use FILL  FILL_962
timestamp 1745462530
transform 1 0 3600 0 1 3170
box -8 -3 16 105
use FILL  FILL_963
timestamp 1745462530
transform 1 0 3560 0 1 3170
box -8 -3 16 105
use FILL  FILL_964
timestamp 1745462530
transform 1 0 3520 0 1 3170
box -8 -3 16 105
use FILL  FILL_965
timestamp 1745462530
transform 1 0 3512 0 1 3170
box -8 -3 16 105
use FILL  FILL_966
timestamp 1745462530
transform 1 0 3464 0 1 3170
box -8 -3 16 105
use FILL  FILL_967
timestamp 1745462530
transform 1 0 3424 0 1 3170
box -8 -3 16 105
use FILL  FILL_968
timestamp 1745462530
transform 1 0 3384 0 1 3170
box -8 -3 16 105
use FILL  FILL_969
timestamp 1745462530
transform 1 0 3376 0 1 3170
box -8 -3 16 105
use FILL  FILL_970
timestamp 1745462530
transform 1 0 3328 0 1 3170
box -8 -3 16 105
use FILL  FILL_971
timestamp 1745462530
transform 1 0 3280 0 1 3170
box -8 -3 16 105
use FILL  FILL_972
timestamp 1745462530
transform 1 0 3272 0 1 3170
box -8 -3 16 105
use FILL  FILL_973
timestamp 1745462530
transform 1 0 3208 0 1 3170
box -8 -3 16 105
use FILL  FILL_974
timestamp 1745462530
transform 1 0 3200 0 1 3170
box -8 -3 16 105
use FILL  FILL_975
timestamp 1745462530
transform 1 0 3144 0 1 3170
box -8 -3 16 105
use FILL  FILL_976
timestamp 1745462530
transform 1 0 3136 0 1 3170
box -8 -3 16 105
use FILL  FILL_977
timestamp 1745462530
transform 1 0 3128 0 1 3170
box -8 -3 16 105
use FILL  FILL_978
timestamp 1745462530
transform 1 0 3056 0 1 3170
box -8 -3 16 105
use FILL  FILL_979
timestamp 1745462530
transform 1 0 3048 0 1 3170
box -8 -3 16 105
use FILL  FILL_980
timestamp 1745462530
transform 1 0 3040 0 1 3170
box -8 -3 16 105
use FILL  FILL_981
timestamp 1745462530
transform 1 0 2984 0 1 3170
box -8 -3 16 105
use FILL  FILL_982
timestamp 1745462530
transform 1 0 2960 0 1 3170
box -8 -3 16 105
use FILL  FILL_983
timestamp 1745462530
transform 1 0 2920 0 1 3170
box -8 -3 16 105
use FILL  FILL_984
timestamp 1745462530
transform 1 0 2912 0 1 3170
box -8 -3 16 105
use FILL  FILL_985
timestamp 1745462530
transform 1 0 2864 0 1 3170
box -8 -3 16 105
use FILL  FILL_986
timestamp 1745462530
transform 1 0 2856 0 1 3170
box -8 -3 16 105
use FILL  FILL_987
timestamp 1745462530
transform 1 0 2816 0 1 3170
box -8 -3 16 105
use FILL  FILL_988
timestamp 1745462530
transform 1 0 2808 0 1 3170
box -8 -3 16 105
use FILL  FILL_989
timestamp 1745462530
transform 1 0 2800 0 1 3170
box -8 -3 16 105
use FILL  FILL_990
timestamp 1745462530
transform 1 0 2752 0 1 3170
box -8 -3 16 105
use FILL  FILL_991
timestamp 1745462530
transform 1 0 2744 0 1 3170
box -8 -3 16 105
use FILL  FILL_992
timestamp 1745462530
transform 1 0 2696 0 1 3170
box -8 -3 16 105
use FILL  FILL_993
timestamp 1745462530
transform 1 0 2688 0 1 3170
box -8 -3 16 105
use FILL  FILL_994
timestamp 1745462530
transform 1 0 2648 0 1 3170
box -8 -3 16 105
use FILL  FILL_995
timestamp 1745462530
transform 1 0 2640 0 1 3170
box -8 -3 16 105
use FILL  FILL_996
timestamp 1745462530
transform 1 0 2632 0 1 3170
box -8 -3 16 105
use FILL  FILL_997
timestamp 1745462530
transform 1 0 2592 0 1 3170
box -8 -3 16 105
use FILL  FILL_998
timestamp 1745462530
transform 1 0 2584 0 1 3170
box -8 -3 16 105
use FILL  FILL_999
timestamp 1745462530
transform 1 0 2576 0 1 3170
box -8 -3 16 105
use FILL  FILL_1000
timestamp 1745462530
transform 1 0 2528 0 1 3170
box -8 -3 16 105
use FILL  FILL_1001
timestamp 1745462530
transform 1 0 2520 0 1 3170
box -8 -3 16 105
use FILL  FILL_1002
timestamp 1745462530
transform 1 0 2512 0 1 3170
box -8 -3 16 105
use FILL  FILL_1003
timestamp 1745462530
transform 1 0 2472 0 1 3170
box -8 -3 16 105
use FILL  FILL_1004
timestamp 1745462530
transform 1 0 2464 0 1 3170
box -8 -3 16 105
use FILL  FILL_1005
timestamp 1745462530
transform 1 0 2456 0 1 3170
box -8 -3 16 105
use FILL  FILL_1006
timestamp 1745462530
transform 1 0 2408 0 1 3170
box -8 -3 16 105
use FILL  FILL_1007
timestamp 1745462530
transform 1 0 2400 0 1 3170
box -8 -3 16 105
use FILL  FILL_1008
timestamp 1745462530
transform 1 0 2392 0 1 3170
box -8 -3 16 105
use FILL  FILL_1009
timestamp 1745462530
transform 1 0 2352 0 1 3170
box -8 -3 16 105
use FILL  FILL_1010
timestamp 1745462530
transform 1 0 2344 0 1 3170
box -8 -3 16 105
use FILL  FILL_1011
timestamp 1745462530
transform 1 0 2304 0 1 3170
box -8 -3 16 105
use FILL  FILL_1012
timestamp 1745462530
transform 1 0 2296 0 1 3170
box -8 -3 16 105
use FILL  FILL_1013
timestamp 1745462530
transform 1 0 2288 0 1 3170
box -8 -3 16 105
use FILL  FILL_1014
timestamp 1745462530
transform 1 0 2256 0 1 3170
box -8 -3 16 105
use FILL  FILL_1015
timestamp 1745462530
transform 1 0 2224 0 1 3170
box -8 -3 16 105
use FILL  FILL_1016
timestamp 1745462530
transform 1 0 2216 0 1 3170
box -8 -3 16 105
use FILL  FILL_1017
timestamp 1745462530
transform 1 0 2176 0 1 3170
box -8 -3 16 105
use FILL  FILL_1018
timestamp 1745462530
transform 1 0 2168 0 1 3170
box -8 -3 16 105
use FILL  FILL_1019
timestamp 1745462530
transform 1 0 2160 0 1 3170
box -8 -3 16 105
use FILL  FILL_1020
timestamp 1745462530
transform 1 0 2120 0 1 3170
box -8 -3 16 105
use FILL  FILL_1021
timestamp 1745462530
transform 1 0 2112 0 1 3170
box -8 -3 16 105
use FILL  FILL_1022
timestamp 1745462530
transform 1 0 2080 0 1 3170
box -8 -3 16 105
use FILL  FILL_1023
timestamp 1745462530
transform 1 0 2072 0 1 3170
box -8 -3 16 105
use FILL  FILL_1024
timestamp 1745462530
transform 1 0 2040 0 1 3170
box -8 -3 16 105
use FILL  FILL_1025
timestamp 1745462530
transform 1 0 2008 0 1 3170
box -8 -3 16 105
use FILL  FILL_1026
timestamp 1745462530
transform 1 0 2000 0 1 3170
box -8 -3 16 105
use FILL  FILL_1027
timestamp 1745462530
transform 1 0 1992 0 1 3170
box -8 -3 16 105
use FILL  FILL_1028
timestamp 1745462530
transform 1 0 1952 0 1 3170
box -8 -3 16 105
use FILL  FILL_1029
timestamp 1745462530
transform 1 0 1944 0 1 3170
box -8 -3 16 105
use FILL  FILL_1030
timestamp 1745462530
transform 1 0 1904 0 1 3170
box -8 -3 16 105
use FILL  FILL_1031
timestamp 1745462530
transform 1 0 1896 0 1 3170
box -8 -3 16 105
use FILL  FILL_1032
timestamp 1745462530
transform 1 0 1888 0 1 3170
box -8 -3 16 105
use FILL  FILL_1033
timestamp 1745462530
transform 1 0 1856 0 1 3170
box -8 -3 16 105
use FILL  FILL_1034
timestamp 1745462530
transform 1 0 1848 0 1 3170
box -8 -3 16 105
use FILL  FILL_1035
timestamp 1745462530
transform 1 0 1808 0 1 3170
box -8 -3 16 105
use FILL  FILL_1036
timestamp 1745462530
transform 1 0 1800 0 1 3170
box -8 -3 16 105
use FILL  FILL_1037
timestamp 1745462530
transform 1 0 1760 0 1 3170
box -8 -3 16 105
use FILL  FILL_1038
timestamp 1745462530
transform 1 0 1720 0 1 3170
box -8 -3 16 105
use FILL  FILL_1039
timestamp 1745462530
transform 1 0 1680 0 1 3170
box -8 -3 16 105
use FILL  FILL_1040
timestamp 1745462530
transform 1 0 1640 0 1 3170
box -8 -3 16 105
use FILL  FILL_1041
timestamp 1745462530
transform 1 0 1632 0 1 3170
box -8 -3 16 105
use FILL  FILL_1042
timestamp 1745462530
transform 1 0 1576 0 1 3170
box -8 -3 16 105
use FILL  FILL_1043
timestamp 1745462530
transform 1 0 1552 0 1 3170
box -8 -3 16 105
use FILL  FILL_1044
timestamp 1745462530
transform 1 0 1496 0 1 3170
box -8 -3 16 105
use FILL  FILL_1045
timestamp 1745462530
transform 1 0 1488 0 1 3170
box -8 -3 16 105
use FILL  FILL_1046
timestamp 1745462530
transform 1 0 1384 0 1 3170
box -8 -3 16 105
use FILL  FILL_1047
timestamp 1745462530
transform 1 0 1344 0 1 3170
box -8 -3 16 105
use FILL  FILL_1048
timestamp 1745462530
transform 1 0 1304 0 1 3170
box -8 -3 16 105
use FILL  FILL_1049
timestamp 1745462530
transform 1 0 1296 0 1 3170
box -8 -3 16 105
use FILL  FILL_1050
timestamp 1745462530
transform 1 0 1240 0 1 3170
box -8 -3 16 105
use FILL  FILL_1051
timestamp 1745462530
transform 1 0 1232 0 1 3170
box -8 -3 16 105
use FILL  FILL_1052
timestamp 1745462530
transform 1 0 1128 0 1 3170
box -8 -3 16 105
use FILL  FILL_1053
timestamp 1745462530
transform 1 0 1120 0 1 3170
box -8 -3 16 105
use FILL  FILL_1054
timestamp 1745462530
transform 1 0 1080 0 1 3170
box -8 -3 16 105
use FILL  FILL_1055
timestamp 1745462530
transform 1 0 1056 0 1 3170
box -8 -3 16 105
use FILL  FILL_1056
timestamp 1745462530
transform 1 0 1016 0 1 3170
box -8 -3 16 105
use FILL  FILL_1057
timestamp 1745462530
transform 1 0 1008 0 1 3170
box -8 -3 16 105
use FILL  FILL_1058
timestamp 1745462530
transform 1 0 960 0 1 3170
box -8 -3 16 105
use FILL  FILL_1059
timestamp 1745462530
transform 1 0 952 0 1 3170
box -8 -3 16 105
use FILL  FILL_1060
timestamp 1745462530
transform 1 0 944 0 1 3170
box -8 -3 16 105
use FILL  FILL_1061
timestamp 1745462530
transform 1 0 904 0 1 3170
box -8 -3 16 105
use FILL  FILL_1062
timestamp 1745462530
transform 1 0 896 0 1 3170
box -8 -3 16 105
use FILL  FILL_1063
timestamp 1745462530
transform 1 0 848 0 1 3170
box -8 -3 16 105
use FILL  FILL_1064
timestamp 1745462530
transform 1 0 840 0 1 3170
box -8 -3 16 105
use FILL  FILL_1065
timestamp 1745462530
transform 1 0 832 0 1 3170
box -8 -3 16 105
use FILL  FILL_1066
timestamp 1745462530
transform 1 0 768 0 1 3170
box -8 -3 16 105
use FILL  FILL_1067
timestamp 1745462530
transform 1 0 760 0 1 3170
box -8 -3 16 105
use FILL  FILL_1068
timestamp 1745462530
transform 1 0 752 0 1 3170
box -8 -3 16 105
use FILL  FILL_1069
timestamp 1745462530
transform 1 0 744 0 1 3170
box -8 -3 16 105
use FILL  FILL_1070
timestamp 1745462530
transform 1 0 688 0 1 3170
box -8 -3 16 105
use FILL  FILL_1071
timestamp 1745462530
transform 1 0 680 0 1 3170
box -8 -3 16 105
use FILL  FILL_1072
timestamp 1745462530
transform 1 0 640 0 1 3170
box -8 -3 16 105
use FILL  FILL_1073
timestamp 1745462530
transform 1 0 632 0 1 3170
box -8 -3 16 105
use FILL  FILL_1074
timestamp 1745462530
transform 1 0 592 0 1 3170
box -8 -3 16 105
use FILL  FILL_1075
timestamp 1745462530
transform 1 0 584 0 1 3170
box -8 -3 16 105
use FILL  FILL_1076
timestamp 1745462530
transform 1 0 536 0 1 3170
box -8 -3 16 105
use FILL  FILL_1077
timestamp 1745462530
transform 1 0 528 0 1 3170
box -8 -3 16 105
use FILL  FILL_1078
timestamp 1745462530
transform 1 0 496 0 1 3170
box -8 -3 16 105
use FILL  FILL_1079
timestamp 1745462530
transform 1 0 488 0 1 3170
box -8 -3 16 105
use FILL  FILL_1080
timestamp 1745462530
transform 1 0 480 0 1 3170
box -8 -3 16 105
use FILL  FILL_1081
timestamp 1745462530
transform 1 0 432 0 1 3170
box -8 -3 16 105
use FILL  FILL_1082
timestamp 1745462530
transform 1 0 424 0 1 3170
box -8 -3 16 105
use FILL  FILL_1083
timestamp 1745462530
transform 1 0 400 0 1 3170
box -8 -3 16 105
use FILL  FILL_1084
timestamp 1745462530
transform 1 0 392 0 1 3170
box -8 -3 16 105
use FILL  FILL_1085
timestamp 1745462530
transform 1 0 384 0 1 3170
box -8 -3 16 105
use FILL  FILL_1086
timestamp 1745462530
transform 1 0 336 0 1 3170
box -8 -3 16 105
use FILL  FILL_1087
timestamp 1745462530
transform 1 0 328 0 1 3170
box -8 -3 16 105
use FILL  FILL_1088
timestamp 1745462530
transform 1 0 320 0 1 3170
box -8 -3 16 105
use FILL  FILL_1089
timestamp 1745462530
transform 1 0 296 0 1 3170
box -8 -3 16 105
use FILL  FILL_1090
timestamp 1745462530
transform 1 0 288 0 1 3170
box -8 -3 16 105
use FILL  FILL_1091
timestamp 1745462530
transform 1 0 280 0 1 3170
box -8 -3 16 105
use FILL  FILL_1092
timestamp 1745462530
transform 1 0 272 0 1 3170
box -8 -3 16 105
use FILL  FILL_1093
timestamp 1745462530
transform 1 0 224 0 1 3170
box -8 -3 16 105
use FILL  FILL_1094
timestamp 1745462530
transform 1 0 200 0 1 3170
box -8 -3 16 105
use FILL  FILL_1095
timestamp 1745462530
transform 1 0 192 0 1 3170
box -8 -3 16 105
use FILL  FILL_1096
timestamp 1745462530
transform 1 0 184 0 1 3170
box -8 -3 16 105
use FILL  FILL_1097
timestamp 1745462530
transform 1 0 176 0 1 3170
box -8 -3 16 105
use FILL  FILL_1098
timestamp 1745462530
transform 1 0 72 0 1 3170
box -8 -3 16 105
use FILL  FILL_1099
timestamp 1745462530
transform 1 0 4368 0 -1 3170
box -8 -3 16 105
use FILL  FILL_1100
timestamp 1745462530
transform 1 0 4264 0 -1 3170
box -8 -3 16 105
use FILL  FILL_1101
timestamp 1745462530
transform 1 0 4256 0 -1 3170
box -8 -3 16 105
use FILL  FILL_1102
timestamp 1745462530
transform 1 0 4192 0 -1 3170
box -8 -3 16 105
use FILL  FILL_1103
timestamp 1745462530
transform 1 0 4168 0 -1 3170
box -8 -3 16 105
use FILL  FILL_1104
timestamp 1745462530
transform 1 0 4064 0 -1 3170
box -8 -3 16 105
use FILL  FILL_1105
timestamp 1745462530
transform 1 0 4056 0 -1 3170
box -8 -3 16 105
use FILL  FILL_1106
timestamp 1745462530
transform 1 0 4048 0 -1 3170
box -8 -3 16 105
use FILL  FILL_1107
timestamp 1745462530
transform 1 0 3992 0 -1 3170
box -8 -3 16 105
use FILL  FILL_1108
timestamp 1745462530
transform 1 0 3984 0 -1 3170
box -8 -3 16 105
use FILL  FILL_1109
timestamp 1745462530
transform 1 0 3976 0 -1 3170
box -8 -3 16 105
use FILL  FILL_1110
timestamp 1745462530
transform 1 0 3920 0 -1 3170
box -8 -3 16 105
use FILL  FILL_1111
timestamp 1745462530
transform 1 0 3912 0 -1 3170
box -8 -3 16 105
use FILL  FILL_1112
timestamp 1745462530
transform 1 0 3904 0 -1 3170
box -8 -3 16 105
use FILL  FILL_1113
timestamp 1745462530
transform 1 0 3800 0 -1 3170
box -8 -3 16 105
use FILL  FILL_1114
timestamp 1745462530
transform 1 0 3792 0 -1 3170
box -8 -3 16 105
use FILL  FILL_1115
timestamp 1745462530
transform 1 0 3784 0 -1 3170
box -8 -3 16 105
use FILL  FILL_1116
timestamp 1745462530
transform 1 0 3752 0 -1 3170
box -8 -3 16 105
use FILL  FILL_1117
timestamp 1745462530
transform 1 0 3744 0 -1 3170
box -8 -3 16 105
use FILL  FILL_1118
timestamp 1745462530
transform 1 0 3736 0 -1 3170
box -8 -3 16 105
use FILL  FILL_1119
timestamp 1745462530
transform 1 0 3632 0 -1 3170
box -8 -3 16 105
use FILL  FILL_1120
timestamp 1745462530
transform 1 0 3624 0 -1 3170
box -8 -3 16 105
use FILL  FILL_1121
timestamp 1745462530
transform 1 0 3616 0 -1 3170
box -8 -3 16 105
use FILL  FILL_1122
timestamp 1745462530
transform 1 0 3576 0 -1 3170
box -8 -3 16 105
use FILL  FILL_1123
timestamp 1745462530
transform 1 0 3568 0 -1 3170
box -8 -3 16 105
use FILL  FILL_1124
timestamp 1745462530
transform 1 0 3528 0 -1 3170
box -8 -3 16 105
use FILL  FILL_1125
timestamp 1745462530
transform 1 0 3520 0 -1 3170
box -8 -3 16 105
use FILL  FILL_1126
timestamp 1745462530
transform 1 0 3472 0 -1 3170
box -8 -3 16 105
use FILL  FILL_1127
timestamp 1745462530
transform 1 0 3464 0 -1 3170
box -8 -3 16 105
use FILL  FILL_1128
timestamp 1745462530
transform 1 0 3416 0 -1 3170
box -8 -3 16 105
use FILL  FILL_1129
timestamp 1745462530
transform 1 0 3408 0 -1 3170
box -8 -3 16 105
use FILL  FILL_1130
timestamp 1745462530
transform 1 0 3360 0 -1 3170
box -8 -3 16 105
use FILL  FILL_1131
timestamp 1745462530
transform 1 0 3352 0 -1 3170
box -8 -3 16 105
use FILL  FILL_1132
timestamp 1745462530
transform 1 0 3312 0 -1 3170
box -8 -3 16 105
use FILL  FILL_1133
timestamp 1745462530
transform 1 0 3304 0 -1 3170
box -8 -3 16 105
use FILL  FILL_1134
timestamp 1745462530
transform 1 0 3256 0 -1 3170
box -8 -3 16 105
use FILL  FILL_1135
timestamp 1745462530
transform 1 0 3248 0 -1 3170
box -8 -3 16 105
use FILL  FILL_1136
timestamp 1745462530
transform 1 0 3200 0 -1 3170
box -8 -3 16 105
use FILL  FILL_1137
timestamp 1745462530
transform 1 0 3192 0 -1 3170
box -8 -3 16 105
use FILL  FILL_1138
timestamp 1745462530
transform 1 0 3168 0 -1 3170
box -8 -3 16 105
use FILL  FILL_1139
timestamp 1745462530
transform 1 0 3128 0 -1 3170
box -8 -3 16 105
use FILL  FILL_1140
timestamp 1745462530
transform 1 0 3104 0 -1 3170
box -8 -3 16 105
use FILL  FILL_1141
timestamp 1745462530
transform 1 0 3096 0 -1 3170
box -8 -3 16 105
use FILL  FILL_1142
timestamp 1745462530
transform 1 0 3056 0 -1 3170
box -8 -3 16 105
use FILL  FILL_1143
timestamp 1745462530
transform 1 0 3016 0 -1 3170
box -8 -3 16 105
use FILL  FILL_1144
timestamp 1745462530
transform 1 0 3008 0 -1 3170
box -8 -3 16 105
use FILL  FILL_1145
timestamp 1745462530
transform 1 0 2968 0 -1 3170
box -8 -3 16 105
use FILL  FILL_1146
timestamp 1745462530
transform 1 0 2944 0 -1 3170
box -8 -3 16 105
use FILL  FILL_1147
timestamp 1745462530
transform 1 0 2936 0 -1 3170
box -8 -3 16 105
use FILL  FILL_1148
timestamp 1745462530
transform 1 0 2896 0 -1 3170
box -8 -3 16 105
use FILL  FILL_1149
timestamp 1745462530
transform 1 0 2888 0 -1 3170
box -8 -3 16 105
use FILL  FILL_1150
timestamp 1745462530
transform 1 0 2880 0 -1 3170
box -8 -3 16 105
use FILL  FILL_1151
timestamp 1745462530
transform 1 0 2832 0 -1 3170
box -8 -3 16 105
use FILL  FILL_1152
timestamp 1745462530
transform 1 0 2824 0 -1 3170
box -8 -3 16 105
use FILL  FILL_1153
timestamp 1745462530
transform 1 0 2816 0 -1 3170
box -8 -3 16 105
use FILL  FILL_1154
timestamp 1745462530
transform 1 0 2760 0 -1 3170
box -8 -3 16 105
use FILL  FILL_1155
timestamp 1745462530
transform 1 0 2752 0 -1 3170
box -8 -3 16 105
use FILL  FILL_1156
timestamp 1745462530
transform 1 0 2712 0 -1 3170
box -8 -3 16 105
use FILL  FILL_1157
timestamp 1745462530
transform 1 0 2704 0 -1 3170
box -8 -3 16 105
use FILL  FILL_1158
timestamp 1745462530
transform 1 0 2648 0 -1 3170
box -8 -3 16 105
use FILL  FILL_1159
timestamp 1745462530
transform 1 0 2640 0 -1 3170
box -8 -3 16 105
use FILL  FILL_1160
timestamp 1745462530
transform 1 0 2632 0 -1 3170
box -8 -3 16 105
use FILL  FILL_1161
timestamp 1745462530
transform 1 0 2560 0 -1 3170
box -8 -3 16 105
use FILL  FILL_1162
timestamp 1745462530
transform 1 0 2552 0 -1 3170
box -8 -3 16 105
use FILL  FILL_1163
timestamp 1745462530
transform 1 0 2544 0 -1 3170
box -8 -3 16 105
use FILL  FILL_1164
timestamp 1745462530
transform 1 0 2496 0 -1 3170
box -8 -3 16 105
use FILL  FILL_1165
timestamp 1745462530
transform 1 0 2488 0 -1 3170
box -8 -3 16 105
use FILL  FILL_1166
timestamp 1745462530
transform 1 0 2464 0 -1 3170
box -8 -3 16 105
use FILL  FILL_1167
timestamp 1745462530
transform 1 0 2416 0 -1 3170
box -8 -3 16 105
use FILL  FILL_1168
timestamp 1745462530
transform 1 0 2408 0 -1 3170
box -8 -3 16 105
use FILL  FILL_1169
timestamp 1745462530
transform 1 0 2400 0 -1 3170
box -8 -3 16 105
use FILL  FILL_1170
timestamp 1745462530
transform 1 0 2368 0 -1 3170
box -8 -3 16 105
use FILL  FILL_1171
timestamp 1745462530
transform 1 0 2328 0 -1 3170
box -8 -3 16 105
use FILL  FILL_1172
timestamp 1745462530
transform 1 0 2320 0 -1 3170
box -8 -3 16 105
use FILL  FILL_1173
timestamp 1745462530
transform 1 0 2312 0 -1 3170
box -8 -3 16 105
use FILL  FILL_1174
timestamp 1745462530
transform 1 0 2304 0 -1 3170
box -8 -3 16 105
use FILL  FILL_1175
timestamp 1745462530
transform 1 0 2264 0 -1 3170
box -8 -3 16 105
use FILL  FILL_1176
timestamp 1745462530
transform 1 0 2256 0 -1 3170
box -8 -3 16 105
use FILL  FILL_1177
timestamp 1745462530
transform 1 0 2224 0 -1 3170
box -8 -3 16 105
use FILL  FILL_1178
timestamp 1745462530
transform 1 0 2192 0 -1 3170
box -8 -3 16 105
use FILL  FILL_1179
timestamp 1745462530
transform 1 0 2160 0 -1 3170
box -8 -3 16 105
use FILL  FILL_1180
timestamp 1745462530
transform 1 0 2152 0 -1 3170
box -8 -3 16 105
use FILL  FILL_1181
timestamp 1745462530
transform 1 0 2096 0 -1 3170
box -8 -3 16 105
use FILL  FILL_1182
timestamp 1745462530
transform 1 0 2088 0 -1 3170
box -8 -3 16 105
use FILL  FILL_1183
timestamp 1745462530
transform 1 0 2008 0 -1 3170
box -8 -3 16 105
use FILL  FILL_1184
timestamp 1745462530
transform 1 0 2000 0 -1 3170
box -8 -3 16 105
use FILL  FILL_1185
timestamp 1745462530
transform 1 0 1944 0 -1 3170
box -8 -3 16 105
use FILL  FILL_1186
timestamp 1745462530
transform 1 0 1936 0 -1 3170
box -8 -3 16 105
use FILL  FILL_1187
timestamp 1745462530
transform 1 0 1880 0 -1 3170
box -8 -3 16 105
use FILL  FILL_1188
timestamp 1745462530
transform 1 0 1872 0 -1 3170
box -8 -3 16 105
use FILL  FILL_1189
timestamp 1745462530
transform 1 0 1864 0 -1 3170
box -8 -3 16 105
use FILL  FILL_1190
timestamp 1745462530
transform 1 0 1808 0 -1 3170
box -8 -3 16 105
use FILL  FILL_1191
timestamp 1745462530
transform 1 0 1744 0 -1 3170
box -8 -3 16 105
use FILL  FILL_1192
timestamp 1745462530
transform 1 0 1736 0 -1 3170
box -8 -3 16 105
use FILL  FILL_1193
timestamp 1745462530
transform 1 0 1728 0 -1 3170
box -8 -3 16 105
use FILL  FILL_1194
timestamp 1745462530
transform 1 0 1648 0 -1 3170
box -8 -3 16 105
use FILL  FILL_1195
timestamp 1745462530
transform 1 0 1600 0 -1 3170
box -8 -3 16 105
use FILL  FILL_1196
timestamp 1745462530
transform 1 0 1552 0 -1 3170
box -8 -3 16 105
use FILL  FILL_1197
timestamp 1745462530
transform 1 0 1448 0 -1 3170
box -8 -3 16 105
use FILL  FILL_1198
timestamp 1745462530
transform 1 0 1408 0 -1 3170
box -8 -3 16 105
use FILL  FILL_1199
timestamp 1745462530
transform 1 0 1368 0 -1 3170
box -8 -3 16 105
use FILL  FILL_1200
timestamp 1745462530
transform 1 0 1344 0 -1 3170
box -8 -3 16 105
use FILL  FILL_1201
timestamp 1745462530
transform 1 0 1296 0 -1 3170
box -8 -3 16 105
use FILL  FILL_1202
timestamp 1745462530
transform 1 0 1264 0 -1 3170
box -8 -3 16 105
use FILL  FILL_1203
timestamp 1745462530
transform 1 0 1160 0 -1 3170
box -8 -3 16 105
use FILL  FILL_1204
timestamp 1745462530
transform 1 0 1128 0 -1 3170
box -8 -3 16 105
use FILL  FILL_1205
timestamp 1745462530
transform 1 0 1024 0 -1 3170
box -8 -3 16 105
use FILL  FILL_1206
timestamp 1745462530
transform 1 0 968 0 -1 3170
box -8 -3 16 105
use FILL  FILL_1207
timestamp 1745462530
transform 1 0 936 0 -1 3170
box -8 -3 16 105
use FILL  FILL_1208
timestamp 1745462530
transform 1 0 880 0 -1 3170
box -8 -3 16 105
use FILL  FILL_1209
timestamp 1745462530
transform 1 0 816 0 -1 3170
box -8 -3 16 105
use FILL  FILL_1210
timestamp 1745462530
transform 1 0 776 0 -1 3170
box -8 -3 16 105
use FILL  FILL_1211
timestamp 1745462530
transform 1 0 672 0 -1 3170
box -8 -3 16 105
use FILL  FILL_1212
timestamp 1745462530
transform 1 0 664 0 -1 3170
box -8 -3 16 105
use FILL  FILL_1213
timestamp 1745462530
transform 1 0 600 0 -1 3170
box -8 -3 16 105
use FILL  FILL_1214
timestamp 1745462530
transform 1 0 560 0 -1 3170
box -8 -3 16 105
use FILL  FILL_1215
timestamp 1745462530
transform 1 0 472 0 -1 3170
box -8 -3 16 105
use FILL  FILL_1216
timestamp 1745462530
transform 1 0 384 0 -1 3170
box -8 -3 16 105
use FILL  FILL_1217
timestamp 1745462530
transform 1 0 376 0 -1 3170
box -8 -3 16 105
use FILL  FILL_1218
timestamp 1745462530
transform 1 0 368 0 -1 3170
box -8 -3 16 105
use FILL  FILL_1219
timestamp 1745462530
transform 1 0 280 0 -1 3170
box -8 -3 16 105
use FILL  FILL_1220
timestamp 1745462530
transform 1 0 272 0 -1 3170
box -8 -3 16 105
use FILL  FILL_1221
timestamp 1745462530
transform 1 0 208 0 -1 3170
box -8 -3 16 105
use FILL  FILL_1222
timestamp 1745462530
transform 1 0 200 0 -1 3170
box -8 -3 16 105
use FILL  FILL_1223
timestamp 1745462530
transform 1 0 192 0 -1 3170
box -8 -3 16 105
use FILL  FILL_1224
timestamp 1745462530
transform 1 0 184 0 -1 3170
box -8 -3 16 105
use FILL  FILL_1225
timestamp 1745462530
transform 1 0 80 0 -1 3170
box -8 -3 16 105
use FILL  FILL_1226
timestamp 1745462530
transform 1 0 72 0 -1 3170
box -8 -3 16 105
use FILL  FILL_1227
timestamp 1745462530
transform 1 0 4368 0 1 2970
box -8 -3 16 105
use FILL  FILL_1228
timestamp 1745462530
transform 1 0 4360 0 1 2970
box -8 -3 16 105
use FILL  FILL_1229
timestamp 1745462530
transform 1 0 4352 0 1 2970
box -8 -3 16 105
use FILL  FILL_1230
timestamp 1745462530
transform 1 0 4344 0 1 2970
box -8 -3 16 105
use FILL  FILL_1231
timestamp 1745462530
transform 1 0 4336 0 1 2970
box -8 -3 16 105
use FILL  FILL_1232
timestamp 1745462530
transform 1 0 4232 0 1 2970
box -8 -3 16 105
use FILL  FILL_1233
timestamp 1745462530
transform 1 0 4224 0 1 2970
box -8 -3 16 105
use FILL  FILL_1234
timestamp 1745462530
transform 1 0 4216 0 1 2970
box -8 -3 16 105
use FILL  FILL_1235
timestamp 1745462530
transform 1 0 4152 0 1 2970
box -8 -3 16 105
use FILL  FILL_1236
timestamp 1745462530
transform 1 0 4144 0 1 2970
box -8 -3 16 105
use FILL  FILL_1237
timestamp 1745462530
transform 1 0 4080 0 1 2970
box -8 -3 16 105
use FILL  FILL_1238
timestamp 1745462530
transform 1 0 3976 0 1 2970
box -8 -3 16 105
use FILL  FILL_1239
timestamp 1745462530
transform 1 0 3968 0 1 2970
box -8 -3 16 105
use FILL  FILL_1240
timestamp 1745462530
transform 1 0 3944 0 1 2970
box -8 -3 16 105
use FILL  FILL_1241
timestamp 1745462530
transform 1 0 3880 0 1 2970
box -8 -3 16 105
use FILL  FILL_1242
timestamp 1745462530
transform 1 0 3872 0 1 2970
box -8 -3 16 105
use FILL  FILL_1243
timestamp 1745462530
transform 1 0 3808 0 1 2970
box -8 -3 16 105
use FILL  FILL_1244
timestamp 1745462530
transform 1 0 3800 0 1 2970
box -8 -3 16 105
use FILL  FILL_1245
timestamp 1745462530
transform 1 0 3792 0 1 2970
box -8 -3 16 105
use FILL  FILL_1246
timestamp 1745462530
transform 1 0 3728 0 1 2970
box -8 -3 16 105
use FILL  FILL_1247
timestamp 1745462530
transform 1 0 3664 0 1 2970
box -8 -3 16 105
use FILL  FILL_1248
timestamp 1745462530
transform 1 0 3656 0 1 2970
box -8 -3 16 105
use FILL  FILL_1249
timestamp 1745462530
transform 1 0 3552 0 1 2970
box -8 -3 16 105
use FILL  FILL_1250
timestamp 1745462530
transform 1 0 3448 0 1 2970
box -8 -3 16 105
use FILL  FILL_1251
timestamp 1745462530
transform 1 0 3344 0 1 2970
box -8 -3 16 105
use FILL  FILL_1252
timestamp 1745462530
transform 1 0 3336 0 1 2970
box -8 -3 16 105
use FILL  FILL_1253
timestamp 1745462530
transform 1 0 3232 0 1 2970
box -8 -3 16 105
use FILL  FILL_1254
timestamp 1745462530
transform 1 0 3168 0 1 2970
box -8 -3 16 105
use FILL  FILL_1255
timestamp 1745462530
transform 1 0 3064 0 1 2970
box -8 -3 16 105
use FILL  FILL_1256
timestamp 1745462530
transform 1 0 2992 0 1 2970
box -8 -3 16 105
use FILL  FILL_1257
timestamp 1745462530
transform 1 0 2936 0 1 2970
box -8 -3 16 105
use FILL  FILL_1258
timestamp 1745462530
transform 1 0 2928 0 1 2970
box -8 -3 16 105
use FILL  FILL_1259
timestamp 1745462530
transform 1 0 2920 0 1 2970
box -8 -3 16 105
use FILL  FILL_1260
timestamp 1745462530
transform 1 0 2864 0 1 2970
box -8 -3 16 105
use FILL  FILL_1261
timestamp 1745462530
transform 1 0 2824 0 1 2970
box -8 -3 16 105
use FILL  FILL_1262
timestamp 1745462530
transform 1 0 2792 0 1 2970
box -8 -3 16 105
use FILL  FILL_1263
timestamp 1745462530
transform 1 0 2784 0 1 2970
box -8 -3 16 105
use FILL  FILL_1264
timestamp 1745462530
transform 1 0 2712 0 1 2970
box -8 -3 16 105
use FILL  FILL_1265
timestamp 1745462530
transform 1 0 2704 0 1 2970
box -8 -3 16 105
use FILL  FILL_1266
timestamp 1745462530
transform 1 0 2648 0 1 2970
box -8 -3 16 105
use FILL  FILL_1267
timestamp 1745462530
transform 1 0 2640 0 1 2970
box -8 -3 16 105
use FILL  FILL_1268
timestamp 1745462530
transform 1 0 2600 0 1 2970
box -8 -3 16 105
use FILL  FILL_1269
timestamp 1745462530
transform 1 0 2560 0 1 2970
box -8 -3 16 105
use FILL  FILL_1270
timestamp 1745462530
transform 1 0 2512 0 1 2970
box -8 -3 16 105
use FILL  FILL_1271
timestamp 1745462530
transform 1 0 2504 0 1 2970
box -8 -3 16 105
use FILL  FILL_1272
timestamp 1745462530
transform 1 0 2440 0 1 2970
box -8 -3 16 105
use FILL  FILL_1273
timestamp 1745462530
transform 1 0 2432 0 1 2970
box -8 -3 16 105
use FILL  FILL_1274
timestamp 1745462530
transform 1 0 2352 0 1 2970
box -8 -3 16 105
use FILL  FILL_1275
timestamp 1745462530
transform 1 0 2248 0 1 2970
box -8 -3 16 105
use FILL  FILL_1276
timestamp 1745462530
transform 1 0 2208 0 1 2970
box -8 -3 16 105
use FILL  FILL_1277
timestamp 1745462530
transform 1 0 2200 0 1 2970
box -8 -3 16 105
use FILL  FILL_1278
timestamp 1745462530
transform 1 0 2152 0 1 2970
box -8 -3 16 105
use FILL  FILL_1279
timestamp 1745462530
transform 1 0 2104 0 1 2970
box -8 -3 16 105
use FILL  FILL_1280
timestamp 1745462530
transform 1 0 2096 0 1 2970
box -8 -3 16 105
use FILL  FILL_1281
timestamp 1745462530
transform 1 0 2048 0 1 2970
box -8 -3 16 105
use FILL  FILL_1282
timestamp 1745462530
transform 1 0 2008 0 1 2970
box -8 -3 16 105
use FILL  FILL_1283
timestamp 1745462530
transform 1 0 2000 0 1 2970
box -8 -3 16 105
use FILL  FILL_1284
timestamp 1745462530
transform 1 0 1880 0 1 2970
box -8 -3 16 105
use FILL  FILL_1285
timestamp 1745462530
transform 1 0 1816 0 1 2970
box -8 -3 16 105
use FILL  FILL_1286
timestamp 1745462530
transform 1 0 1728 0 1 2970
box -8 -3 16 105
use FILL  FILL_1287
timestamp 1745462530
transform 1 0 1688 0 1 2970
box -8 -3 16 105
use FILL  FILL_1288
timestamp 1745462530
transform 1 0 1624 0 1 2970
box -8 -3 16 105
use FILL  FILL_1289
timestamp 1745462530
transform 1 0 1616 0 1 2970
box -8 -3 16 105
use FILL  FILL_1290
timestamp 1745462530
transform 1 0 1560 0 1 2970
box -8 -3 16 105
use FILL  FILL_1291
timestamp 1745462530
transform 1 0 1552 0 1 2970
box -8 -3 16 105
use FILL  FILL_1292
timestamp 1745462530
transform 1 0 1544 0 1 2970
box -8 -3 16 105
use FILL  FILL_1293
timestamp 1745462530
transform 1 0 1496 0 1 2970
box -8 -3 16 105
use FILL  FILL_1294
timestamp 1745462530
transform 1 0 1392 0 1 2970
box -8 -3 16 105
use FILL  FILL_1295
timestamp 1745462530
transform 1 0 1384 0 1 2970
box -8 -3 16 105
use FILL  FILL_1296
timestamp 1745462530
transform 1 0 1320 0 1 2970
box -8 -3 16 105
use FILL  FILL_1297
timestamp 1745462530
transform 1 0 1312 0 1 2970
box -8 -3 16 105
use FILL  FILL_1298
timestamp 1745462530
transform 1 0 1304 0 1 2970
box -8 -3 16 105
use FILL  FILL_1299
timestamp 1745462530
transform 1 0 1248 0 1 2970
box -8 -3 16 105
use FILL  FILL_1300
timestamp 1745462530
transform 1 0 1240 0 1 2970
box -8 -3 16 105
use FILL  FILL_1301
timestamp 1745462530
transform 1 0 1168 0 1 2970
box -8 -3 16 105
use FILL  FILL_1302
timestamp 1745462530
transform 1 0 1160 0 1 2970
box -8 -3 16 105
use FILL  FILL_1303
timestamp 1745462530
transform 1 0 1096 0 1 2970
box -8 -3 16 105
use FILL  FILL_1304
timestamp 1745462530
transform 1 0 1072 0 1 2970
box -8 -3 16 105
use FILL  FILL_1305
timestamp 1745462530
transform 1 0 1064 0 1 2970
box -8 -3 16 105
use FILL  FILL_1306
timestamp 1745462530
transform 1 0 960 0 1 2970
box -8 -3 16 105
use FILL  FILL_1307
timestamp 1745462530
transform 1 0 952 0 1 2970
box -8 -3 16 105
use FILL  FILL_1308
timestamp 1745462530
transform 1 0 848 0 1 2970
box -8 -3 16 105
use FILL  FILL_1309
timestamp 1745462530
transform 1 0 840 0 1 2970
box -8 -3 16 105
use FILL  FILL_1310
timestamp 1745462530
transform 1 0 736 0 1 2970
box -8 -3 16 105
use FILL  FILL_1311
timestamp 1745462530
transform 1 0 632 0 1 2970
box -8 -3 16 105
use FILL  FILL_1312
timestamp 1745462530
transform 1 0 624 0 1 2970
box -8 -3 16 105
use FILL  FILL_1313
timestamp 1745462530
transform 1 0 560 0 1 2970
box -8 -3 16 105
use FILL  FILL_1314
timestamp 1745462530
transform 1 0 520 0 1 2970
box -8 -3 16 105
use FILL  FILL_1315
timestamp 1745462530
transform 1 0 456 0 1 2970
box -8 -3 16 105
use FILL  FILL_1316
timestamp 1745462530
transform 1 0 448 0 1 2970
box -8 -3 16 105
use FILL  FILL_1317
timestamp 1745462530
transform 1 0 352 0 1 2970
box -8 -3 16 105
use FILL  FILL_1318
timestamp 1745462530
transform 1 0 344 0 1 2970
box -8 -3 16 105
use FILL  FILL_1319
timestamp 1745462530
transform 1 0 304 0 1 2970
box -8 -3 16 105
use FILL  FILL_1320
timestamp 1745462530
transform 1 0 296 0 1 2970
box -8 -3 16 105
use FILL  FILL_1321
timestamp 1745462530
transform 1 0 232 0 1 2970
box -8 -3 16 105
use FILL  FILL_1322
timestamp 1745462530
transform 1 0 144 0 1 2970
box -8 -3 16 105
use FILL  FILL_1323
timestamp 1745462530
transform 1 0 136 0 1 2970
box -8 -3 16 105
use FILL  FILL_1324
timestamp 1745462530
transform 1 0 72 0 1 2970
box -8 -3 16 105
use FILL  FILL_1325
timestamp 1745462530
transform 1 0 4272 0 -1 2970
box -8 -3 16 105
use FILL  FILL_1326
timestamp 1745462530
transform 1 0 3944 0 -1 2970
box -8 -3 16 105
use FILL  FILL_1327
timestamp 1745462530
transform 1 0 3880 0 -1 2970
box -8 -3 16 105
use FILL  FILL_1328
timestamp 1745462530
transform 1 0 3776 0 -1 2970
box -8 -3 16 105
use FILL  FILL_1329
timestamp 1745462530
transform 1 0 3712 0 -1 2970
box -8 -3 16 105
use FILL  FILL_1330
timestamp 1745462530
transform 1 0 3688 0 -1 2970
box -8 -3 16 105
use FILL  FILL_1331
timestamp 1745462530
transform 1 0 3584 0 -1 2970
box -8 -3 16 105
use FILL  FILL_1332
timestamp 1745462530
transform 1 0 3576 0 -1 2970
box -8 -3 16 105
use FILL  FILL_1333
timestamp 1745462530
transform 1 0 3512 0 -1 2970
box -8 -3 16 105
use FILL  FILL_1334
timestamp 1745462530
transform 1 0 3352 0 -1 2970
box -8 -3 16 105
use FILL  FILL_1335
timestamp 1745462530
transform 1 0 3344 0 -1 2970
box -8 -3 16 105
use FILL  FILL_1336
timestamp 1745462530
transform 1 0 3336 0 -1 2970
box -8 -3 16 105
use FILL  FILL_1337
timestamp 1745462530
transform 1 0 3272 0 -1 2970
box -8 -3 16 105
use FILL  FILL_1338
timestamp 1745462530
transform 1 0 3208 0 -1 2970
box -8 -3 16 105
use FILL  FILL_1339
timestamp 1745462530
transform 1 0 3144 0 -1 2970
box -8 -3 16 105
use FILL  FILL_1340
timestamp 1745462530
transform 1 0 3040 0 -1 2970
box -8 -3 16 105
use FILL  FILL_1341
timestamp 1745462530
transform 1 0 3032 0 -1 2970
box -8 -3 16 105
use FILL  FILL_1342
timestamp 1745462530
transform 1 0 2968 0 -1 2970
box -8 -3 16 105
use FILL  FILL_1343
timestamp 1745462530
transform 1 0 2864 0 -1 2970
box -8 -3 16 105
use FILL  FILL_1344
timestamp 1745462530
transform 1 0 2856 0 -1 2970
box -8 -3 16 105
use FILL  FILL_1345
timestamp 1745462530
transform 1 0 2752 0 -1 2970
box -8 -3 16 105
use FILL  FILL_1346
timestamp 1745462530
transform 1 0 2744 0 -1 2970
box -8 -3 16 105
use FILL  FILL_1347
timestamp 1745462530
transform 1 0 2640 0 -1 2970
box -8 -3 16 105
use FILL  FILL_1348
timestamp 1745462530
transform 1 0 2632 0 -1 2970
box -8 -3 16 105
use FILL  FILL_1349
timestamp 1745462530
transform 1 0 2592 0 -1 2970
box -8 -3 16 105
use FILL  FILL_1350
timestamp 1745462530
transform 1 0 2488 0 -1 2970
box -8 -3 16 105
use FILL  FILL_1351
timestamp 1745462530
transform 1 0 2480 0 -1 2970
box -8 -3 16 105
use FILL  FILL_1352
timestamp 1745462530
transform 1 0 2376 0 -1 2970
box -8 -3 16 105
use FILL  FILL_1353
timestamp 1745462530
transform 1 0 2368 0 -1 2970
box -8 -3 16 105
use FILL  FILL_1354
timestamp 1745462530
transform 1 0 2264 0 -1 2970
box -8 -3 16 105
use FILL  FILL_1355
timestamp 1745462530
transform 1 0 2256 0 -1 2970
box -8 -3 16 105
use FILL  FILL_1356
timestamp 1745462530
transform 1 0 2216 0 -1 2970
box -8 -3 16 105
use FILL  FILL_1357
timestamp 1745462530
transform 1 0 2208 0 -1 2970
box -8 -3 16 105
use FILL  FILL_1358
timestamp 1745462530
transform 1 0 2200 0 -1 2970
box -8 -3 16 105
use FILL  FILL_1359
timestamp 1745462530
transform 1 0 2152 0 -1 2970
box -8 -3 16 105
use FILL  FILL_1360
timestamp 1745462530
transform 1 0 2144 0 -1 2970
box -8 -3 16 105
use FILL  FILL_1361
timestamp 1745462530
transform 1 0 2136 0 -1 2970
box -8 -3 16 105
use FILL  FILL_1362
timestamp 1745462530
transform 1 0 2088 0 -1 2970
box -8 -3 16 105
use FILL  FILL_1363
timestamp 1745462530
transform 1 0 2080 0 -1 2970
box -8 -3 16 105
use FILL  FILL_1364
timestamp 1745462530
transform 1 0 2072 0 -1 2970
box -8 -3 16 105
use FILL  FILL_1365
timestamp 1745462530
transform 1 0 2024 0 -1 2970
box -8 -3 16 105
use FILL  FILL_1366
timestamp 1745462530
transform 1 0 2016 0 -1 2970
box -8 -3 16 105
use FILL  FILL_1367
timestamp 1745462530
transform 1 0 1968 0 -1 2970
box -8 -3 16 105
use FILL  FILL_1368
timestamp 1745462530
transform 1 0 1960 0 -1 2970
box -8 -3 16 105
use FILL  FILL_1369
timestamp 1745462530
transform 1 0 1912 0 -1 2970
box -8 -3 16 105
use FILL  FILL_1370
timestamp 1745462530
transform 1 0 1904 0 -1 2970
box -8 -3 16 105
use FILL  FILL_1371
timestamp 1745462530
transform 1 0 1800 0 -1 2970
box -8 -3 16 105
use FILL  FILL_1372
timestamp 1745462530
transform 1 0 1792 0 -1 2970
box -8 -3 16 105
use FILL  FILL_1373
timestamp 1745462530
transform 1 0 1688 0 -1 2970
box -8 -3 16 105
use FILL  FILL_1374
timestamp 1745462530
transform 1 0 1640 0 -1 2970
box -8 -3 16 105
use FILL  FILL_1375
timestamp 1745462530
transform 1 0 1632 0 -1 2970
box -8 -3 16 105
use FILL  FILL_1376
timestamp 1745462530
transform 1 0 1528 0 -1 2970
box -8 -3 16 105
use FILL  FILL_1377
timestamp 1745462530
transform 1 0 1480 0 -1 2970
box -8 -3 16 105
use FILL  FILL_1378
timestamp 1745462530
transform 1 0 1472 0 -1 2970
box -8 -3 16 105
use FILL  FILL_1379
timestamp 1745462530
transform 1 0 1424 0 -1 2970
box -8 -3 16 105
use FILL  FILL_1380
timestamp 1745462530
transform 1 0 1320 0 -1 2970
box -8 -3 16 105
use FILL  FILL_1381
timestamp 1745462530
transform 1 0 1312 0 -1 2970
box -8 -3 16 105
use FILL  FILL_1382
timestamp 1745462530
transform 1 0 1208 0 -1 2970
box -8 -3 16 105
use FILL  FILL_1383
timestamp 1745462530
transform 1 0 1104 0 -1 2970
box -8 -3 16 105
use FILL  FILL_1384
timestamp 1745462530
transform 1 0 1096 0 -1 2970
box -8 -3 16 105
use FILL  FILL_1385
timestamp 1745462530
transform 1 0 992 0 -1 2970
box -8 -3 16 105
use FILL  FILL_1386
timestamp 1745462530
transform 1 0 984 0 -1 2970
box -8 -3 16 105
use FILL  FILL_1387
timestamp 1745462530
transform 1 0 936 0 -1 2970
box -8 -3 16 105
use FILL  FILL_1388
timestamp 1745462530
transform 1 0 888 0 -1 2970
box -8 -3 16 105
use FILL  FILL_1389
timestamp 1745462530
transform 1 0 880 0 -1 2970
box -8 -3 16 105
use FILL  FILL_1390
timestamp 1745462530
transform 1 0 816 0 -1 2970
box -8 -3 16 105
use FILL  FILL_1391
timestamp 1745462530
transform 1 0 808 0 -1 2970
box -8 -3 16 105
use FILL  FILL_1392
timestamp 1745462530
transform 1 0 784 0 -1 2970
box -8 -3 16 105
use FILL  FILL_1393
timestamp 1745462530
transform 1 0 736 0 -1 2970
box -8 -3 16 105
use FILL  FILL_1394
timestamp 1745462530
transform 1 0 728 0 -1 2970
box -8 -3 16 105
use FILL  FILL_1395
timestamp 1745462530
transform 1 0 664 0 -1 2970
box -8 -3 16 105
use FILL  FILL_1396
timestamp 1745462530
transform 1 0 656 0 -1 2970
box -8 -3 16 105
use FILL  FILL_1397
timestamp 1745462530
transform 1 0 648 0 -1 2970
box -8 -3 16 105
use FILL  FILL_1398
timestamp 1745462530
transform 1 0 544 0 -1 2970
box -8 -3 16 105
use FILL  FILL_1399
timestamp 1745462530
transform 1 0 536 0 -1 2970
box -8 -3 16 105
use FILL  FILL_1400
timestamp 1745462530
transform 1 0 528 0 -1 2970
box -8 -3 16 105
use FILL  FILL_1401
timestamp 1745462530
transform 1 0 424 0 -1 2970
box -8 -3 16 105
use FILL  FILL_1402
timestamp 1745462530
transform 1 0 416 0 -1 2970
box -8 -3 16 105
use FILL  FILL_1403
timestamp 1745462530
transform 1 0 312 0 -1 2970
box -8 -3 16 105
use FILL  FILL_1404
timestamp 1745462530
transform 1 0 304 0 -1 2970
box -8 -3 16 105
use FILL  FILL_1405
timestamp 1745462530
transform 1 0 280 0 -1 2970
box -8 -3 16 105
use FILL  FILL_1406
timestamp 1745462530
transform 1 0 272 0 -1 2970
box -8 -3 16 105
use FILL  FILL_1407
timestamp 1745462530
transform 1 0 168 0 -1 2970
box -8 -3 16 105
use FILL  FILL_1408
timestamp 1745462530
transform 1 0 160 0 -1 2970
box -8 -3 16 105
use FILL  FILL_1409
timestamp 1745462530
transform 1 0 152 0 -1 2970
box -8 -3 16 105
use FILL  FILL_1410
timestamp 1745462530
transform 1 0 144 0 -1 2970
box -8 -3 16 105
use FILL  FILL_1411
timestamp 1745462530
transform 1 0 136 0 -1 2970
box -8 -3 16 105
use FILL  FILL_1412
timestamp 1745462530
transform 1 0 128 0 -1 2970
box -8 -3 16 105
use FILL  FILL_1413
timestamp 1745462530
transform 1 0 120 0 -1 2970
box -8 -3 16 105
use FILL  FILL_1414
timestamp 1745462530
transform 1 0 112 0 -1 2970
box -8 -3 16 105
use FILL  FILL_1415
timestamp 1745462530
transform 1 0 104 0 -1 2970
box -8 -3 16 105
use FILL  FILL_1416
timestamp 1745462530
transform 1 0 96 0 -1 2970
box -8 -3 16 105
use FILL  FILL_1417
timestamp 1745462530
transform 1 0 88 0 -1 2970
box -8 -3 16 105
use FILL  FILL_1418
timestamp 1745462530
transform 1 0 80 0 -1 2970
box -8 -3 16 105
use FILL  FILL_1419
timestamp 1745462530
transform 1 0 72 0 -1 2970
box -8 -3 16 105
use FILL  FILL_1420
timestamp 1745462530
transform 1 0 4272 0 1 2770
box -8 -3 16 105
use FILL  FILL_1421
timestamp 1745462530
transform 1 0 4128 0 1 2770
box -8 -3 16 105
use FILL  FILL_1422
timestamp 1745462530
transform 1 0 4064 0 1 2770
box -8 -3 16 105
use FILL  FILL_1423
timestamp 1745462530
transform 1 0 4000 0 1 2770
box -8 -3 16 105
use FILL  FILL_1424
timestamp 1745462530
transform 1 0 3992 0 1 2770
box -8 -3 16 105
use FILL  FILL_1425
timestamp 1745462530
transform 1 0 3888 0 1 2770
box -8 -3 16 105
use FILL  FILL_1426
timestamp 1745462530
transform 1 0 3840 0 1 2770
box -8 -3 16 105
use FILL  FILL_1427
timestamp 1745462530
transform 1 0 3776 0 1 2770
box -8 -3 16 105
use FILL  FILL_1428
timestamp 1745462530
transform 1 0 3768 0 1 2770
box -8 -3 16 105
use FILL  FILL_1429
timestamp 1745462530
transform 1 0 3664 0 1 2770
box -8 -3 16 105
use FILL  FILL_1430
timestamp 1745462530
transform 1 0 3656 0 1 2770
box -8 -3 16 105
use FILL  FILL_1431
timestamp 1745462530
transform 1 0 3592 0 1 2770
box -8 -3 16 105
use FILL  FILL_1432
timestamp 1745462530
transform 1 0 3584 0 1 2770
box -8 -3 16 105
use FILL  FILL_1433
timestamp 1745462530
transform 1 0 3536 0 1 2770
box -8 -3 16 105
use FILL  FILL_1434
timestamp 1745462530
transform 1 0 3432 0 1 2770
box -8 -3 16 105
use FILL  FILL_1435
timestamp 1745462530
transform 1 0 3424 0 1 2770
box -8 -3 16 105
use FILL  FILL_1436
timestamp 1745462530
transform 1 0 3360 0 1 2770
box -8 -3 16 105
use FILL  FILL_1437
timestamp 1745462530
transform 1 0 3352 0 1 2770
box -8 -3 16 105
use FILL  FILL_1438
timestamp 1745462530
transform 1 0 3304 0 1 2770
box -8 -3 16 105
use FILL  FILL_1439
timestamp 1745462530
transform 1 0 3296 0 1 2770
box -8 -3 16 105
use FILL  FILL_1440
timestamp 1745462530
transform 1 0 3232 0 1 2770
box -8 -3 16 105
use FILL  FILL_1441
timestamp 1745462530
transform 1 0 3224 0 1 2770
box -8 -3 16 105
use FILL  FILL_1442
timestamp 1745462530
transform 1 0 3160 0 1 2770
box -8 -3 16 105
use FILL  FILL_1443
timestamp 1745462530
transform 1 0 3152 0 1 2770
box -8 -3 16 105
use FILL  FILL_1444
timestamp 1745462530
transform 1 0 3048 0 1 2770
box -8 -3 16 105
use FILL  FILL_1445
timestamp 1745462530
transform 1 0 3040 0 1 2770
box -8 -3 16 105
use FILL  FILL_1446
timestamp 1745462530
transform 1 0 2992 0 1 2770
box -8 -3 16 105
use FILL  FILL_1447
timestamp 1745462530
transform 1 0 2984 0 1 2770
box -8 -3 16 105
use FILL  FILL_1448
timestamp 1745462530
transform 1 0 2944 0 1 2770
box -8 -3 16 105
use FILL  FILL_1449
timestamp 1745462530
transform 1 0 2936 0 1 2770
box -8 -3 16 105
use FILL  FILL_1450
timestamp 1745462530
transform 1 0 2928 0 1 2770
box -8 -3 16 105
use FILL  FILL_1451
timestamp 1745462530
transform 1 0 2824 0 1 2770
box -8 -3 16 105
use FILL  FILL_1452
timestamp 1745462530
transform 1 0 2816 0 1 2770
box -8 -3 16 105
use FILL  FILL_1453
timestamp 1745462530
transform 1 0 2808 0 1 2770
box -8 -3 16 105
use FILL  FILL_1454
timestamp 1745462530
transform 1 0 2800 0 1 2770
box -8 -3 16 105
use FILL  FILL_1455
timestamp 1745462530
transform 1 0 2736 0 1 2770
box -8 -3 16 105
use FILL  FILL_1456
timestamp 1745462530
transform 1 0 2728 0 1 2770
box -8 -3 16 105
use FILL  FILL_1457
timestamp 1745462530
transform 1 0 2720 0 1 2770
box -8 -3 16 105
use FILL  FILL_1458
timestamp 1745462530
transform 1 0 2672 0 1 2770
box -8 -3 16 105
use FILL  FILL_1459
timestamp 1745462530
transform 1 0 2648 0 1 2770
box -8 -3 16 105
use FILL  FILL_1460
timestamp 1745462530
transform 1 0 2640 0 1 2770
box -8 -3 16 105
use FILL  FILL_1461
timestamp 1745462530
transform 1 0 2592 0 1 2770
box -8 -3 16 105
use FILL  FILL_1462
timestamp 1745462530
transform 1 0 2584 0 1 2770
box -8 -3 16 105
use FILL  FILL_1463
timestamp 1745462530
transform 1 0 2544 0 1 2770
box -8 -3 16 105
use FILL  FILL_1464
timestamp 1745462530
transform 1 0 2536 0 1 2770
box -8 -3 16 105
use FILL  FILL_1465
timestamp 1745462530
transform 1 0 2528 0 1 2770
box -8 -3 16 105
use FILL  FILL_1466
timestamp 1745462530
transform 1 0 2480 0 1 2770
box -8 -3 16 105
use FILL  FILL_1467
timestamp 1745462530
transform 1 0 2456 0 1 2770
box -8 -3 16 105
use FILL  FILL_1468
timestamp 1745462530
transform 1 0 2448 0 1 2770
box -8 -3 16 105
use FILL  FILL_1469
timestamp 1745462530
transform 1 0 2344 0 1 2770
box -8 -3 16 105
use FILL  FILL_1470
timestamp 1745462530
transform 1 0 2336 0 1 2770
box -8 -3 16 105
use FILL  FILL_1471
timestamp 1745462530
transform 1 0 2296 0 1 2770
box -8 -3 16 105
use FILL  FILL_1472
timestamp 1745462530
transform 1 0 2288 0 1 2770
box -8 -3 16 105
use FILL  FILL_1473
timestamp 1745462530
transform 1 0 2280 0 1 2770
box -8 -3 16 105
use FILL  FILL_1474
timestamp 1745462530
transform 1 0 2176 0 1 2770
box -8 -3 16 105
use FILL  FILL_1475
timestamp 1745462530
transform 1 0 2136 0 1 2770
box -8 -3 16 105
use FILL  FILL_1476
timestamp 1745462530
transform 1 0 2128 0 1 2770
box -8 -3 16 105
use FILL  FILL_1477
timestamp 1745462530
transform 1 0 2088 0 1 2770
box -8 -3 16 105
use FILL  FILL_1478
timestamp 1745462530
transform 1 0 2080 0 1 2770
box -8 -3 16 105
use FILL  FILL_1479
timestamp 1745462530
transform 1 0 2040 0 1 2770
box -8 -3 16 105
use FILL  FILL_1480
timestamp 1745462530
transform 1 0 2032 0 1 2770
box -8 -3 16 105
use FILL  FILL_1481
timestamp 1745462530
transform 1 0 2024 0 1 2770
box -8 -3 16 105
use FILL  FILL_1482
timestamp 1745462530
transform 1 0 1920 0 1 2770
box -8 -3 16 105
use FILL  FILL_1483
timestamp 1745462530
transform 1 0 1912 0 1 2770
box -8 -3 16 105
use FILL  FILL_1484
timestamp 1745462530
transform 1 0 1864 0 1 2770
box -8 -3 16 105
use FILL  FILL_1485
timestamp 1745462530
transform 1 0 1856 0 1 2770
box -8 -3 16 105
use FILL  FILL_1486
timestamp 1745462530
transform 1 0 1792 0 1 2770
box -8 -3 16 105
use FILL  FILL_1487
timestamp 1745462530
transform 1 0 1784 0 1 2770
box -8 -3 16 105
use FILL  FILL_1488
timestamp 1745462530
transform 1 0 1776 0 1 2770
box -8 -3 16 105
use FILL  FILL_1489
timestamp 1745462530
transform 1 0 1728 0 1 2770
box -8 -3 16 105
use FILL  FILL_1490
timestamp 1745462530
transform 1 0 1704 0 1 2770
box -8 -3 16 105
use FILL  FILL_1491
timestamp 1745462530
transform 1 0 1696 0 1 2770
box -8 -3 16 105
use FILL  FILL_1492
timestamp 1745462530
transform 1 0 1632 0 1 2770
box -8 -3 16 105
use FILL  FILL_1493
timestamp 1745462530
transform 1 0 1624 0 1 2770
box -8 -3 16 105
use FILL  FILL_1494
timestamp 1745462530
transform 1 0 1576 0 1 2770
box -8 -3 16 105
use FILL  FILL_1495
timestamp 1745462530
transform 1 0 1552 0 1 2770
box -8 -3 16 105
use FILL  FILL_1496
timestamp 1745462530
transform 1 0 1504 0 1 2770
box -8 -3 16 105
use FILL  FILL_1497
timestamp 1745462530
transform 1 0 1496 0 1 2770
box -8 -3 16 105
use FILL  FILL_1498
timestamp 1745462530
transform 1 0 1456 0 1 2770
box -8 -3 16 105
use FILL  FILL_1499
timestamp 1745462530
transform 1 0 1408 0 1 2770
box -8 -3 16 105
use FILL  FILL_1500
timestamp 1745462530
transform 1 0 1400 0 1 2770
box -8 -3 16 105
use FILL  FILL_1501
timestamp 1745462530
transform 1 0 1392 0 1 2770
box -8 -3 16 105
use FILL  FILL_1502
timestamp 1745462530
transform 1 0 1328 0 1 2770
box -8 -3 16 105
use FILL  FILL_1503
timestamp 1745462530
transform 1 0 1280 0 1 2770
box -8 -3 16 105
use FILL  FILL_1504
timestamp 1745462530
transform 1 0 1272 0 1 2770
box -8 -3 16 105
use FILL  FILL_1505
timestamp 1745462530
transform 1 0 1224 0 1 2770
box -8 -3 16 105
use FILL  FILL_1506
timestamp 1745462530
transform 1 0 1216 0 1 2770
box -8 -3 16 105
use FILL  FILL_1507
timestamp 1745462530
transform 1 0 1168 0 1 2770
box -8 -3 16 105
use FILL  FILL_1508
timestamp 1745462530
transform 1 0 1144 0 1 2770
box -8 -3 16 105
use FILL  FILL_1509
timestamp 1745462530
transform 1 0 1136 0 1 2770
box -8 -3 16 105
use FILL  FILL_1510
timestamp 1745462530
transform 1 0 1032 0 1 2770
box -8 -3 16 105
use FILL  FILL_1511
timestamp 1745462530
transform 1 0 992 0 1 2770
box -8 -3 16 105
use FILL  FILL_1512
timestamp 1745462530
transform 1 0 984 0 1 2770
box -8 -3 16 105
use FILL  FILL_1513
timestamp 1745462530
transform 1 0 936 0 1 2770
box -8 -3 16 105
use FILL  FILL_1514
timestamp 1745462530
transform 1 0 896 0 1 2770
box -8 -3 16 105
use FILL  FILL_1515
timestamp 1745462530
transform 1 0 848 0 1 2770
box -8 -3 16 105
use FILL  FILL_1516
timestamp 1745462530
transform 1 0 816 0 1 2770
box -8 -3 16 105
use FILL  FILL_1517
timestamp 1745462530
transform 1 0 768 0 1 2770
box -8 -3 16 105
use FILL  FILL_1518
timestamp 1745462530
transform 1 0 720 0 1 2770
box -8 -3 16 105
use FILL  FILL_1519
timestamp 1745462530
transform 1 0 688 0 1 2770
box -8 -3 16 105
use FILL  FILL_1520
timestamp 1745462530
transform 1 0 640 0 1 2770
box -8 -3 16 105
use FILL  FILL_1521
timestamp 1745462530
transform 1 0 616 0 1 2770
box -8 -3 16 105
use FILL  FILL_1522
timestamp 1745462530
transform 1 0 568 0 1 2770
box -8 -3 16 105
use FILL  FILL_1523
timestamp 1745462530
transform 1 0 560 0 1 2770
box -8 -3 16 105
use FILL  FILL_1524
timestamp 1745462530
transform 1 0 496 0 1 2770
box -8 -3 16 105
use FILL  FILL_1525
timestamp 1745462530
transform 1 0 488 0 1 2770
box -8 -3 16 105
use FILL  FILL_1526
timestamp 1745462530
transform 1 0 424 0 1 2770
box -8 -3 16 105
use FILL  FILL_1527
timestamp 1745462530
transform 1 0 416 0 1 2770
box -8 -3 16 105
use FILL  FILL_1528
timestamp 1745462530
transform 1 0 352 0 1 2770
box -8 -3 16 105
use FILL  FILL_1529
timestamp 1745462530
transform 1 0 328 0 1 2770
box -8 -3 16 105
use FILL  FILL_1530
timestamp 1745462530
transform 1 0 320 0 1 2770
box -8 -3 16 105
use FILL  FILL_1531
timestamp 1745462530
transform 1 0 256 0 1 2770
box -8 -3 16 105
use FILL  FILL_1532
timestamp 1745462530
transform 1 0 248 0 1 2770
box -8 -3 16 105
use FILL  FILL_1533
timestamp 1745462530
transform 1 0 200 0 1 2770
box -8 -3 16 105
use FILL  FILL_1534
timestamp 1745462530
transform 1 0 176 0 1 2770
box -8 -3 16 105
use FILL  FILL_1535
timestamp 1745462530
transform 1 0 72 0 1 2770
box -8 -3 16 105
use FILL  FILL_1536
timestamp 1745462530
transform 1 0 4368 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1537
timestamp 1745462530
transform 1 0 4360 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1538
timestamp 1745462530
transform 1 0 4352 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1539
timestamp 1745462530
transform 1 0 4344 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1540
timestamp 1745462530
transform 1 0 4336 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1541
timestamp 1745462530
transform 1 0 4328 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1542
timestamp 1745462530
transform 1 0 4224 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1543
timestamp 1745462530
transform 1 0 4216 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1544
timestamp 1745462530
transform 1 0 4152 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1545
timestamp 1745462530
transform 1 0 4144 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1546
timestamp 1745462530
transform 1 0 4080 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1547
timestamp 1745462530
transform 1 0 4032 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1548
timestamp 1745462530
transform 1 0 4024 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1549
timestamp 1745462530
transform 1 0 4016 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1550
timestamp 1745462530
transform 1 0 3976 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1551
timestamp 1745462530
transform 1 0 3968 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1552
timestamp 1745462530
transform 1 0 3920 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1553
timestamp 1745462530
transform 1 0 3912 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1554
timestamp 1745462530
transform 1 0 3904 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1555
timestamp 1745462530
transform 1 0 3896 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1556
timestamp 1745462530
transform 1 0 3848 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1557
timestamp 1745462530
transform 1 0 3840 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1558
timestamp 1745462530
transform 1 0 3816 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1559
timestamp 1745462530
transform 1 0 3808 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1560
timestamp 1745462530
transform 1 0 3800 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1561
timestamp 1745462530
transform 1 0 3752 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1562
timestamp 1745462530
transform 1 0 3728 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1563
timestamp 1745462530
transform 1 0 3720 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1564
timestamp 1745462530
transform 1 0 3712 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1565
timestamp 1745462530
transform 1 0 3704 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1566
timestamp 1745462530
transform 1 0 3656 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1567
timestamp 1745462530
transform 1 0 3648 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1568
timestamp 1745462530
transform 1 0 3624 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1569
timestamp 1745462530
transform 1 0 3616 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1570
timestamp 1745462530
transform 1 0 3568 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1571
timestamp 1745462530
transform 1 0 3560 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1572
timestamp 1745462530
transform 1 0 3552 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1573
timestamp 1745462530
transform 1 0 3504 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1574
timestamp 1745462530
transform 1 0 3496 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1575
timestamp 1745462530
transform 1 0 3472 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1576
timestamp 1745462530
transform 1 0 3424 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1577
timestamp 1745462530
transform 1 0 3416 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1578
timestamp 1745462530
transform 1 0 3408 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1579
timestamp 1745462530
transform 1 0 3360 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1580
timestamp 1745462530
transform 1 0 3352 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1581
timestamp 1745462530
transform 1 0 3312 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1582
timestamp 1745462530
transform 1 0 3304 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1583
timestamp 1745462530
transform 1 0 3256 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1584
timestamp 1745462530
transform 1 0 3248 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1585
timestamp 1745462530
transform 1 0 3144 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1586
timestamp 1745462530
transform 1 0 3136 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1587
timestamp 1745462530
transform 1 0 3096 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1588
timestamp 1745462530
transform 1 0 3056 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1589
timestamp 1745462530
transform 1 0 3048 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1590
timestamp 1745462530
transform 1 0 3008 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1591
timestamp 1745462530
transform 1 0 2976 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1592
timestamp 1745462530
transform 1 0 2872 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1593
timestamp 1745462530
transform 1 0 2848 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1594
timestamp 1745462530
transform 1 0 2840 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1595
timestamp 1745462530
transform 1 0 2664 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1596
timestamp 1745462530
transform 1 0 2656 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1597
timestamp 1745462530
transform 1 0 2608 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1598
timestamp 1745462530
transform 1 0 2504 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1599
timestamp 1745462530
transform 1 0 2424 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1600
timestamp 1745462530
transform 1 0 2384 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1601
timestamp 1745462530
transform 1 0 2376 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1602
timestamp 1745462530
transform 1 0 2320 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1603
timestamp 1745462530
transform 1 0 2288 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1604
timestamp 1745462530
transform 1 0 2248 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1605
timestamp 1745462530
transform 1 0 2184 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1606
timestamp 1745462530
transform 1 0 2080 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1607
timestamp 1745462530
transform 1 0 1960 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1608
timestamp 1745462530
transform 1 0 1856 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1609
timestamp 1745462530
transform 1 0 1808 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1610
timestamp 1745462530
transform 1 0 1664 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1611
timestamp 1745462530
transform 1 0 1608 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1612
timestamp 1745462530
transform 1 0 1504 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1613
timestamp 1745462530
transform 1 0 1464 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1614
timestamp 1745462530
transform 1 0 1360 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1615
timestamp 1745462530
transform 1 0 1320 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1616
timestamp 1745462530
transform 1 0 1256 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1617
timestamp 1745462530
transform 1 0 1064 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1618
timestamp 1745462530
transform 1 0 824 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1619
timestamp 1745462530
transform 1 0 736 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1620
timestamp 1745462530
transform 1 0 664 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1621
timestamp 1745462530
transform 1 0 560 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1622
timestamp 1745462530
transform 1 0 456 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1623
timestamp 1745462530
transform 1 0 392 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1624
timestamp 1745462530
transform 1 0 248 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1625
timestamp 1745462530
transform 1 0 168 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1626
timestamp 1745462530
transform 1 0 4368 0 1 2570
box -8 -3 16 105
use FILL  FILL_1627
timestamp 1745462530
transform 1 0 4360 0 1 2570
box -8 -3 16 105
use FILL  FILL_1628
timestamp 1745462530
transform 1 0 4352 0 1 2570
box -8 -3 16 105
use FILL  FILL_1629
timestamp 1745462530
transform 1 0 4344 0 1 2570
box -8 -3 16 105
use FILL  FILL_1630
timestamp 1745462530
transform 1 0 4336 0 1 2570
box -8 -3 16 105
use FILL  FILL_1631
timestamp 1745462530
transform 1 0 4232 0 1 2570
box -8 -3 16 105
use FILL  FILL_1632
timestamp 1745462530
transform 1 0 4224 0 1 2570
box -8 -3 16 105
use FILL  FILL_1633
timestamp 1745462530
transform 1 0 4160 0 1 2570
box -8 -3 16 105
use FILL  FILL_1634
timestamp 1745462530
transform 1 0 4152 0 1 2570
box -8 -3 16 105
use FILL  FILL_1635
timestamp 1745462530
transform 1 0 4104 0 1 2570
box -8 -3 16 105
use FILL  FILL_1636
timestamp 1745462530
transform 1 0 4064 0 1 2570
box -8 -3 16 105
use FILL  FILL_1637
timestamp 1745462530
transform 1 0 4024 0 1 2570
box -8 -3 16 105
use FILL  FILL_1638
timestamp 1745462530
transform 1 0 4016 0 1 2570
box -8 -3 16 105
use FILL  FILL_1639
timestamp 1745462530
transform 1 0 3968 0 1 2570
box -8 -3 16 105
use FILL  FILL_1640
timestamp 1745462530
transform 1 0 3960 0 1 2570
box -8 -3 16 105
use FILL  FILL_1641
timestamp 1745462530
transform 1 0 3856 0 1 2570
box -8 -3 16 105
use FILL  FILL_1642
timestamp 1745462530
transform 1 0 3816 0 1 2570
box -8 -3 16 105
use FILL  FILL_1643
timestamp 1745462530
transform 1 0 3776 0 1 2570
box -8 -3 16 105
use FILL  FILL_1644
timestamp 1745462530
transform 1 0 3728 0 1 2570
box -8 -3 16 105
use FILL  FILL_1645
timestamp 1745462530
transform 1 0 3720 0 1 2570
box -8 -3 16 105
use FILL  FILL_1646
timestamp 1745462530
transform 1 0 3616 0 1 2570
box -8 -3 16 105
use FILL  FILL_1647
timestamp 1745462530
transform 1 0 3608 0 1 2570
box -8 -3 16 105
use FILL  FILL_1648
timestamp 1745462530
transform 1 0 3560 0 1 2570
box -8 -3 16 105
use FILL  FILL_1649
timestamp 1745462530
transform 1 0 3552 0 1 2570
box -8 -3 16 105
use FILL  FILL_1650
timestamp 1745462530
transform 1 0 3512 0 1 2570
box -8 -3 16 105
use FILL  FILL_1651
timestamp 1745462530
transform 1 0 3504 0 1 2570
box -8 -3 16 105
use FILL  FILL_1652
timestamp 1745462530
transform 1 0 3464 0 1 2570
box -8 -3 16 105
use FILL  FILL_1653
timestamp 1745462530
transform 1 0 3456 0 1 2570
box -8 -3 16 105
use FILL  FILL_1654
timestamp 1745462530
transform 1 0 3416 0 1 2570
box -8 -3 16 105
use FILL  FILL_1655
timestamp 1745462530
transform 1 0 3408 0 1 2570
box -8 -3 16 105
use FILL  FILL_1656
timestamp 1745462530
transform 1 0 3400 0 1 2570
box -8 -3 16 105
use FILL  FILL_1657
timestamp 1745462530
transform 1 0 3368 0 1 2570
box -8 -3 16 105
use FILL  FILL_1658
timestamp 1745462530
transform 1 0 3360 0 1 2570
box -8 -3 16 105
use FILL  FILL_1659
timestamp 1745462530
transform 1 0 3320 0 1 2570
box -8 -3 16 105
use FILL  FILL_1660
timestamp 1745462530
transform 1 0 3312 0 1 2570
box -8 -3 16 105
use FILL  FILL_1661
timestamp 1745462530
transform 1 0 3304 0 1 2570
box -8 -3 16 105
use FILL  FILL_1662
timestamp 1745462530
transform 1 0 3256 0 1 2570
box -8 -3 16 105
use FILL  FILL_1663
timestamp 1745462530
transform 1 0 3248 0 1 2570
box -8 -3 16 105
use FILL  FILL_1664
timestamp 1745462530
transform 1 0 3200 0 1 2570
box -8 -3 16 105
use FILL  FILL_1665
timestamp 1745462530
transform 1 0 3176 0 1 2570
box -8 -3 16 105
use FILL  FILL_1666
timestamp 1745462530
transform 1 0 3168 0 1 2570
box -8 -3 16 105
use FILL  FILL_1667
timestamp 1745462530
transform 1 0 3128 0 1 2570
box -8 -3 16 105
use FILL  FILL_1668
timestamp 1745462530
transform 1 0 3080 0 1 2570
box -8 -3 16 105
use FILL  FILL_1669
timestamp 1745462530
transform 1 0 3072 0 1 2570
box -8 -3 16 105
use FILL  FILL_1670
timestamp 1745462530
transform 1 0 3064 0 1 2570
box -8 -3 16 105
use FILL  FILL_1671
timestamp 1745462530
transform 1 0 3024 0 1 2570
box -8 -3 16 105
use FILL  FILL_1672
timestamp 1745462530
transform 1 0 2984 0 1 2570
box -8 -3 16 105
use FILL  FILL_1673
timestamp 1745462530
transform 1 0 2976 0 1 2570
box -8 -3 16 105
use FILL  FILL_1674
timestamp 1745462530
transform 1 0 2968 0 1 2570
box -8 -3 16 105
use FILL  FILL_1675
timestamp 1745462530
transform 1 0 2920 0 1 2570
box -8 -3 16 105
use FILL  FILL_1676
timestamp 1745462530
transform 1 0 2912 0 1 2570
box -8 -3 16 105
use FILL  FILL_1677
timestamp 1745462530
transform 1 0 2904 0 1 2570
box -8 -3 16 105
use FILL  FILL_1678
timestamp 1745462530
transform 1 0 2856 0 1 2570
box -8 -3 16 105
use FILL  FILL_1679
timestamp 1745462530
transform 1 0 2848 0 1 2570
box -8 -3 16 105
use FILL  FILL_1680
timestamp 1745462530
transform 1 0 2824 0 1 2570
box -8 -3 16 105
use FILL  FILL_1681
timestamp 1745462530
transform 1 0 2720 0 1 2570
box -8 -3 16 105
use FILL  FILL_1682
timestamp 1745462530
transform 1 0 2712 0 1 2570
box -8 -3 16 105
use FILL  FILL_1683
timestamp 1745462530
transform 1 0 2656 0 1 2570
box -8 -3 16 105
use FILL  FILL_1684
timestamp 1745462530
transform 1 0 2600 0 1 2570
box -8 -3 16 105
use FILL  FILL_1685
timestamp 1745462530
transform 1 0 2592 0 1 2570
box -8 -3 16 105
use FILL  FILL_1686
timestamp 1745462530
transform 1 0 2536 0 1 2570
box -8 -3 16 105
use FILL  FILL_1687
timestamp 1745462530
transform 1 0 2504 0 1 2570
box -8 -3 16 105
use FILL  FILL_1688
timestamp 1745462530
transform 1 0 2496 0 1 2570
box -8 -3 16 105
use FILL  FILL_1689
timestamp 1745462530
transform 1 0 2432 0 1 2570
box -8 -3 16 105
use FILL  FILL_1690
timestamp 1745462530
transform 1 0 2424 0 1 2570
box -8 -3 16 105
use FILL  FILL_1691
timestamp 1745462530
transform 1 0 2376 0 1 2570
box -8 -3 16 105
use FILL  FILL_1692
timestamp 1745462530
transform 1 0 2368 0 1 2570
box -8 -3 16 105
use FILL  FILL_1693
timestamp 1745462530
transform 1 0 2304 0 1 2570
box -8 -3 16 105
use FILL  FILL_1694
timestamp 1745462530
transform 1 0 2296 0 1 2570
box -8 -3 16 105
use FILL  FILL_1695
timestamp 1745462530
transform 1 0 2232 0 1 2570
box -8 -3 16 105
use FILL  FILL_1696
timestamp 1745462530
transform 1 0 2168 0 1 2570
box -8 -3 16 105
use FILL  FILL_1697
timestamp 1745462530
transform 1 0 2104 0 1 2570
box -8 -3 16 105
use FILL  FILL_1698
timestamp 1745462530
transform 1 0 2096 0 1 2570
box -8 -3 16 105
use FILL  FILL_1699
timestamp 1745462530
transform 1 0 1992 0 1 2570
box -8 -3 16 105
use FILL  FILL_1700
timestamp 1745462530
transform 1 0 1984 0 1 2570
box -8 -3 16 105
use FILL  FILL_1701
timestamp 1745462530
transform 1 0 1936 0 1 2570
box -8 -3 16 105
use FILL  FILL_1702
timestamp 1745462530
transform 1 0 1928 0 1 2570
box -8 -3 16 105
use FILL  FILL_1703
timestamp 1745462530
transform 1 0 1880 0 1 2570
box -8 -3 16 105
use FILL  FILL_1704
timestamp 1745462530
transform 1 0 1856 0 1 2570
box -8 -3 16 105
use FILL  FILL_1705
timestamp 1745462530
transform 1 0 1808 0 1 2570
box -8 -3 16 105
use FILL  FILL_1706
timestamp 1745462530
transform 1 0 1800 0 1 2570
box -8 -3 16 105
use FILL  FILL_1707
timestamp 1745462530
transform 1 0 1696 0 1 2570
box -8 -3 16 105
use FILL  FILL_1708
timestamp 1745462530
transform 1 0 1688 0 1 2570
box -8 -3 16 105
use FILL  FILL_1709
timestamp 1745462530
transform 1 0 1664 0 1 2570
box -8 -3 16 105
use FILL  FILL_1710
timestamp 1745462530
transform 1 0 1616 0 1 2570
box -8 -3 16 105
use FILL  FILL_1711
timestamp 1745462530
transform 1 0 1584 0 1 2570
box -8 -3 16 105
use FILL  FILL_1712
timestamp 1745462530
transform 1 0 1576 0 1 2570
box -8 -3 16 105
use FILL  FILL_1713
timestamp 1745462530
transform 1 0 1512 0 1 2570
box -8 -3 16 105
use FILL  FILL_1714
timestamp 1745462530
transform 1 0 1504 0 1 2570
box -8 -3 16 105
use FILL  FILL_1715
timestamp 1745462530
transform 1 0 1456 0 1 2570
box -8 -3 16 105
use FILL  FILL_1716
timestamp 1745462530
transform 1 0 1448 0 1 2570
box -8 -3 16 105
use FILL  FILL_1717
timestamp 1745462530
transform 1 0 1440 0 1 2570
box -8 -3 16 105
use FILL  FILL_1718
timestamp 1745462530
transform 1 0 1408 0 1 2570
box -8 -3 16 105
use FILL  FILL_1719
timestamp 1745462530
transform 1 0 1384 0 1 2570
box -8 -3 16 105
use FILL  FILL_1720
timestamp 1745462530
transform 1 0 1376 0 1 2570
box -8 -3 16 105
use FILL  FILL_1721
timestamp 1745462530
transform 1 0 1304 0 1 2570
box -8 -3 16 105
use FILL  FILL_1722
timestamp 1745462530
transform 1 0 1296 0 1 2570
box -8 -3 16 105
use FILL  FILL_1723
timestamp 1745462530
transform 1 0 1192 0 1 2570
box -8 -3 16 105
use FILL  FILL_1724
timestamp 1745462530
transform 1 0 1184 0 1 2570
box -8 -3 16 105
use FILL  FILL_1725
timestamp 1745462530
transform 1 0 1136 0 1 2570
box -8 -3 16 105
use FILL  FILL_1726
timestamp 1745462530
transform 1 0 1104 0 1 2570
box -8 -3 16 105
use FILL  FILL_1727
timestamp 1745462530
transform 1 0 1096 0 1 2570
box -8 -3 16 105
use FILL  FILL_1728
timestamp 1745462530
transform 1 0 992 0 1 2570
box -8 -3 16 105
use FILL  FILL_1729
timestamp 1745462530
transform 1 0 984 0 1 2570
box -8 -3 16 105
use FILL  FILL_1730
timestamp 1745462530
transform 1 0 936 0 1 2570
box -8 -3 16 105
use FILL  FILL_1731
timestamp 1745462530
transform 1 0 928 0 1 2570
box -8 -3 16 105
use FILL  FILL_1732
timestamp 1745462530
transform 1 0 880 0 1 2570
box -8 -3 16 105
use FILL  FILL_1733
timestamp 1745462530
transform 1 0 832 0 1 2570
box -8 -3 16 105
use FILL  FILL_1734
timestamp 1745462530
transform 1 0 824 0 1 2570
box -8 -3 16 105
use FILL  FILL_1735
timestamp 1745462530
transform 1 0 760 0 1 2570
box -8 -3 16 105
use FILL  FILL_1736
timestamp 1745462530
transform 1 0 752 0 1 2570
box -8 -3 16 105
use FILL  FILL_1737
timestamp 1745462530
transform 1 0 704 0 1 2570
box -8 -3 16 105
use FILL  FILL_1738
timestamp 1745462530
transform 1 0 672 0 1 2570
box -8 -3 16 105
use FILL  FILL_1739
timestamp 1745462530
transform 1 0 664 0 1 2570
box -8 -3 16 105
use FILL  FILL_1740
timestamp 1745462530
transform 1 0 616 0 1 2570
box -8 -3 16 105
use FILL  FILL_1741
timestamp 1745462530
transform 1 0 568 0 1 2570
box -8 -3 16 105
use FILL  FILL_1742
timestamp 1745462530
transform 1 0 560 0 1 2570
box -8 -3 16 105
use FILL  FILL_1743
timestamp 1745462530
transform 1 0 496 0 1 2570
box -8 -3 16 105
use FILL  FILL_1744
timestamp 1745462530
transform 1 0 488 0 1 2570
box -8 -3 16 105
use FILL  FILL_1745
timestamp 1745462530
transform 1 0 384 0 1 2570
box -8 -3 16 105
use FILL  FILL_1746
timestamp 1745462530
transform 1 0 376 0 1 2570
box -8 -3 16 105
use FILL  FILL_1747
timestamp 1745462530
transform 1 0 368 0 1 2570
box -8 -3 16 105
use FILL  FILL_1748
timestamp 1745462530
transform 1 0 304 0 1 2570
box -8 -3 16 105
use FILL  FILL_1749
timestamp 1745462530
transform 1 0 296 0 1 2570
box -8 -3 16 105
use FILL  FILL_1750
timestamp 1745462530
transform 1 0 192 0 1 2570
box -8 -3 16 105
use FILL  FILL_1751
timestamp 1745462530
transform 1 0 184 0 1 2570
box -8 -3 16 105
use FILL  FILL_1752
timestamp 1745462530
transform 1 0 176 0 1 2570
box -8 -3 16 105
use FILL  FILL_1753
timestamp 1745462530
transform 1 0 72 0 1 2570
box -8 -3 16 105
use FILL  FILL_1754
timestamp 1745462530
transform 1 0 4368 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1755
timestamp 1745462530
transform 1 0 4264 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1756
timestamp 1745462530
transform 1 0 4256 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1757
timestamp 1745462530
transform 1 0 4192 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1758
timestamp 1745462530
transform 1 0 4144 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1759
timestamp 1745462530
transform 1 0 4104 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1760
timestamp 1745462530
transform 1 0 4040 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1761
timestamp 1745462530
transform 1 0 4032 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1762
timestamp 1745462530
transform 1 0 3984 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1763
timestamp 1745462530
transform 1 0 3976 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1764
timestamp 1745462530
transform 1 0 3872 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1765
timestamp 1745462530
transform 1 0 3864 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1766
timestamp 1745462530
transform 1 0 3816 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1767
timestamp 1745462530
transform 1 0 3792 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1768
timestamp 1745462530
transform 1 0 3752 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1769
timestamp 1745462530
transform 1 0 3744 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1770
timestamp 1745462530
transform 1 0 3712 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1771
timestamp 1745462530
transform 1 0 3704 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1772
timestamp 1745462530
transform 1 0 3656 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1773
timestamp 1745462530
transform 1 0 3648 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1774
timestamp 1745462530
transform 1 0 3640 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1775
timestamp 1745462530
transform 1 0 3600 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1776
timestamp 1745462530
transform 1 0 3592 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1777
timestamp 1745462530
transform 1 0 3584 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1778
timestamp 1745462530
transform 1 0 3552 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1779
timestamp 1745462530
transform 1 0 3544 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1780
timestamp 1745462530
transform 1 0 3536 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1781
timestamp 1745462530
transform 1 0 3488 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1782
timestamp 1745462530
transform 1 0 3480 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1783
timestamp 1745462530
transform 1 0 3472 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1784
timestamp 1745462530
transform 1 0 3368 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1785
timestamp 1745462530
transform 1 0 3360 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1786
timestamp 1745462530
transform 1 0 3352 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1787
timestamp 1745462530
transform 1 0 3248 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1788
timestamp 1745462530
transform 1 0 3240 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1789
timestamp 1745462530
transform 1 0 3200 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1790
timestamp 1745462530
transform 1 0 3192 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1791
timestamp 1745462530
transform 1 0 3152 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1792
timestamp 1745462530
transform 1 0 3120 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1793
timestamp 1745462530
transform 1 0 3112 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1794
timestamp 1745462530
transform 1 0 3104 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1795
timestamp 1745462530
transform 1 0 3056 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1796
timestamp 1745462530
transform 1 0 3048 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1797
timestamp 1745462530
transform 1 0 2944 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1798
timestamp 1745462530
transform 1 0 2936 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1799
timestamp 1745462530
transform 1 0 2912 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1800
timestamp 1745462530
transform 1 0 2904 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1801
timestamp 1745462530
transform 1 0 2896 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1802
timestamp 1745462530
transform 1 0 2848 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1803
timestamp 1745462530
transform 1 0 2840 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1804
timestamp 1745462530
transform 1 0 2832 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1805
timestamp 1745462530
transform 1 0 2808 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1806
timestamp 1745462530
transform 1 0 2800 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1807
timestamp 1745462530
transform 1 0 2752 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1808
timestamp 1745462530
transform 1 0 2744 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1809
timestamp 1745462530
transform 1 0 2736 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1810
timestamp 1745462530
transform 1 0 2728 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1811
timestamp 1745462530
transform 1 0 2696 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1812
timestamp 1745462530
transform 1 0 2664 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1813
timestamp 1745462530
transform 1 0 2656 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1814
timestamp 1745462530
transform 1 0 2632 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1815
timestamp 1745462530
transform 1 0 2600 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1816
timestamp 1745462530
transform 1 0 2592 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1817
timestamp 1745462530
transform 1 0 2560 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1818
timestamp 1745462530
transform 1 0 2528 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1819
timestamp 1745462530
transform 1 0 2488 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1820
timestamp 1745462530
transform 1 0 2480 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1821
timestamp 1745462530
transform 1 0 2448 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1822
timestamp 1745462530
transform 1 0 2440 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1823
timestamp 1745462530
transform 1 0 2408 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1824
timestamp 1745462530
transform 1 0 2400 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1825
timestamp 1745462530
transform 1 0 2352 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1826
timestamp 1745462530
transform 1 0 2344 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1827
timestamp 1745462530
transform 1 0 2336 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1828
timestamp 1745462530
transform 1 0 2296 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1829
timestamp 1745462530
transform 1 0 2288 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1830
timestamp 1745462530
transform 1 0 2248 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1831
timestamp 1745462530
transform 1 0 2240 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1832
timestamp 1745462530
transform 1 0 2232 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1833
timestamp 1745462530
transform 1 0 2176 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1834
timestamp 1745462530
transform 1 0 2168 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1835
timestamp 1745462530
transform 1 0 2104 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1836
timestamp 1745462530
transform 1 0 2072 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1837
timestamp 1745462530
transform 1 0 2064 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1838
timestamp 1745462530
transform 1 0 2056 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1839
timestamp 1745462530
transform 1 0 2016 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1840
timestamp 1745462530
transform 1 0 1992 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1841
timestamp 1745462530
transform 1 0 1984 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1842
timestamp 1745462530
transform 1 0 1936 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1843
timestamp 1745462530
transform 1 0 1928 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1844
timestamp 1745462530
transform 1 0 1896 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1845
timestamp 1745462530
transform 1 0 1888 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1846
timestamp 1745462530
transform 1 0 1848 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1847
timestamp 1745462530
transform 1 0 1824 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1848
timestamp 1745462530
transform 1 0 1816 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1849
timestamp 1745462530
transform 1 0 1808 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1850
timestamp 1745462530
transform 1 0 1760 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1851
timestamp 1745462530
transform 1 0 1752 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1852
timestamp 1745462530
transform 1 0 1744 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1853
timestamp 1745462530
transform 1 0 1696 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1854
timestamp 1745462530
transform 1 0 1688 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1855
timestamp 1745462530
transform 1 0 1584 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1856
timestamp 1745462530
transform 1 0 1560 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1857
timestamp 1745462530
transform 1 0 1552 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1858
timestamp 1745462530
transform 1 0 1504 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1859
timestamp 1745462530
transform 1 0 1496 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1860
timestamp 1745462530
transform 1 0 1488 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1861
timestamp 1745462530
transform 1 0 1448 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1862
timestamp 1745462530
transform 1 0 1440 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1863
timestamp 1745462530
transform 1 0 1416 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1864
timestamp 1745462530
transform 1 0 1408 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1865
timestamp 1745462530
transform 1 0 1368 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1866
timestamp 1745462530
transform 1 0 1360 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1867
timestamp 1745462530
transform 1 0 1352 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1868
timestamp 1745462530
transform 1 0 1304 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1869
timestamp 1745462530
transform 1 0 1296 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1870
timestamp 1745462530
transform 1 0 1288 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1871
timestamp 1745462530
transform 1 0 1224 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1872
timestamp 1745462530
transform 1 0 1216 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1873
timestamp 1745462530
transform 1 0 1168 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1874
timestamp 1745462530
transform 1 0 1144 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1875
timestamp 1745462530
transform 1 0 1136 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1876
timestamp 1745462530
transform 1 0 1032 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1877
timestamp 1745462530
transform 1 0 1024 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1878
timestamp 1745462530
transform 1 0 984 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1879
timestamp 1745462530
transform 1 0 976 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1880
timestamp 1745462530
transform 1 0 936 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1881
timestamp 1745462530
transform 1 0 904 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1882
timestamp 1745462530
transform 1 0 896 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1883
timestamp 1745462530
transform 1 0 792 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1884
timestamp 1745462530
transform 1 0 752 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1885
timestamp 1745462530
transform 1 0 744 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1886
timestamp 1745462530
transform 1 0 664 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1887
timestamp 1745462530
transform 1 0 656 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1888
timestamp 1745462530
transform 1 0 608 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1889
timestamp 1745462530
transform 1 0 560 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1890
timestamp 1745462530
transform 1 0 504 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1891
timestamp 1745462530
transform 1 0 400 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1892
timestamp 1745462530
transform 1 0 240 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1893
timestamp 1745462530
transform 1 0 192 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1894
timestamp 1745462530
transform 1 0 72 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1895
timestamp 1745462530
transform 1 0 4368 0 1 2370
box -8 -3 16 105
use FILL  FILL_1896
timestamp 1745462530
transform 1 0 4360 0 1 2370
box -8 -3 16 105
use FILL  FILL_1897
timestamp 1745462530
transform 1 0 4256 0 1 2370
box -8 -3 16 105
use FILL  FILL_1898
timestamp 1745462530
transform 1 0 4248 0 1 2370
box -8 -3 16 105
use FILL  FILL_1899
timestamp 1745462530
transform 1 0 4200 0 1 2370
box -8 -3 16 105
use FILL  FILL_1900
timestamp 1745462530
transform 1 0 4176 0 1 2370
box -8 -3 16 105
use FILL  FILL_1901
timestamp 1745462530
transform 1 0 4128 0 1 2370
box -8 -3 16 105
use FILL  FILL_1902
timestamp 1745462530
transform 1 0 4120 0 1 2370
box -8 -3 16 105
use FILL  FILL_1903
timestamp 1745462530
transform 1 0 4112 0 1 2370
box -8 -3 16 105
use FILL  FILL_1904
timestamp 1745462530
transform 1 0 4072 0 1 2370
box -8 -3 16 105
use FILL  FILL_1905
timestamp 1745462530
transform 1 0 4040 0 1 2370
box -8 -3 16 105
use FILL  FILL_1906
timestamp 1745462530
transform 1 0 4032 0 1 2370
box -8 -3 16 105
use FILL  FILL_1907
timestamp 1745462530
transform 1 0 4024 0 1 2370
box -8 -3 16 105
use FILL  FILL_1908
timestamp 1745462530
transform 1 0 3976 0 1 2370
box -8 -3 16 105
use FILL  FILL_1909
timestamp 1745462530
transform 1 0 3968 0 1 2370
box -8 -3 16 105
use FILL  FILL_1910
timestamp 1745462530
transform 1 0 3960 0 1 2370
box -8 -3 16 105
use FILL  FILL_1911
timestamp 1745462530
transform 1 0 3936 0 1 2370
box -8 -3 16 105
use FILL  FILL_1912
timestamp 1745462530
transform 1 0 3928 0 1 2370
box -8 -3 16 105
use FILL  FILL_1913
timestamp 1745462530
transform 1 0 3920 0 1 2370
box -8 -3 16 105
use FILL  FILL_1914
timestamp 1745462530
transform 1 0 3872 0 1 2370
box -8 -3 16 105
use FILL  FILL_1915
timestamp 1745462530
transform 1 0 3864 0 1 2370
box -8 -3 16 105
use FILL  FILL_1916
timestamp 1745462530
transform 1 0 3856 0 1 2370
box -8 -3 16 105
use FILL  FILL_1917
timestamp 1745462530
transform 1 0 3816 0 1 2370
box -8 -3 16 105
use FILL  FILL_1918
timestamp 1745462530
transform 1 0 3808 0 1 2370
box -8 -3 16 105
use FILL  FILL_1919
timestamp 1745462530
transform 1 0 3800 0 1 2370
box -8 -3 16 105
use FILL  FILL_1920
timestamp 1745462530
transform 1 0 3696 0 1 2370
box -8 -3 16 105
use FILL  FILL_1921
timestamp 1745462530
transform 1 0 3688 0 1 2370
box -8 -3 16 105
use FILL  FILL_1922
timestamp 1745462530
transform 1 0 3640 0 1 2370
box -8 -3 16 105
use FILL  FILL_1923
timestamp 1745462530
transform 1 0 3632 0 1 2370
box -8 -3 16 105
use FILL  FILL_1924
timestamp 1745462530
transform 1 0 3624 0 1 2370
box -8 -3 16 105
use FILL  FILL_1925
timestamp 1745462530
transform 1 0 3584 0 1 2370
box -8 -3 16 105
use FILL  FILL_1926
timestamp 1745462530
transform 1 0 3576 0 1 2370
box -8 -3 16 105
use FILL  FILL_1927
timestamp 1745462530
transform 1 0 3568 0 1 2370
box -8 -3 16 105
use FILL  FILL_1928
timestamp 1745462530
transform 1 0 3560 0 1 2370
box -8 -3 16 105
use FILL  FILL_1929
timestamp 1745462530
transform 1 0 3512 0 1 2370
box -8 -3 16 105
use FILL  FILL_1930
timestamp 1745462530
transform 1 0 3504 0 1 2370
box -8 -3 16 105
use FILL  FILL_1931
timestamp 1745462530
transform 1 0 3496 0 1 2370
box -8 -3 16 105
use FILL  FILL_1932
timestamp 1745462530
transform 1 0 3488 0 1 2370
box -8 -3 16 105
use FILL  FILL_1933
timestamp 1745462530
transform 1 0 3424 0 1 2370
box -8 -3 16 105
use FILL  FILL_1934
timestamp 1745462530
transform 1 0 3416 0 1 2370
box -8 -3 16 105
use FILL  FILL_1935
timestamp 1745462530
transform 1 0 3408 0 1 2370
box -8 -3 16 105
use FILL  FILL_1936
timestamp 1745462530
transform 1 0 3360 0 1 2370
box -8 -3 16 105
use FILL  FILL_1937
timestamp 1745462530
transform 1 0 3352 0 1 2370
box -8 -3 16 105
use FILL  FILL_1938
timestamp 1745462530
transform 1 0 3328 0 1 2370
box -8 -3 16 105
use FILL  FILL_1939
timestamp 1745462530
transform 1 0 3320 0 1 2370
box -8 -3 16 105
use FILL  FILL_1940
timestamp 1745462530
transform 1 0 3312 0 1 2370
box -8 -3 16 105
use FILL  FILL_1941
timestamp 1745462530
transform 1 0 3264 0 1 2370
box -8 -3 16 105
use FILL  FILL_1942
timestamp 1745462530
transform 1 0 3240 0 1 2370
box -8 -3 16 105
use FILL  FILL_1943
timestamp 1745462530
transform 1 0 3232 0 1 2370
box -8 -3 16 105
use FILL  FILL_1944
timestamp 1745462530
transform 1 0 3184 0 1 2370
box -8 -3 16 105
use FILL  FILL_1945
timestamp 1745462530
transform 1 0 3160 0 1 2370
box -8 -3 16 105
use FILL  FILL_1946
timestamp 1745462530
transform 1 0 3152 0 1 2370
box -8 -3 16 105
use FILL  FILL_1947
timestamp 1745462530
transform 1 0 3144 0 1 2370
box -8 -3 16 105
use FILL  FILL_1948
timestamp 1745462530
transform 1 0 3040 0 1 2370
box -8 -3 16 105
use FILL  FILL_1949
timestamp 1745462530
transform 1 0 3016 0 1 2370
box -8 -3 16 105
use FILL  FILL_1950
timestamp 1745462530
transform 1 0 3008 0 1 2370
box -8 -3 16 105
use FILL  FILL_1951
timestamp 1745462530
transform 1 0 3000 0 1 2370
box -8 -3 16 105
use FILL  FILL_1952
timestamp 1745462530
transform 1 0 2952 0 1 2370
box -8 -3 16 105
use FILL  FILL_1953
timestamp 1745462530
transform 1 0 2944 0 1 2370
box -8 -3 16 105
use FILL  FILL_1954
timestamp 1745462530
transform 1 0 2936 0 1 2370
box -8 -3 16 105
use FILL  FILL_1955
timestamp 1745462530
transform 1 0 2928 0 1 2370
box -8 -3 16 105
use FILL  FILL_1956
timestamp 1745462530
transform 1 0 2880 0 1 2370
box -8 -3 16 105
use FILL  FILL_1957
timestamp 1745462530
transform 1 0 2872 0 1 2370
box -8 -3 16 105
use FILL  FILL_1958
timestamp 1745462530
transform 1 0 2864 0 1 2370
box -8 -3 16 105
use FILL  FILL_1959
timestamp 1745462530
transform 1 0 2856 0 1 2370
box -8 -3 16 105
use FILL  FILL_1960
timestamp 1745462530
transform 1 0 2808 0 1 2370
box -8 -3 16 105
use FILL  FILL_1961
timestamp 1745462530
transform 1 0 2800 0 1 2370
box -8 -3 16 105
use FILL  FILL_1962
timestamp 1745462530
transform 1 0 2792 0 1 2370
box -8 -3 16 105
use FILL  FILL_1963
timestamp 1745462530
transform 1 0 2784 0 1 2370
box -8 -3 16 105
use FILL  FILL_1964
timestamp 1745462530
transform 1 0 2736 0 1 2370
box -8 -3 16 105
use FILL  FILL_1965
timestamp 1745462530
transform 1 0 2728 0 1 2370
box -8 -3 16 105
use FILL  FILL_1966
timestamp 1745462530
transform 1 0 2720 0 1 2370
box -8 -3 16 105
use FILL  FILL_1967
timestamp 1745462530
transform 1 0 2712 0 1 2370
box -8 -3 16 105
use FILL  FILL_1968
timestamp 1745462530
transform 1 0 2664 0 1 2370
box -8 -3 16 105
use FILL  FILL_1969
timestamp 1745462530
transform 1 0 2656 0 1 2370
box -8 -3 16 105
use FILL  FILL_1970
timestamp 1745462530
transform 1 0 2648 0 1 2370
box -8 -3 16 105
use FILL  FILL_1971
timestamp 1745462530
transform 1 0 2616 0 1 2370
box -8 -3 16 105
use FILL  FILL_1972
timestamp 1745462530
transform 1 0 2584 0 1 2370
box -8 -3 16 105
use FILL  FILL_1973
timestamp 1745462530
transform 1 0 2576 0 1 2370
box -8 -3 16 105
use FILL  FILL_1974
timestamp 1745462530
transform 1 0 2536 0 1 2370
box -8 -3 16 105
use FILL  FILL_1975
timestamp 1745462530
transform 1 0 2528 0 1 2370
box -8 -3 16 105
use FILL  FILL_1976
timestamp 1745462530
transform 1 0 2496 0 1 2370
box -8 -3 16 105
use FILL  FILL_1977
timestamp 1745462530
transform 1 0 2464 0 1 2370
box -8 -3 16 105
use FILL  FILL_1978
timestamp 1745462530
transform 1 0 2432 0 1 2370
box -8 -3 16 105
use FILL  FILL_1979
timestamp 1745462530
transform 1 0 2400 0 1 2370
box -8 -3 16 105
use FILL  FILL_1980
timestamp 1745462530
transform 1 0 2392 0 1 2370
box -8 -3 16 105
use FILL  FILL_1981
timestamp 1745462530
transform 1 0 2352 0 1 2370
box -8 -3 16 105
use FILL  FILL_1982
timestamp 1745462530
transform 1 0 2344 0 1 2370
box -8 -3 16 105
use FILL  FILL_1983
timestamp 1745462530
transform 1 0 2336 0 1 2370
box -8 -3 16 105
use FILL  FILL_1984
timestamp 1745462530
transform 1 0 2296 0 1 2370
box -8 -3 16 105
use FILL  FILL_1985
timestamp 1745462530
transform 1 0 2288 0 1 2370
box -8 -3 16 105
use FILL  FILL_1986
timestamp 1745462530
transform 1 0 2248 0 1 2370
box -8 -3 16 105
use FILL  FILL_1987
timestamp 1745462530
transform 1 0 2240 0 1 2370
box -8 -3 16 105
use FILL  FILL_1988
timestamp 1745462530
transform 1 0 2232 0 1 2370
box -8 -3 16 105
use FILL  FILL_1989
timestamp 1745462530
transform 1 0 2224 0 1 2370
box -8 -3 16 105
use FILL  FILL_1990
timestamp 1745462530
transform 1 0 2176 0 1 2370
box -8 -3 16 105
use FILL  FILL_1991
timestamp 1745462530
transform 1 0 2168 0 1 2370
box -8 -3 16 105
use FILL  FILL_1992
timestamp 1745462530
transform 1 0 2160 0 1 2370
box -8 -3 16 105
use FILL  FILL_1993
timestamp 1745462530
transform 1 0 2112 0 1 2370
box -8 -3 16 105
use FILL  FILL_1994
timestamp 1745462530
transform 1 0 2104 0 1 2370
box -8 -3 16 105
use FILL  FILL_1995
timestamp 1745462530
transform 1 0 2072 0 1 2370
box -8 -3 16 105
use FILL  FILL_1996
timestamp 1745462530
transform 1 0 2064 0 1 2370
box -8 -3 16 105
use FILL  FILL_1997
timestamp 1745462530
transform 1 0 2016 0 1 2370
box -8 -3 16 105
use FILL  FILL_1998
timestamp 1745462530
transform 1 0 2008 0 1 2370
box -8 -3 16 105
use FILL  FILL_1999
timestamp 1745462530
transform 1 0 2000 0 1 2370
box -8 -3 16 105
use FILL  FILL_2000
timestamp 1745462530
transform 1 0 1952 0 1 2370
box -8 -3 16 105
use FILL  FILL_2001
timestamp 1745462530
transform 1 0 1944 0 1 2370
box -8 -3 16 105
use FILL  FILL_2002
timestamp 1745462530
transform 1 0 1936 0 1 2370
box -8 -3 16 105
use FILL  FILL_2003
timestamp 1745462530
transform 1 0 1888 0 1 2370
box -8 -3 16 105
use FILL  FILL_2004
timestamp 1745462530
transform 1 0 1880 0 1 2370
box -8 -3 16 105
use FILL  FILL_2005
timestamp 1745462530
transform 1 0 1840 0 1 2370
box -8 -3 16 105
use FILL  FILL_2006
timestamp 1745462530
transform 1 0 1832 0 1 2370
box -8 -3 16 105
use FILL  FILL_2007
timestamp 1745462530
transform 1 0 1808 0 1 2370
box -8 -3 16 105
use FILL  FILL_2008
timestamp 1745462530
transform 1 0 1704 0 1 2370
box -8 -3 16 105
use FILL  FILL_2009
timestamp 1745462530
transform 1 0 1696 0 1 2370
box -8 -3 16 105
use FILL  FILL_2010
timestamp 1745462530
transform 1 0 1688 0 1 2370
box -8 -3 16 105
use FILL  FILL_2011
timestamp 1745462530
transform 1 0 1640 0 1 2370
box -8 -3 16 105
use FILL  FILL_2012
timestamp 1745462530
transform 1 0 1632 0 1 2370
box -8 -3 16 105
use FILL  FILL_2013
timestamp 1745462530
transform 1 0 1624 0 1 2370
box -8 -3 16 105
use FILL  FILL_2014
timestamp 1745462530
transform 1 0 1584 0 1 2370
box -8 -3 16 105
use FILL  FILL_2015
timestamp 1745462530
transform 1 0 1576 0 1 2370
box -8 -3 16 105
use FILL  FILL_2016
timestamp 1745462530
transform 1 0 1568 0 1 2370
box -8 -3 16 105
use FILL  FILL_2017
timestamp 1745462530
transform 1 0 1520 0 1 2370
box -8 -3 16 105
use FILL  FILL_2018
timestamp 1745462530
transform 1 0 1512 0 1 2370
box -8 -3 16 105
use FILL  FILL_2019
timestamp 1745462530
transform 1 0 1504 0 1 2370
box -8 -3 16 105
use FILL  FILL_2020
timestamp 1745462530
transform 1 0 1464 0 1 2370
box -8 -3 16 105
use FILL  FILL_2021
timestamp 1745462530
transform 1 0 1456 0 1 2370
box -8 -3 16 105
use FILL  FILL_2022
timestamp 1745462530
transform 1 0 1448 0 1 2370
box -8 -3 16 105
use FILL  FILL_2023
timestamp 1745462530
transform 1 0 1408 0 1 2370
box -8 -3 16 105
use FILL  FILL_2024
timestamp 1745462530
transform 1 0 1400 0 1 2370
box -8 -3 16 105
use FILL  FILL_2025
timestamp 1745462530
transform 1 0 1392 0 1 2370
box -8 -3 16 105
use FILL  FILL_2026
timestamp 1745462530
transform 1 0 1384 0 1 2370
box -8 -3 16 105
use FILL  FILL_2027
timestamp 1745462530
transform 1 0 1336 0 1 2370
box -8 -3 16 105
use FILL  FILL_2028
timestamp 1745462530
transform 1 0 1328 0 1 2370
box -8 -3 16 105
use FILL  FILL_2029
timestamp 1745462530
transform 1 0 1296 0 1 2370
box -8 -3 16 105
use FILL  FILL_2030
timestamp 1745462530
transform 1 0 1288 0 1 2370
box -8 -3 16 105
use FILL  FILL_2031
timestamp 1745462530
transform 1 0 1280 0 1 2370
box -8 -3 16 105
use FILL  FILL_2032
timestamp 1745462530
transform 1 0 1232 0 1 2370
box -8 -3 16 105
use FILL  FILL_2033
timestamp 1745462530
transform 1 0 1224 0 1 2370
box -8 -3 16 105
use FILL  FILL_2034
timestamp 1745462530
transform 1 0 1216 0 1 2370
box -8 -3 16 105
use FILL  FILL_2035
timestamp 1745462530
transform 1 0 1168 0 1 2370
box -8 -3 16 105
use FILL  FILL_2036
timestamp 1745462530
transform 1 0 1160 0 1 2370
box -8 -3 16 105
use FILL  FILL_2037
timestamp 1745462530
transform 1 0 1128 0 1 2370
box -8 -3 16 105
use FILL  FILL_2038
timestamp 1745462530
transform 1 0 1120 0 1 2370
box -8 -3 16 105
use FILL  FILL_2039
timestamp 1745462530
transform 1 0 1080 0 1 2370
box -8 -3 16 105
use FILL  FILL_2040
timestamp 1745462530
transform 1 0 1072 0 1 2370
box -8 -3 16 105
use FILL  FILL_2041
timestamp 1745462530
transform 1 0 1048 0 1 2370
box -8 -3 16 105
use FILL  FILL_2042
timestamp 1745462530
transform 1 0 1000 0 1 2370
box -8 -3 16 105
use FILL  FILL_2043
timestamp 1745462530
transform 1 0 992 0 1 2370
box -8 -3 16 105
use FILL  FILL_2044
timestamp 1745462530
transform 1 0 944 0 1 2370
box -8 -3 16 105
use FILL  FILL_2045
timestamp 1745462530
transform 1 0 936 0 1 2370
box -8 -3 16 105
use FILL  FILL_2046
timestamp 1745462530
transform 1 0 888 0 1 2370
box -8 -3 16 105
use FILL  FILL_2047
timestamp 1745462530
transform 1 0 832 0 1 2370
box -8 -3 16 105
use FILL  FILL_2048
timestamp 1745462530
transform 1 0 824 0 1 2370
box -8 -3 16 105
use FILL  FILL_2049
timestamp 1745462530
transform 1 0 816 0 1 2370
box -8 -3 16 105
use FILL  FILL_2050
timestamp 1745462530
transform 1 0 784 0 1 2370
box -8 -3 16 105
use FILL  FILL_2051
timestamp 1745462530
transform 1 0 736 0 1 2370
box -8 -3 16 105
use FILL  FILL_2052
timestamp 1745462530
transform 1 0 728 0 1 2370
box -8 -3 16 105
use FILL  FILL_2053
timestamp 1745462530
transform 1 0 680 0 1 2370
box -8 -3 16 105
use FILL  FILL_2054
timestamp 1745462530
transform 1 0 672 0 1 2370
box -8 -3 16 105
use FILL  FILL_2055
timestamp 1745462530
transform 1 0 640 0 1 2370
box -8 -3 16 105
use FILL  FILL_2056
timestamp 1745462530
transform 1 0 600 0 1 2370
box -8 -3 16 105
use FILL  FILL_2057
timestamp 1745462530
transform 1 0 592 0 1 2370
box -8 -3 16 105
use FILL  FILL_2058
timestamp 1745462530
transform 1 0 488 0 1 2370
box -8 -3 16 105
use FILL  FILL_2059
timestamp 1745462530
transform 1 0 480 0 1 2370
box -8 -3 16 105
use FILL  FILL_2060
timestamp 1745462530
transform 1 0 424 0 1 2370
box -8 -3 16 105
use FILL  FILL_2061
timestamp 1745462530
transform 1 0 376 0 1 2370
box -8 -3 16 105
use FILL  FILL_2062
timestamp 1745462530
transform 1 0 368 0 1 2370
box -8 -3 16 105
use FILL  FILL_2063
timestamp 1745462530
transform 1 0 264 0 1 2370
box -8 -3 16 105
use FILL  FILL_2064
timestamp 1745462530
transform 1 0 240 0 1 2370
box -8 -3 16 105
use FILL  FILL_2065
timestamp 1745462530
transform 1 0 176 0 1 2370
box -8 -3 16 105
use FILL  FILL_2066
timestamp 1745462530
transform 1 0 72 0 1 2370
box -8 -3 16 105
use FILL  FILL_2067
timestamp 1745462530
transform 1 0 4272 0 -1 2370
box -8 -3 16 105
use FILL  FILL_2068
timestamp 1745462530
transform 1 0 4208 0 -1 2370
box -8 -3 16 105
use FILL  FILL_2069
timestamp 1745462530
transform 1 0 4144 0 -1 2370
box -8 -3 16 105
use FILL  FILL_2070
timestamp 1745462530
transform 1 0 4136 0 -1 2370
box -8 -3 16 105
use FILL  FILL_2071
timestamp 1745462530
transform 1 0 4064 0 -1 2370
box -8 -3 16 105
use FILL  FILL_2072
timestamp 1745462530
transform 1 0 3960 0 -1 2370
box -8 -3 16 105
use FILL  FILL_2073
timestamp 1745462530
transform 1 0 3896 0 -1 2370
box -8 -3 16 105
use FILL  FILL_2074
timestamp 1745462530
transform 1 0 3888 0 -1 2370
box -8 -3 16 105
use FILL  FILL_2075
timestamp 1745462530
transform 1 0 3848 0 -1 2370
box -8 -3 16 105
use FILL  FILL_2076
timestamp 1745462530
transform 1 0 3840 0 -1 2370
box -8 -3 16 105
use FILL  FILL_2077
timestamp 1745462530
transform 1 0 3792 0 -1 2370
box -8 -3 16 105
use FILL  FILL_2078
timestamp 1745462530
transform 1 0 3760 0 -1 2370
box -8 -3 16 105
use FILL  FILL_2079
timestamp 1745462530
transform 1 0 3752 0 -1 2370
box -8 -3 16 105
use FILL  FILL_2080
timestamp 1745462530
transform 1 0 3648 0 -1 2370
box -8 -3 16 105
use FILL  FILL_2081
timestamp 1745462530
transform 1 0 3600 0 -1 2370
box -8 -3 16 105
use FILL  FILL_2082
timestamp 1745462530
transform 1 0 3592 0 -1 2370
box -8 -3 16 105
use FILL  FILL_2083
timestamp 1745462530
transform 1 0 3584 0 -1 2370
box -8 -3 16 105
use FILL  FILL_2084
timestamp 1745462530
transform 1 0 3536 0 -1 2370
box -8 -3 16 105
use FILL  FILL_2085
timestamp 1745462530
transform 1 0 3528 0 -1 2370
box -8 -3 16 105
use FILL  FILL_2086
timestamp 1745462530
transform 1 0 3400 0 -1 2370
box -8 -3 16 105
use FILL  FILL_2087
timestamp 1745462530
transform 1 0 3352 0 -1 2370
box -8 -3 16 105
use FILL  FILL_2088
timestamp 1745462530
transform 1 0 3344 0 -1 2370
box -8 -3 16 105
use FILL  FILL_2089
timestamp 1745462530
transform 1 0 3336 0 -1 2370
box -8 -3 16 105
use FILL  FILL_2090
timestamp 1745462530
transform 1 0 3288 0 -1 2370
box -8 -3 16 105
use FILL  FILL_2091
timestamp 1745462530
transform 1 0 3280 0 -1 2370
box -8 -3 16 105
use FILL  FILL_2092
timestamp 1745462530
transform 1 0 3272 0 -1 2370
box -8 -3 16 105
use FILL  FILL_2093
timestamp 1745462530
transform 1 0 3224 0 -1 2370
box -8 -3 16 105
use FILL  FILL_2094
timestamp 1745462530
transform 1 0 3216 0 -1 2370
box -8 -3 16 105
use FILL  FILL_2095
timestamp 1745462530
transform 1 0 3112 0 -1 2370
box -8 -3 16 105
use FILL  FILL_2096
timestamp 1745462530
transform 1 0 3104 0 -1 2370
box -8 -3 16 105
use FILL  FILL_2097
timestamp 1745462530
transform 1 0 3064 0 -1 2370
box -8 -3 16 105
use FILL  FILL_2098
timestamp 1745462530
transform 1 0 3056 0 -1 2370
box -8 -3 16 105
use FILL  FILL_2099
timestamp 1745462530
transform 1 0 3016 0 -1 2370
box -8 -3 16 105
use FILL  FILL_2100
timestamp 1745462530
transform 1 0 3008 0 -1 2370
box -8 -3 16 105
use FILL  FILL_2101
timestamp 1745462530
transform 1 0 3000 0 -1 2370
box -8 -3 16 105
use FILL  FILL_2102
timestamp 1745462530
transform 1 0 2960 0 -1 2370
box -8 -3 16 105
use FILL  FILL_2103
timestamp 1745462530
transform 1 0 2952 0 -1 2370
box -8 -3 16 105
use FILL  FILL_2104
timestamp 1745462530
transform 1 0 2912 0 -1 2370
box -8 -3 16 105
use FILL  FILL_2105
timestamp 1745462530
transform 1 0 2904 0 -1 2370
box -8 -3 16 105
use FILL  FILL_2106
timestamp 1745462530
transform 1 0 2872 0 -1 2370
box -8 -3 16 105
use FILL  FILL_2107
timestamp 1745462530
transform 1 0 2768 0 -1 2370
box -8 -3 16 105
use FILL  FILL_2108
timestamp 1745462530
transform 1 0 2664 0 -1 2370
box -8 -3 16 105
use FILL  FILL_2109
timestamp 1745462530
transform 1 0 2632 0 -1 2370
box -8 -3 16 105
use FILL  FILL_2110
timestamp 1745462530
transform 1 0 2624 0 -1 2370
box -8 -3 16 105
use FILL  FILL_2111
timestamp 1745462530
transform 1 0 2576 0 -1 2370
box -8 -3 16 105
use FILL  FILL_2112
timestamp 1745462530
transform 1 0 2568 0 -1 2370
box -8 -3 16 105
use FILL  FILL_2113
timestamp 1745462530
transform 1 0 2512 0 -1 2370
box -8 -3 16 105
use FILL  FILL_2114
timestamp 1745462530
transform 1 0 2456 0 -1 2370
box -8 -3 16 105
use FILL  FILL_2115
timestamp 1745462530
transform 1 0 2424 0 -1 2370
box -8 -3 16 105
use FILL  FILL_2116
timestamp 1745462530
transform 1 0 2416 0 -1 2370
box -8 -3 16 105
use FILL  FILL_2117
timestamp 1745462530
transform 1 0 2384 0 -1 2370
box -8 -3 16 105
use FILL  FILL_2118
timestamp 1745462530
transform 1 0 2344 0 -1 2370
box -8 -3 16 105
use FILL  FILL_2119
timestamp 1745462530
transform 1 0 2336 0 -1 2370
box -8 -3 16 105
use FILL  FILL_2120
timestamp 1745462530
transform 1 0 2328 0 -1 2370
box -8 -3 16 105
use FILL  FILL_2121
timestamp 1745462530
transform 1 0 2288 0 -1 2370
box -8 -3 16 105
use FILL  FILL_2122
timestamp 1745462530
transform 1 0 2248 0 -1 2370
box -8 -3 16 105
use FILL  FILL_2123
timestamp 1745462530
transform 1 0 2240 0 -1 2370
box -8 -3 16 105
use FILL  FILL_2124
timestamp 1745462530
transform 1 0 2200 0 -1 2370
box -8 -3 16 105
use FILL  FILL_2125
timestamp 1745462530
transform 1 0 2192 0 -1 2370
box -8 -3 16 105
use FILL  FILL_2126
timestamp 1745462530
transform 1 0 2152 0 -1 2370
box -8 -3 16 105
use FILL  FILL_2127
timestamp 1745462530
transform 1 0 2120 0 -1 2370
box -8 -3 16 105
use FILL  FILL_2128
timestamp 1745462530
transform 1 0 2112 0 -1 2370
box -8 -3 16 105
use FILL  FILL_2129
timestamp 1745462530
transform 1 0 2080 0 -1 2370
box -8 -3 16 105
use FILL  FILL_2130
timestamp 1745462530
transform 1 0 2040 0 -1 2370
box -8 -3 16 105
use FILL  FILL_2131
timestamp 1745462530
transform 1 0 2032 0 -1 2370
box -8 -3 16 105
use FILL  FILL_2132
timestamp 1745462530
transform 1 0 1984 0 -1 2370
box -8 -3 16 105
use FILL  FILL_2133
timestamp 1745462530
transform 1 0 1976 0 -1 2370
box -8 -3 16 105
use FILL  FILL_2134
timestamp 1745462530
transform 1 0 1912 0 -1 2370
box -8 -3 16 105
use FILL  FILL_2135
timestamp 1745462530
transform 1 0 1904 0 -1 2370
box -8 -3 16 105
use FILL  FILL_2136
timestamp 1745462530
transform 1 0 1896 0 -1 2370
box -8 -3 16 105
use FILL  FILL_2137
timestamp 1745462530
transform 1 0 1848 0 -1 2370
box -8 -3 16 105
use FILL  FILL_2138
timestamp 1745462530
transform 1 0 1816 0 -1 2370
box -8 -3 16 105
use FILL  FILL_2139
timestamp 1745462530
transform 1 0 1808 0 -1 2370
box -8 -3 16 105
use FILL  FILL_2140
timestamp 1745462530
transform 1 0 1760 0 -1 2370
box -8 -3 16 105
use FILL  FILL_2141
timestamp 1745462530
transform 1 0 1752 0 -1 2370
box -8 -3 16 105
use FILL  FILL_2142
timestamp 1745462530
transform 1 0 1744 0 -1 2370
box -8 -3 16 105
use FILL  FILL_2143
timestamp 1745462530
transform 1 0 1696 0 -1 2370
box -8 -3 16 105
use FILL  FILL_2144
timestamp 1745462530
transform 1 0 1688 0 -1 2370
box -8 -3 16 105
use FILL  FILL_2145
timestamp 1745462530
transform 1 0 1640 0 -1 2370
box -8 -3 16 105
use FILL  FILL_2146
timestamp 1745462530
transform 1 0 1632 0 -1 2370
box -8 -3 16 105
use FILL  FILL_2147
timestamp 1745462530
transform 1 0 1600 0 -1 2370
box -8 -3 16 105
use FILL  FILL_2148
timestamp 1745462530
transform 1 0 1592 0 -1 2370
box -8 -3 16 105
use FILL  FILL_2149
timestamp 1745462530
transform 1 0 1544 0 -1 2370
box -8 -3 16 105
use FILL  FILL_2150
timestamp 1745462530
transform 1 0 1536 0 -1 2370
box -8 -3 16 105
use FILL  FILL_2151
timestamp 1745462530
transform 1 0 1496 0 -1 2370
box -8 -3 16 105
use FILL  FILL_2152
timestamp 1745462530
transform 1 0 1488 0 -1 2370
box -8 -3 16 105
use FILL  FILL_2153
timestamp 1745462530
transform 1 0 1480 0 -1 2370
box -8 -3 16 105
use FILL  FILL_2154
timestamp 1745462530
transform 1 0 1432 0 -1 2370
box -8 -3 16 105
use FILL  FILL_2155
timestamp 1745462530
transform 1 0 1400 0 -1 2370
box -8 -3 16 105
use FILL  FILL_2156
timestamp 1745462530
transform 1 0 1392 0 -1 2370
box -8 -3 16 105
use FILL  FILL_2157
timestamp 1745462530
transform 1 0 1384 0 -1 2370
box -8 -3 16 105
use FILL  FILL_2158
timestamp 1745462530
transform 1 0 1336 0 -1 2370
box -8 -3 16 105
use FILL  FILL_2159
timestamp 1745462530
transform 1 0 1328 0 -1 2370
box -8 -3 16 105
use FILL  FILL_2160
timestamp 1745462530
transform 1 0 1296 0 -1 2370
box -8 -3 16 105
use FILL  FILL_2161
timestamp 1745462530
transform 1 0 1288 0 -1 2370
box -8 -3 16 105
use FILL  FILL_2162
timestamp 1745462530
transform 1 0 1240 0 -1 2370
box -8 -3 16 105
use FILL  FILL_2163
timestamp 1745462530
transform 1 0 1232 0 -1 2370
box -8 -3 16 105
use FILL  FILL_2164
timestamp 1745462530
transform 1 0 1224 0 -1 2370
box -8 -3 16 105
use FILL  FILL_2165
timestamp 1745462530
transform 1 0 1176 0 -1 2370
box -8 -3 16 105
use FILL  FILL_2166
timestamp 1745462530
transform 1 0 1168 0 -1 2370
box -8 -3 16 105
use FILL  FILL_2167
timestamp 1745462530
transform 1 0 1160 0 -1 2370
box -8 -3 16 105
use FILL  FILL_2168
timestamp 1745462530
transform 1 0 1112 0 -1 2370
box -8 -3 16 105
use FILL  FILL_2169
timestamp 1745462530
transform 1 0 1104 0 -1 2370
box -8 -3 16 105
use FILL  FILL_2170
timestamp 1745462530
transform 1 0 1000 0 -1 2370
box -8 -3 16 105
use FILL  FILL_2171
timestamp 1745462530
transform 1 0 992 0 -1 2370
box -8 -3 16 105
use FILL  FILL_2172
timestamp 1745462530
transform 1 0 888 0 -1 2370
box -8 -3 16 105
use FILL  FILL_2173
timestamp 1745462530
transform 1 0 880 0 -1 2370
box -8 -3 16 105
use FILL  FILL_2174
timestamp 1745462530
transform 1 0 840 0 -1 2370
box -8 -3 16 105
use FILL  FILL_2175
timestamp 1745462530
transform 1 0 808 0 -1 2370
box -8 -3 16 105
use FILL  FILL_2176
timestamp 1745462530
transform 1 0 768 0 -1 2370
box -8 -3 16 105
use FILL  FILL_2177
timestamp 1745462530
transform 1 0 760 0 -1 2370
box -8 -3 16 105
use FILL  FILL_2178
timestamp 1745462530
transform 1 0 752 0 -1 2370
box -8 -3 16 105
use FILL  FILL_2179
timestamp 1745462530
transform 1 0 704 0 -1 2370
box -8 -3 16 105
use FILL  FILL_2180
timestamp 1745462530
transform 1 0 672 0 -1 2370
box -8 -3 16 105
use FILL  FILL_2181
timestamp 1745462530
transform 1 0 664 0 -1 2370
box -8 -3 16 105
use FILL  FILL_2182
timestamp 1745462530
transform 1 0 616 0 -1 2370
box -8 -3 16 105
use FILL  FILL_2183
timestamp 1745462530
transform 1 0 608 0 -1 2370
box -8 -3 16 105
use FILL  FILL_2184
timestamp 1745462530
transform 1 0 568 0 -1 2370
box -8 -3 16 105
use FILL  FILL_2185
timestamp 1745462530
transform 1 0 528 0 -1 2370
box -8 -3 16 105
use FILL  FILL_2186
timestamp 1745462530
transform 1 0 520 0 -1 2370
box -8 -3 16 105
use FILL  FILL_2187
timestamp 1745462530
transform 1 0 512 0 -1 2370
box -8 -3 16 105
use FILL  FILL_2188
timestamp 1745462530
transform 1 0 408 0 -1 2370
box -8 -3 16 105
use FILL  FILL_2189
timestamp 1745462530
transform 1 0 400 0 -1 2370
box -8 -3 16 105
use FILL  FILL_2190
timestamp 1745462530
transform 1 0 336 0 -1 2370
box -8 -3 16 105
use FILL  FILL_2191
timestamp 1745462530
transform 1 0 328 0 -1 2370
box -8 -3 16 105
use FILL  FILL_2192
timestamp 1745462530
transform 1 0 320 0 -1 2370
box -8 -3 16 105
use FILL  FILL_2193
timestamp 1745462530
transform 1 0 256 0 -1 2370
box -8 -3 16 105
use FILL  FILL_2194
timestamp 1745462530
transform 1 0 248 0 -1 2370
box -8 -3 16 105
use FILL  FILL_2195
timestamp 1745462530
transform 1 0 240 0 -1 2370
box -8 -3 16 105
use FILL  FILL_2196
timestamp 1745462530
transform 1 0 232 0 -1 2370
box -8 -3 16 105
use FILL  FILL_2197
timestamp 1745462530
transform 1 0 168 0 -1 2370
box -8 -3 16 105
use FILL  FILL_2198
timestamp 1745462530
transform 1 0 160 0 -1 2370
box -8 -3 16 105
use FILL  FILL_2199
timestamp 1745462530
transform 1 0 152 0 -1 2370
box -8 -3 16 105
use FILL  FILL_2200
timestamp 1745462530
transform 1 0 144 0 -1 2370
box -8 -3 16 105
use FILL  FILL_2201
timestamp 1745462530
transform 1 0 136 0 -1 2370
box -8 -3 16 105
use FILL  FILL_2202
timestamp 1745462530
transform 1 0 128 0 -1 2370
box -8 -3 16 105
use FILL  FILL_2203
timestamp 1745462530
transform 1 0 120 0 -1 2370
box -8 -3 16 105
use FILL  FILL_2204
timestamp 1745462530
transform 1 0 112 0 -1 2370
box -8 -3 16 105
use FILL  FILL_2205
timestamp 1745462530
transform 1 0 104 0 -1 2370
box -8 -3 16 105
use FILL  FILL_2206
timestamp 1745462530
transform 1 0 96 0 -1 2370
box -8 -3 16 105
use FILL  FILL_2207
timestamp 1745462530
transform 1 0 88 0 -1 2370
box -8 -3 16 105
use FILL  FILL_2208
timestamp 1745462530
transform 1 0 80 0 -1 2370
box -8 -3 16 105
use FILL  FILL_2209
timestamp 1745462530
transform 1 0 72 0 -1 2370
box -8 -3 16 105
use FILL  FILL_2210
timestamp 1745462530
transform 1 0 4368 0 1 2170
box -8 -3 16 105
use FILL  FILL_2211
timestamp 1745462530
transform 1 0 4248 0 1 2170
box -8 -3 16 105
use FILL  FILL_2212
timestamp 1745462530
transform 1 0 4128 0 1 2170
box -8 -3 16 105
use FILL  FILL_2213
timestamp 1745462530
transform 1 0 4080 0 1 2170
box -8 -3 16 105
use FILL  FILL_2214
timestamp 1745462530
transform 1 0 4048 0 1 2170
box -8 -3 16 105
use FILL  FILL_2215
timestamp 1745462530
transform 1 0 4040 0 1 2170
box -8 -3 16 105
use FILL  FILL_2216
timestamp 1745462530
transform 1 0 3936 0 1 2170
box -8 -3 16 105
use FILL  FILL_2217
timestamp 1745462530
transform 1 0 3928 0 1 2170
box -8 -3 16 105
use FILL  FILL_2218
timestamp 1745462530
transform 1 0 3880 0 1 2170
box -8 -3 16 105
use FILL  FILL_2219
timestamp 1745462530
transform 1 0 3832 0 1 2170
box -8 -3 16 105
use FILL  FILL_2220
timestamp 1745462530
transform 1 0 3824 0 1 2170
box -8 -3 16 105
use FILL  FILL_2221
timestamp 1745462530
transform 1 0 3792 0 1 2170
box -8 -3 16 105
use FILL  FILL_2222
timestamp 1745462530
transform 1 0 3752 0 1 2170
box -8 -3 16 105
use FILL  FILL_2223
timestamp 1745462530
transform 1 0 3728 0 1 2170
box -8 -3 16 105
use FILL  FILL_2224
timestamp 1745462530
transform 1 0 3624 0 1 2170
box -8 -3 16 105
use FILL  FILL_2225
timestamp 1745462530
transform 1 0 3616 0 1 2170
box -8 -3 16 105
use FILL  FILL_2226
timestamp 1745462530
transform 1 0 3608 0 1 2170
box -8 -3 16 105
use FILL  FILL_2227
timestamp 1745462530
transform 1 0 3560 0 1 2170
box -8 -3 16 105
use FILL  FILL_2228
timestamp 1745462530
transform 1 0 3552 0 1 2170
box -8 -3 16 105
use FILL  FILL_2229
timestamp 1745462530
transform 1 0 3544 0 1 2170
box -8 -3 16 105
use FILL  FILL_2230
timestamp 1745462530
transform 1 0 3520 0 1 2170
box -8 -3 16 105
use FILL  FILL_2231
timestamp 1745462530
transform 1 0 3416 0 1 2170
box -8 -3 16 105
use FILL  FILL_2232
timestamp 1745462530
transform 1 0 3408 0 1 2170
box -8 -3 16 105
use FILL  FILL_2233
timestamp 1745462530
transform 1 0 3360 0 1 2170
box -8 -3 16 105
use FILL  FILL_2234
timestamp 1745462530
transform 1 0 3352 0 1 2170
box -8 -3 16 105
use FILL  FILL_2235
timestamp 1745462530
transform 1 0 3344 0 1 2170
box -8 -3 16 105
use FILL  FILL_2236
timestamp 1745462530
transform 1 0 3336 0 1 2170
box -8 -3 16 105
use FILL  FILL_2237
timestamp 1745462530
transform 1 0 3288 0 1 2170
box -8 -3 16 105
use FILL  FILL_2238
timestamp 1745462530
transform 1 0 3280 0 1 2170
box -8 -3 16 105
use FILL  FILL_2239
timestamp 1745462530
transform 1 0 3160 0 1 2170
box -8 -3 16 105
use FILL  FILL_2240
timestamp 1745462530
transform 1 0 3152 0 1 2170
box -8 -3 16 105
use FILL  FILL_2241
timestamp 1745462530
transform 1 0 3144 0 1 2170
box -8 -3 16 105
use FILL  FILL_2242
timestamp 1745462530
transform 1 0 3096 0 1 2170
box -8 -3 16 105
use FILL  FILL_2243
timestamp 1745462530
transform 1 0 3088 0 1 2170
box -8 -3 16 105
use FILL  FILL_2244
timestamp 1745462530
transform 1 0 2968 0 1 2170
box -8 -3 16 105
use FILL  FILL_2245
timestamp 1745462530
transform 1 0 2960 0 1 2170
box -8 -3 16 105
use FILL  FILL_2246
timestamp 1745462530
transform 1 0 2912 0 1 2170
box -8 -3 16 105
use FILL  FILL_2247
timestamp 1745462530
transform 1 0 2904 0 1 2170
box -8 -3 16 105
use FILL  FILL_2248
timestamp 1745462530
transform 1 0 2896 0 1 2170
box -8 -3 16 105
use FILL  FILL_2249
timestamp 1745462530
transform 1 0 2832 0 1 2170
box -8 -3 16 105
use FILL  FILL_2250
timestamp 1745462530
transform 1 0 2824 0 1 2170
box -8 -3 16 105
use FILL  FILL_2251
timestamp 1745462530
transform 1 0 2816 0 1 2170
box -8 -3 16 105
use FILL  FILL_2252
timestamp 1745462530
transform 1 0 2768 0 1 2170
box -8 -3 16 105
use FILL  FILL_2253
timestamp 1745462530
transform 1 0 2760 0 1 2170
box -8 -3 16 105
use FILL  FILL_2254
timestamp 1745462530
transform 1 0 2656 0 1 2170
box -8 -3 16 105
use FILL  FILL_2255
timestamp 1745462530
transform 1 0 2608 0 1 2170
box -8 -3 16 105
use FILL  FILL_2256
timestamp 1745462530
transform 1 0 2600 0 1 2170
box -8 -3 16 105
use FILL  FILL_2257
timestamp 1745462530
transform 1 0 2576 0 1 2170
box -8 -3 16 105
use FILL  FILL_2258
timestamp 1745462530
transform 1 0 2472 0 1 2170
box -8 -3 16 105
use FILL  FILL_2259
timestamp 1745462530
transform 1 0 2440 0 1 2170
box -8 -3 16 105
use FILL  FILL_2260
timestamp 1745462530
transform 1 0 2408 0 1 2170
box -8 -3 16 105
use FILL  FILL_2261
timestamp 1745462530
transform 1 0 2376 0 1 2170
box -8 -3 16 105
use FILL  FILL_2262
timestamp 1745462530
transform 1 0 2368 0 1 2170
box -8 -3 16 105
use FILL  FILL_2263
timestamp 1745462530
transform 1 0 2312 0 1 2170
box -8 -3 16 105
use FILL  FILL_2264
timestamp 1745462530
transform 1 0 2304 0 1 2170
box -8 -3 16 105
use FILL  FILL_2265
timestamp 1745462530
transform 1 0 2264 0 1 2170
box -8 -3 16 105
use FILL  FILL_2266
timestamp 1745462530
transform 1 0 2256 0 1 2170
box -8 -3 16 105
use FILL  FILL_2267
timestamp 1745462530
transform 1 0 2248 0 1 2170
box -8 -3 16 105
use FILL  FILL_2268
timestamp 1745462530
transform 1 0 2208 0 1 2170
box -8 -3 16 105
use FILL  FILL_2269
timestamp 1745462530
transform 1 0 2184 0 1 2170
box -8 -3 16 105
use FILL  FILL_2270
timestamp 1745462530
transform 1 0 2144 0 1 2170
box -8 -3 16 105
use FILL  FILL_2271
timestamp 1745462530
transform 1 0 2136 0 1 2170
box -8 -3 16 105
use FILL  FILL_2272
timestamp 1745462530
transform 1 0 2032 0 1 2170
box -8 -3 16 105
use FILL  FILL_2273
timestamp 1745462530
transform 1 0 2008 0 1 2170
box -8 -3 16 105
use FILL  FILL_2274
timestamp 1745462530
transform 1 0 1960 0 1 2170
box -8 -3 16 105
use FILL  FILL_2275
timestamp 1745462530
transform 1 0 1952 0 1 2170
box -8 -3 16 105
use FILL  FILL_2276
timestamp 1745462530
transform 1 0 1944 0 1 2170
box -8 -3 16 105
use FILL  FILL_2277
timestamp 1745462530
transform 1 0 1880 0 1 2170
box -8 -3 16 105
use FILL  FILL_2278
timestamp 1745462530
transform 1 0 1872 0 1 2170
box -8 -3 16 105
use FILL  FILL_2279
timestamp 1745462530
transform 1 0 1816 0 1 2170
box -8 -3 16 105
use FILL  FILL_2280
timestamp 1745462530
transform 1 0 1808 0 1 2170
box -8 -3 16 105
use FILL  FILL_2281
timestamp 1745462530
transform 1 0 1744 0 1 2170
box -8 -3 16 105
use FILL  FILL_2282
timestamp 1745462530
transform 1 0 1736 0 1 2170
box -8 -3 16 105
use FILL  FILL_2283
timestamp 1745462530
transform 1 0 1728 0 1 2170
box -8 -3 16 105
use FILL  FILL_2284
timestamp 1745462530
transform 1 0 1680 0 1 2170
box -8 -3 16 105
use FILL  FILL_2285
timestamp 1745462530
transform 1 0 1672 0 1 2170
box -8 -3 16 105
use FILL  FILL_2286
timestamp 1745462530
transform 1 0 1632 0 1 2170
box -8 -3 16 105
use FILL  FILL_2287
timestamp 1745462530
transform 1 0 1600 0 1 2170
box -8 -3 16 105
use FILL  FILL_2288
timestamp 1745462530
transform 1 0 1592 0 1 2170
box -8 -3 16 105
use FILL  FILL_2289
timestamp 1745462530
transform 1 0 1584 0 1 2170
box -8 -3 16 105
use FILL  FILL_2290
timestamp 1745462530
transform 1 0 1536 0 1 2170
box -8 -3 16 105
use FILL  FILL_2291
timestamp 1745462530
transform 1 0 1528 0 1 2170
box -8 -3 16 105
use FILL  FILL_2292
timestamp 1745462530
transform 1 0 1480 0 1 2170
box -8 -3 16 105
use FILL  FILL_2293
timestamp 1745462530
transform 1 0 1472 0 1 2170
box -8 -3 16 105
use FILL  FILL_2294
timestamp 1745462530
transform 1 0 1432 0 1 2170
box -8 -3 16 105
use FILL  FILL_2295
timestamp 1745462530
transform 1 0 1424 0 1 2170
box -8 -3 16 105
use FILL  FILL_2296
timestamp 1745462530
transform 1 0 1416 0 1 2170
box -8 -3 16 105
use FILL  FILL_2297
timestamp 1745462530
transform 1 0 1352 0 1 2170
box -8 -3 16 105
use FILL  FILL_2298
timestamp 1745462530
transform 1 0 1328 0 1 2170
box -8 -3 16 105
use FILL  FILL_2299
timestamp 1745462530
transform 1 0 1320 0 1 2170
box -8 -3 16 105
use FILL  FILL_2300
timestamp 1745462530
transform 1 0 1272 0 1 2170
box -8 -3 16 105
use FILL  FILL_2301
timestamp 1745462530
transform 1 0 1264 0 1 2170
box -8 -3 16 105
use FILL  FILL_2302
timestamp 1745462530
transform 1 0 1256 0 1 2170
box -8 -3 16 105
use FILL  FILL_2303
timestamp 1745462530
transform 1 0 1208 0 1 2170
box -8 -3 16 105
use FILL  FILL_2304
timestamp 1745462530
transform 1 0 1200 0 1 2170
box -8 -3 16 105
use FILL  FILL_2305
timestamp 1745462530
transform 1 0 1152 0 1 2170
box -8 -3 16 105
use FILL  FILL_2306
timestamp 1745462530
transform 1 0 1144 0 1 2170
box -8 -3 16 105
use FILL  FILL_2307
timestamp 1745462530
transform 1 0 1136 0 1 2170
box -8 -3 16 105
use FILL  FILL_2308
timestamp 1745462530
transform 1 0 1096 0 1 2170
box -8 -3 16 105
use FILL  FILL_2309
timestamp 1745462530
transform 1 0 1064 0 1 2170
box -8 -3 16 105
use FILL  FILL_2310
timestamp 1745462530
transform 1 0 1056 0 1 2170
box -8 -3 16 105
use FILL  FILL_2311
timestamp 1745462530
transform 1 0 1008 0 1 2170
box -8 -3 16 105
use FILL  FILL_2312
timestamp 1745462530
transform 1 0 1000 0 1 2170
box -8 -3 16 105
use FILL  FILL_2313
timestamp 1745462530
transform 1 0 944 0 1 2170
box -8 -3 16 105
use FILL  FILL_2314
timestamp 1745462530
transform 1 0 896 0 1 2170
box -8 -3 16 105
use FILL  FILL_2315
timestamp 1745462530
transform 1 0 888 0 1 2170
box -8 -3 16 105
use FILL  FILL_2316
timestamp 1745462530
transform 1 0 848 0 1 2170
box -8 -3 16 105
use FILL  FILL_2317
timestamp 1745462530
transform 1 0 800 0 1 2170
box -8 -3 16 105
use FILL  FILL_2318
timestamp 1745462530
transform 1 0 792 0 1 2170
box -8 -3 16 105
use FILL  FILL_2319
timestamp 1745462530
transform 1 0 784 0 1 2170
box -8 -3 16 105
use FILL  FILL_2320
timestamp 1745462530
transform 1 0 744 0 1 2170
box -8 -3 16 105
use FILL  FILL_2321
timestamp 1745462530
transform 1 0 696 0 1 2170
box -8 -3 16 105
use FILL  FILL_2322
timestamp 1745462530
transform 1 0 688 0 1 2170
box -8 -3 16 105
use FILL  FILL_2323
timestamp 1745462530
transform 1 0 648 0 1 2170
box -8 -3 16 105
use FILL  FILL_2324
timestamp 1745462530
transform 1 0 640 0 1 2170
box -8 -3 16 105
use FILL  FILL_2325
timestamp 1745462530
transform 1 0 592 0 1 2170
box -8 -3 16 105
use FILL  FILL_2326
timestamp 1745462530
transform 1 0 584 0 1 2170
box -8 -3 16 105
use FILL  FILL_2327
timestamp 1745462530
transform 1 0 552 0 1 2170
box -8 -3 16 105
use FILL  FILL_2328
timestamp 1745462530
transform 1 0 544 0 1 2170
box -8 -3 16 105
use FILL  FILL_2329
timestamp 1745462530
transform 1 0 496 0 1 2170
box -8 -3 16 105
use FILL  FILL_2330
timestamp 1745462530
transform 1 0 488 0 1 2170
box -8 -3 16 105
use FILL  FILL_2331
timestamp 1745462530
transform 1 0 384 0 1 2170
box -8 -3 16 105
use FILL  FILL_2332
timestamp 1745462530
transform 1 0 376 0 1 2170
box -8 -3 16 105
use FILL  FILL_2333
timestamp 1745462530
transform 1 0 352 0 1 2170
box -8 -3 16 105
use FILL  FILL_2334
timestamp 1745462530
transform 1 0 304 0 1 2170
box -8 -3 16 105
use FILL  FILL_2335
timestamp 1745462530
transform 1 0 296 0 1 2170
box -8 -3 16 105
use FILL  FILL_2336
timestamp 1745462530
transform 1 0 192 0 1 2170
box -8 -3 16 105
use FILL  FILL_2337
timestamp 1745462530
transform 1 0 184 0 1 2170
box -8 -3 16 105
use FILL  FILL_2338
timestamp 1745462530
transform 1 0 176 0 1 2170
box -8 -3 16 105
use FILL  FILL_2339
timestamp 1745462530
transform 1 0 72 0 1 2170
box -8 -3 16 105
use FILL  FILL_2340
timestamp 1745462530
transform 1 0 4080 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2341
timestamp 1745462530
transform 1 0 4032 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2342
timestamp 1745462530
transform 1 0 4024 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2343
timestamp 1745462530
transform 1 0 3984 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2344
timestamp 1745462530
transform 1 0 3952 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2345
timestamp 1745462530
transform 1 0 3944 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2346
timestamp 1745462530
transform 1 0 3896 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2347
timestamp 1745462530
transform 1 0 3856 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2348
timestamp 1745462530
transform 1 0 3808 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2349
timestamp 1745462530
transform 1 0 3800 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2350
timestamp 1745462530
transform 1 0 3696 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2351
timestamp 1745462530
transform 1 0 3592 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2352
timestamp 1745462530
transform 1 0 3584 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2353
timestamp 1745462530
transform 1 0 3576 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2354
timestamp 1745462530
transform 1 0 3528 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2355
timestamp 1745462530
transform 1 0 3520 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2356
timestamp 1745462530
transform 1 0 3488 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2357
timestamp 1745462530
transform 1 0 3480 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2358
timestamp 1745462530
transform 1 0 3472 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2359
timestamp 1745462530
transform 1 0 3424 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2360
timestamp 1745462530
transform 1 0 3416 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2361
timestamp 1745462530
transform 1 0 3408 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2362
timestamp 1745462530
transform 1 0 3400 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2363
timestamp 1745462530
transform 1 0 3352 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2364
timestamp 1745462530
transform 1 0 3344 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2365
timestamp 1745462530
transform 1 0 3336 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2366
timestamp 1745462530
transform 1 0 3288 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2367
timestamp 1745462530
transform 1 0 3280 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2368
timestamp 1745462530
transform 1 0 3272 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2369
timestamp 1745462530
transform 1 0 3240 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2370
timestamp 1745462530
transform 1 0 3232 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2371
timestamp 1745462530
transform 1 0 3160 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2372
timestamp 1745462530
transform 1 0 3152 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2373
timestamp 1745462530
transform 1 0 3144 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2374
timestamp 1745462530
transform 1 0 3104 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2375
timestamp 1745462530
transform 1 0 3096 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2376
timestamp 1745462530
transform 1 0 3088 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2377
timestamp 1745462530
transform 1 0 3048 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2378
timestamp 1745462530
transform 1 0 3040 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2379
timestamp 1745462530
transform 1 0 3032 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2380
timestamp 1745462530
transform 1 0 3024 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2381
timestamp 1745462530
transform 1 0 2976 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2382
timestamp 1745462530
transform 1 0 2968 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2383
timestamp 1745462530
transform 1 0 2960 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2384
timestamp 1745462530
transform 1 0 2952 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2385
timestamp 1745462530
transform 1 0 2912 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2386
timestamp 1745462530
transform 1 0 2888 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2387
timestamp 1745462530
transform 1 0 2880 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2388
timestamp 1745462530
transform 1 0 2872 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2389
timestamp 1745462530
transform 1 0 2864 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2390
timestamp 1745462530
transform 1 0 2816 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2391
timestamp 1745462530
transform 1 0 2808 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2392
timestamp 1745462530
transform 1 0 2800 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2393
timestamp 1745462530
transform 1 0 2776 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2394
timestamp 1745462530
transform 1 0 2768 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2395
timestamp 1745462530
transform 1 0 2728 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2396
timestamp 1745462530
transform 1 0 2720 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2397
timestamp 1745462530
transform 1 0 2712 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2398
timestamp 1745462530
transform 1 0 2672 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2399
timestamp 1745462530
transform 1 0 2664 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2400
timestamp 1745462530
transform 1 0 2616 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2401
timestamp 1745462530
transform 1 0 2608 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2402
timestamp 1745462530
transform 1 0 2600 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2403
timestamp 1745462530
transform 1 0 2568 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2404
timestamp 1745462530
transform 1 0 2528 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2405
timestamp 1745462530
transform 1 0 2520 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2406
timestamp 1745462530
transform 1 0 2512 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2407
timestamp 1745462530
transform 1 0 2456 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2408
timestamp 1745462530
transform 1 0 2448 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2409
timestamp 1745462530
transform 1 0 2400 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2410
timestamp 1745462530
transform 1 0 2344 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2411
timestamp 1745462530
transform 1 0 2312 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2412
timestamp 1745462530
transform 1 0 2272 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2413
timestamp 1745462530
transform 1 0 2264 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2414
timestamp 1745462530
transform 1 0 2224 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2415
timestamp 1745462530
transform 1 0 2216 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2416
timestamp 1745462530
transform 1 0 2176 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2417
timestamp 1745462530
transform 1 0 2168 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2418
timestamp 1745462530
transform 1 0 2128 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2419
timestamp 1745462530
transform 1 0 2120 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2420
timestamp 1745462530
transform 1 0 2080 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2421
timestamp 1745462530
transform 1 0 2072 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2422
timestamp 1745462530
transform 1 0 2024 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2423
timestamp 1745462530
transform 1 0 2016 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2424
timestamp 1745462530
transform 1 0 1896 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2425
timestamp 1745462530
transform 1 0 1888 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2426
timestamp 1745462530
transform 1 0 1832 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2427
timestamp 1745462530
transform 1 0 1824 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2428
timestamp 1745462530
transform 1 0 1776 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2429
timestamp 1745462530
transform 1 0 1768 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2430
timestamp 1745462530
transform 1 0 1736 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2431
timestamp 1745462530
transform 1 0 1632 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2432
timestamp 1745462530
transform 1 0 1528 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2433
timestamp 1745462530
transform 1 0 1520 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2434
timestamp 1745462530
transform 1 0 1480 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2435
timestamp 1745462530
transform 1 0 1472 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2436
timestamp 1745462530
transform 1 0 1440 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2437
timestamp 1745462530
transform 1 0 1432 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2438
timestamp 1745462530
transform 1 0 1400 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2439
timestamp 1745462530
transform 1 0 1368 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2440
timestamp 1745462530
transform 1 0 1240 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2441
timestamp 1745462530
transform 1 0 1232 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2442
timestamp 1745462530
transform 1 0 1184 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2443
timestamp 1745462530
transform 1 0 1176 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2444
timestamp 1745462530
transform 1 0 1168 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2445
timestamp 1745462530
transform 1 0 1120 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2446
timestamp 1745462530
transform 1 0 1072 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2447
timestamp 1745462530
transform 1 0 1064 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2448
timestamp 1745462530
transform 1 0 960 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2449
timestamp 1745462530
transform 1 0 928 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2450
timestamp 1745462530
transform 1 0 920 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2451
timestamp 1745462530
transform 1 0 872 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2452
timestamp 1745462530
transform 1 0 864 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2453
timestamp 1745462530
transform 1 0 824 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2454
timestamp 1745462530
transform 1 0 816 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2455
timestamp 1745462530
transform 1 0 768 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2456
timestamp 1745462530
transform 1 0 760 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2457
timestamp 1745462530
transform 1 0 720 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2458
timestamp 1745462530
transform 1 0 712 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2459
timestamp 1745462530
transform 1 0 672 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2460
timestamp 1745462530
transform 1 0 624 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2461
timestamp 1745462530
transform 1 0 616 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2462
timestamp 1745462530
transform 1 0 568 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2463
timestamp 1745462530
transform 1 0 560 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2464
timestamp 1745462530
transform 1 0 520 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2465
timestamp 1745462530
transform 1 0 512 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2466
timestamp 1745462530
transform 1 0 448 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2467
timestamp 1745462530
transform 1 0 440 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2468
timestamp 1745462530
transform 1 0 336 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2469
timestamp 1745462530
transform 1 0 328 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2470
timestamp 1745462530
transform 1 0 264 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2471
timestamp 1745462530
transform 1 0 240 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2472
timestamp 1745462530
transform 1 0 176 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2473
timestamp 1745462530
transform 1 0 72 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2474
timestamp 1745462530
transform 1 0 4368 0 1 1970
box -8 -3 16 105
use FILL  FILL_2475
timestamp 1745462530
transform 1 0 4360 0 1 1970
box -8 -3 16 105
use FILL  FILL_2476
timestamp 1745462530
transform 1 0 4352 0 1 1970
box -8 -3 16 105
use FILL  FILL_2477
timestamp 1745462530
transform 1 0 4344 0 1 1970
box -8 -3 16 105
use FILL  FILL_2478
timestamp 1745462530
transform 1 0 4336 0 1 1970
box -8 -3 16 105
use FILL  FILL_2479
timestamp 1745462530
transform 1 0 4272 0 1 1970
box -8 -3 16 105
use FILL  FILL_2480
timestamp 1745462530
transform 1 0 4264 0 1 1970
box -8 -3 16 105
use FILL  FILL_2481
timestamp 1745462530
transform 1 0 4256 0 1 1970
box -8 -3 16 105
use FILL  FILL_2482
timestamp 1745462530
transform 1 0 4248 0 1 1970
box -8 -3 16 105
use FILL  FILL_2483
timestamp 1745462530
transform 1 0 4184 0 1 1970
box -8 -3 16 105
use FILL  FILL_2484
timestamp 1745462530
transform 1 0 4176 0 1 1970
box -8 -3 16 105
use FILL  FILL_2485
timestamp 1745462530
transform 1 0 4168 0 1 1970
box -8 -3 16 105
use FILL  FILL_2486
timestamp 1745462530
transform 1 0 4104 0 1 1970
box -8 -3 16 105
use FILL  FILL_2487
timestamp 1745462530
transform 1 0 4096 0 1 1970
box -8 -3 16 105
use FILL  FILL_2488
timestamp 1745462530
transform 1 0 3992 0 1 1970
box -8 -3 16 105
use FILL  FILL_2489
timestamp 1745462530
transform 1 0 3984 0 1 1970
box -8 -3 16 105
use FILL  FILL_2490
timestamp 1745462530
transform 1 0 3976 0 1 1970
box -8 -3 16 105
use FILL  FILL_2491
timestamp 1745462530
transform 1 0 3928 0 1 1970
box -8 -3 16 105
use FILL  FILL_2492
timestamp 1745462530
transform 1 0 3920 0 1 1970
box -8 -3 16 105
use FILL  FILL_2493
timestamp 1745462530
transform 1 0 3912 0 1 1970
box -8 -3 16 105
use FILL  FILL_2494
timestamp 1745462530
transform 1 0 3888 0 1 1970
box -8 -3 16 105
use FILL  FILL_2495
timestamp 1745462530
transform 1 0 3880 0 1 1970
box -8 -3 16 105
use FILL  FILL_2496
timestamp 1745462530
transform 1 0 3832 0 1 1970
box -8 -3 16 105
use FILL  FILL_2497
timestamp 1745462530
transform 1 0 3824 0 1 1970
box -8 -3 16 105
use FILL  FILL_2498
timestamp 1745462530
transform 1 0 3816 0 1 1970
box -8 -3 16 105
use FILL  FILL_2499
timestamp 1745462530
transform 1 0 3808 0 1 1970
box -8 -3 16 105
use FILL  FILL_2500
timestamp 1745462530
transform 1 0 3760 0 1 1970
box -8 -3 16 105
use FILL  FILL_2501
timestamp 1745462530
transform 1 0 3752 0 1 1970
box -8 -3 16 105
use FILL  FILL_2502
timestamp 1745462530
transform 1 0 3728 0 1 1970
box -8 -3 16 105
use FILL  FILL_2503
timestamp 1745462530
transform 1 0 3720 0 1 1970
box -8 -3 16 105
use FILL  FILL_2504
timestamp 1745462530
transform 1 0 3712 0 1 1970
box -8 -3 16 105
use FILL  FILL_2505
timestamp 1745462530
transform 1 0 3664 0 1 1970
box -8 -3 16 105
use FILL  FILL_2506
timestamp 1745462530
transform 1 0 3656 0 1 1970
box -8 -3 16 105
use FILL  FILL_2507
timestamp 1745462530
transform 1 0 3632 0 1 1970
box -8 -3 16 105
use FILL  FILL_2508
timestamp 1745462530
transform 1 0 3624 0 1 1970
box -8 -3 16 105
use FILL  FILL_2509
timestamp 1745462530
transform 1 0 3616 0 1 1970
box -8 -3 16 105
use FILL  FILL_2510
timestamp 1745462530
transform 1 0 3608 0 1 1970
box -8 -3 16 105
use FILL  FILL_2511
timestamp 1745462530
transform 1 0 3560 0 1 1970
box -8 -3 16 105
use FILL  FILL_2512
timestamp 1745462530
transform 1 0 3552 0 1 1970
box -8 -3 16 105
use FILL  FILL_2513
timestamp 1745462530
transform 1 0 3544 0 1 1970
box -8 -3 16 105
use FILL  FILL_2514
timestamp 1745462530
transform 1 0 3536 0 1 1970
box -8 -3 16 105
use FILL  FILL_2515
timestamp 1745462530
transform 1 0 3496 0 1 1970
box -8 -3 16 105
use FILL  FILL_2516
timestamp 1745462530
transform 1 0 3488 0 1 1970
box -8 -3 16 105
use FILL  FILL_2517
timestamp 1745462530
transform 1 0 3480 0 1 1970
box -8 -3 16 105
use FILL  FILL_2518
timestamp 1745462530
transform 1 0 3472 0 1 1970
box -8 -3 16 105
use FILL  FILL_2519
timestamp 1745462530
transform 1 0 3432 0 1 1970
box -8 -3 16 105
use FILL  FILL_2520
timestamp 1745462530
transform 1 0 3424 0 1 1970
box -8 -3 16 105
use FILL  FILL_2521
timestamp 1745462530
transform 1 0 3416 0 1 1970
box -8 -3 16 105
use FILL  FILL_2522
timestamp 1745462530
transform 1 0 3408 0 1 1970
box -8 -3 16 105
use FILL  FILL_2523
timestamp 1745462530
transform 1 0 3400 0 1 1970
box -8 -3 16 105
use FILL  FILL_2524
timestamp 1745462530
transform 1 0 3352 0 1 1970
box -8 -3 16 105
use FILL  FILL_2525
timestamp 1745462530
transform 1 0 3344 0 1 1970
box -8 -3 16 105
use FILL  FILL_2526
timestamp 1745462530
transform 1 0 3336 0 1 1970
box -8 -3 16 105
use FILL  FILL_2527
timestamp 1745462530
transform 1 0 3328 0 1 1970
box -8 -3 16 105
use FILL  FILL_2528
timestamp 1745462530
transform 1 0 3288 0 1 1970
box -8 -3 16 105
use FILL  FILL_2529
timestamp 1745462530
transform 1 0 3256 0 1 1970
box -8 -3 16 105
use FILL  FILL_2530
timestamp 1745462530
transform 1 0 3248 0 1 1970
box -8 -3 16 105
use FILL  FILL_2531
timestamp 1745462530
transform 1 0 3240 0 1 1970
box -8 -3 16 105
use FILL  FILL_2532
timestamp 1745462530
transform 1 0 3192 0 1 1970
box -8 -3 16 105
use FILL  FILL_2533
timestamp 1745462530
transform 1 0 3184 0 1 1970
box -8 -3 16 105
use FILL  FILL_2534
timestamp 1745462530
transform 1 0 3176 0 1 1970
box -8 -3 16 105
use FILL  FILL_2535
timestamp 1745462530
transform 1 0 3168 0 1 1970
box -8 -3 16 105
use FILL  FILL_2536
timestamp 1745462530
transform 1 0 3136 0 1 1970
box -8 -3 16 105
use FILL  FILL_2537
timestamp 1745462530
transform 1 0 3104 0 1 1970
box -8 -3 16 105
use FILL  FILL_2538
timestamp 1745462530
transform 1 0 3096 0 1 1970
box -8 -3 16 105
use FILL  FILL_2539
timestamp 1745462530
transform 1 0 3088 0 1 1970
box -8 -3 16 105
use FILL  FILL_2540
timestamp 1745462530
transform 1 0 3048 0 1 1970
box -8 -3 16 105
use FILL  FILL_2541
timestamp 1745462530
transform 1 0 3040 0 1 1970
box -8 -3 16 105
use FILL  FILL_2542
timestamp 1745462530
transform 1 0 3032 0 1 1970
box -8 -3 16 105
use FILL  FILL_2543
timestamp 1745462530
transform 1 0 2984 0 1 1970
box -8 -3 16 105
use FILL  FILL_2544
timestamp 1745462530
transform 1 0 2976 0 1 1970
box -8 -3 16 105
use FILL  FILL_2545
timestamp 1745462530
transform 1 0 2968 0 1 1970
box -8 -3 16 105
use FILL  FILL_2546
timestamp 1745462530
transform 1 0 2920 0 1 1970
box -8 -3 16 105
use FILL  FILL_2547
timestamp 1745462530
transform 1 0 2912 0 1 1970
box -8 -3 16 105
use FILL  FILL_2548
timestamp 1745462530
transform 1 0 2904 0 1 1970
box -8 -3 16 105
use FILL  FILL_2549
timestamp 1745462530
transform 1 0 2800 0 1 1970
box -8 -3 16 105
use FILL  FILL_2550
timestamp 1745462530
transform 1 0 2768 0 1 1970
box -8 -3 16 105
use FILL  FILL_2551
timestamp 1745462530
transform 1 0 2760 0 1 1970
box -8 -3 16 105
use FILL  FILL_2552
timestamp 1745462530
transform 1 0 2752 0 1 1970
box -8 -3 16 105
use FILL  FILL_2553
timestamp 1745462530
transform 1 0 2712 0 1 1970
box -8 -3 16 105
use FILL  FILL_2554
timestamp 1745462530
transform 1 0 2704 0 1 1970
box -8 -3 16 105
use FILL  FILL_2555
timestamp 1745462530
transform 1 0 2600 0 1 1970
box -8 -3 16 105
use FILL  FILL_2556
timestamp 1745462530
transform 1 0 2544 0 1 1970
box -8 -3 16 105
use FILL  FILL_2557
timestamp 1745462530
transform 1 0 2536 0 1 1970
box -8 -3 16 105
use FILL  FILL_2558
timestamp 1745462530
transform 1 0 2504 0 1 1970
box -8 -3 16 105
use FILL  FILL_2559
timestamp 1745462530
transform 1 0 2448 0 1 1970
box -8 -3 16 105
use FILL  FILL_2560
timestamp 1745462530
transform 1 0 2440 0 1 1970
box -8 -3 16 105
use FILL  FILL_2561
timestamp 1745462530
transform 1 0 2384 0 1 1970
box -8 -3 16 105
use FILL  FILL_2562
timestamp 1745462530
transform 1 0 2352 0 1 1970
box -8 -3 16 105
use FILL  FILL_2563
timestamp 1745462530
transform 1 0 2296 0 1 1970
box -8 -3 16 105
use FILL  FILL_2564
timestamp 1745462530
transform 1 0 2288 0 1 1970
box -8 -3 16 105
use FILL  FILL_2565
timestamp 1745462530
transform 1 0 2240 0 1 1970
box -8 -3 16 105
use FILL  FILL_2566
timestamp 1745462530
transform 1 0 2232 0 1 1970
box -8 -3 16 105
use FILL  FILL_2567
timestamp 1745462530
transform 1 0 2176 0 1 1970
box -8 -3 16 105
use FILL  FILL_2568
timestamp 1745462530
transform 1 0 2168 0 1 1970
box -8 -3 16 105
use FILL  FILL_2569
timestamp 1745462530
transform 1 0 2064 0 1 1970
box -8 -3 16 105
use FILL  FILL_2570
timestamp 1745462530
transform 1 0 1960 0 1 1970
box -8 -3 16 105
use FILL  FILL_2571
timestamp 1745462530
transform 1 0 1952 0 1 1970
box -8 -3 16 105
use FILL  FILL_2572
timestamp 1745462530
transform 1 0 1904 0 1 1970
box -8 -3 16 105
use FILL  FILL_2573
timestamp 1745462530
transform 1 0 1896 0 1 1970
box -8 -3 16 105
use FILL  FILL_2574
timestamp 1745462530
transform 1 0 1872 0 1 1970
box -8 -3 16 105
use FILL  FILL_2575
timestamp 1745462530
transform 1 0 1864 0 1 1970
box -8 -3 16 105
use FILL  FILL_2576
timestamp 1745462530
transform 1 0 1816 0 1 1970
box -8 -3 16 105
use FILL  FILL_2577
timestamp 1745462530
transform 1 0 1808 0 1 1970
box -8 -3 16 105
use FILL  FILL_2578
timestamp 1745462530
transform 1 0 1760 0 1 1970
box -8 -3 16 105
use FILL  FILL_2579
timestamp 1745462530
transform 1 0 1656 0 1 1970
box -8 -3 16 105
use FILL  FILL_2580
timestamp 1745462530
transform 1 0 1632 0 1 1970
box -8 -3 16 105
use FILL  FILL_2581
timestamp 1745462530
transform 1 0 1624 0 1 1970
box -8 -3 16 105
use FILL  FILL_2582
timestamp 1745462530
transform 1 0 1616 0 1 1970
box -8 -3 16 105
use FILL  FILL_2583
timestamp 1745462530
transform 1 0 1568 0 1 1970
box -8 -3 16 105
use FILL  FILL_2584
timestamp 1745462530
transform 1 0 1560 0 1 1970
box -8 -3 16 105
use FILL  FILL_2585
timestamp 1745462530
transform 1 0 1552 0 1 1970
box -8 -3 16 105
use FILL  FILL_2586
timestamp 1745462530
transform 1 0 1480 0 1 1970
box -8 -3 16 105
use FILL  FILL_2587
timestamp 1745462530
transform 1 0 1472 0 1 1970
box -8 -3 16 105
use FILL  FILL_2588
timestamp 1745462530
transform 1 0 1464 0 1 1970
box -8 -3 16 105
use FILL  FILL_2589
timestamp 1745462530
transform 1 0 1456 0 1 1970
box -8 -3 16 105
use FILL  FILL_2590
timestamp 1745462530
transform 1 0 1408 0 1 1970
box -8 -3 16 105
use FILL  FILL_2591
timestamp 1745462530
transform 1 0 1400 0 1 1970
box -8 -3 16 105
use FILL  FILL_2592
timestamp 1745462530
transform 1 0 1392 0 1 1970
box -8 -3 16 105
use FILL  FILL_2593
timestamp 1745462530
transform 1 0 1272 0 1 1970
box -8 -3 16 105
use FILL  FILL_2594
timestamp 1745462530
transform 1 0 1264 0 1 1970
box -8 -3 16 105
use FILL  FILL_2595
timestamp 1745462530
transform 1 0 1256 0 1 1970
box -8 -3 16 105
use FILL  FILL_2596
timestamp 1745462530
transform 1 0 1208 0 1 1970
box -8 -3 16 105
use FILL  FILL_2597
timestamp 1745462530
transform 1 0 1200 0 1 1970
box -8 -3 16 105
use FILL  FILL_2598
timestamp 1745462530
transform 1 0 1192 0 1 1970
box -8 -3 16 105
use FILL  FILL_2599
timestamp 1745462530
transform 1 0 1088 0 1 1970
box -8 -3 16 105
use FILL  FILL_2600
timestamp 1745462530
transform 1 0 1080 0 1 1970
box -8 -3 16 105
use FILL  FILL_2601
timestamp 1745462530
transform 1 0 1032 0 1 1970
box -8 -3 16 105
use FILL  FILL_2602
timestamp 1745462530
transform 1 0 1024 0 1 1970
box -8 -3 16 105
use FILL  FILL_2603
timestamp 1745462530
transform 1 0 1016 0 1 1970
box -8 -3 16 105
use FILL  FILL_2604
timestamp 1745462530
transform 1 0 968 0 1 1970
box -8 -3 16 105
use FILL  FILL_2605
timestamp 1745462530
transform 1 0 920 0 1 1970
box -8 -3 16 105
use FILL  FILL_2606
timestamp 1745462530
transform 1 0 912 0 1 1970
box -8 -3 16 105
use FILL  FILL_2607
timestamp 1745462530
transform 1 0 840 0 1 1970
box -8 -3 16 105
use FILL  FILL_2608
timestamp 1745462530
transform 1 0 832 0 1 1970
box -8 -3 16 105
use FILL  FILL_2609
timestamp 1745462530
transform 1 0 824 0 1 1970
box -8 -3 16 105
use FILL  FILL_2610
timestamp 1745462530
transform 1 0 816 0 1 1970
box -8 -3 16 105
use FILL  FILL_2611
timestamp 1745462530
transform 1 0 768 0 1 1970
box -8 -3 16 105
use FILL  FILL_2612
timestamp 1745462530
transform 1 0 760 0 1 1970
box -8 -3 16 105
use FILL  FILL_2613
timestamp 1745462530
transform 1 0 752 0 1 1970
box -8 -3 16 105
use FILL  FILL_2614
timestamp 1745462530
transform 1 0 704 0 1 1970
box -8 -3 16 105
use FILL  FILL_2615
timestamp 1745462530
transform 1 0 696 0 1 1970
box -8 -3 16 105
use FILL  FILL_2616
timestamp 1745462530
transform 1 0 688 0 1 1970
box -8 -3 16 105
use FILL  FILL_2617
timestamp 1745462530
transform 1 0 624 0 1 1970
box -8 -3 16 105
use FILL  FILL_2618
timestamp 1745462530
transform 1 0 616 0 1 1970
box -8 -3 16 105
use FILL  FILL_2619
timestamp 1745462530
transform 1 0 568 0 1 1970
box -8 -3 16 105
use FILL  FILL_2620
timestamp 1745462530
transform 1 0 560 0 1 1970
box -8 -3 16 105
use FILL  FILL_2621
timestamp 1745462530
transform 1 0 400 0 1 1970
box -8 -3 16 105
use FILL  FILL_2622
timestamp 1745462530
transform 1 0 336 0 1 1970
box -8 -3 16 105
use FILL  FILL_2623
timestamp 1745462530
transform 1 0 232 0 1 1970
box -8 -3 16 105
use FILL  FILL_2624
timestamp 1745462530
transform 1 0 168 0 1 1970
box -8 -3 16 105
use FILL  FILL_2625
timestamp 1745462530
transform 1 0 4256 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2626
timestamp 1745462530
transform 1 0 4248 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2627
timestamp 1745462530
transform 1 0 4160 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2628
timestamp 1745462530
transform 1 0 4152 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2629
timestamp 1745462530
transform 1 0 4144 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2630
timestamp 1745462530
transform 1 0 4080 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2631
timestamp 1745462530
transform 1 0 4032 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2632
timestamp 1745462530
transform 1 0 3992 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2633
timestamp 1745462530
transform 1 0 3952 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2634
timestamp 1745462530
transform 1 0 3944 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2635
timestamp 1745462530
transform 1 0 3896 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2636
timestamp 1745462530
transform 1 0 3864 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2637
timestamp 1745462530
transform 1 0 3856 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2638
timestamp 1745462530
transform 1 0 3792 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2639
timestamp 1745462530
transform 1 0 3784 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2640
timestamp 1745462530
transform 1 0 3776 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2641
timestamp 1745462530
transform 1 0 3728 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2642
timestamp 1745462530
transform 1 0 3696 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2643
timestamp 1745462530
transform 1 0 3688 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2644
timestamp 1745462530
transform 1 0 3680 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2645
timestamp 1745462530
transform 1 0 3632 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2646
timestamp 1745462530
transform 1 0 3624 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2647
timestamp 1745462530
transform 1 0 3616 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2648
timestamp 1745462530
transform 1 0 3568 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2649
timestamp 1745462530
transform 1 0 3560 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2650
timestamp 1745462530
transform 1 0 3552 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2651
timestamp 1745462530
transform 1 0 3504 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2652
timestamp 1745462530
transform 1 0 3496 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2653
timestamp 1745462530
transform 1 0 3488 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2654
timestamp 1745462530
transform 1 0 3440 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2655
timestamp 1745462530
transform 1 0 3432 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2656
timestamp 1745462530
transform 1 0 3424 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2657
timestamp 1745462530
transform 1 0 3384 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2658
timestamp 1745462530
transform 1 0 3376 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2659
timestamp 1745462530
transform 1 0 3272 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2660
timestamp 1745462530
transform 1 0 3240 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2661
timestamp 1745462530
transform 1 0 3232 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2662
timestamp 1745462530
transform 1 0 3184 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2663
timestamp 1745462530
transform 1 0 3176 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2664
timestamp 1745462530
transform 1 0 3168 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2665
timestamp 1745462530
transform 1 0 3120 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2666
timestamp 1745462530
transform 1 0 3112 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2667
timestamp 1745462530
transform 1 0 3104 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2668
timestamp 1745462530
transform 1 0 3072 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2669
timestamp 1745462530
transform 1 0 3064 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2670
timestamp 1745462530
transform 1 0 3016 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2671
timestamp 1745462530
transform 1 0 3008 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2672
timestamp 1745462530
transform 1 0 3000 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2673
timestamp 1745462530
transform 1 0 2992 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2674
timestamp 1745462530
transform 1 0 2944 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2675
timestamp 1745462530
transform 1 0 2936 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2676
timestamp 1745462530
transform 1 0 2832 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2677
timestamp 1745462530
transform 1 0 2728 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2678
timestamp 1745462530
transform 1 0 2704 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2679
timestamp 1745462530
transform 1 0 2696 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2680
timestamp 1745462530
transform 1 0 2648 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2681
timestamp 1745462530
transform 1 0 2640 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2682
timestamp 1745462530
transform 1 0 2536 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2683
timestamp 1745462530
transform 1 0 2528 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2684
timestamp 1745462530
transform 1 0 2480 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2685
timestamp 1745462530
transform 1 0 2472 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2686
timestamp 1745462530
transform 1 0 2464 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2687
timestamp 1745462530
transform 1 0 2432 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2688
timestamp 1745462530
transform 1 0 2424 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2689
timestamp 1745462530
transform 1 0 2384 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2690
timestamp 1745462530
transform 1 0 2376 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2691
timestamp 1745462530
transform 1 0 2368 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2692
timestamp 1745462530
transform 1 0 2336 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2693
timestamp 1745462530
transform 1 0 2328 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2694
timestamp 1745462530
transform 1 0 2320 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2695
timestamp 1745462530
transform 1 0 2280 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2696
timestamp 1745462530
transform 1 0 2272 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2697
timestamp 1745462530
transform 1 0 2216 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2698
timestamp 1745462530
transform 1 0 2208 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2699
timestamp 1745462530
transform 1 0 2176 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2700
timestamp 1745462530
transform 1 0 2168 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2701
timestamp 1745462530
transform 1 0 2160 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2702
timestamp 1745462530
transform 1 0 2120 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2703
timestamp 1745462530
transform 1 0 2112 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2704
timestamp 1745462530
transform 1 0 2080 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2705
timestamp 1745462530
transform 1 0 2048 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2706
timestamp 1745462530
transform 1 0 2040 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2707
timestamp 1745462530
transform 1 0 2032 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2708
timestamp 1745462530
transform 1 0 2024 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2709
timestamp 1745462530
transform 1 0 1976 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2710
timestamp 1745462530
transform 1 0 1968 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2711
timestamp 1745462530
transform 1 0 1864 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2712
timestamp 1745462530
transform 1 0 1840 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2713
timestamp 1745462530
transform 1 0 1832 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2714
timestamp 1745462530
transform 1 0 1824 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2715
timestamp 1745462530
transform 1 0 1776 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2716
timestamp 1745462530
transform 1 0 1768 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2717
timestamp 1745462530
transform 1 0 1760 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2718
timestamp 1745462530
transform 1 0 1752 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2719
timestamp 1745462530
transform 1 0 1704 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2720
timestamp 1745462530
transform 1 0 1696 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2721
timestamp 1745462530
transform 1 0 1688 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2722
timestamp 1745462530
transform 1 0 1680 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2723
timestamp 1745462530
transform 1 0 1672 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2724
timestamp 1745462530
transform 1 0 1624 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2725
timestamp 1745462530
transform 1 0 1616 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2726
timestamp 1745462530
transform 1 0 1608 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2727
timestamp 1745462530
transform 1 0 1600 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2728
timestamp 1745462530
transform 1 0 1592 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2729
timestamp 1745462530
transform 1 0 1544 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2730
timestamp 1745462530
transform 1 0 1536 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2731
timestamp 1745462530
transform 1 0 1528 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2732
timestamp 1745462530
transform 1 0 1520 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2733
timestamp 1745462530
transform 1 0 1472 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2734
timestamp 1745462530
transform 1 0 1464 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2735
timestamp 1745462530
transform 1 0 1360 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2736
timestamp 1745462530
transform 1 0 1352 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2737
timestamp 1745462530
transform 1 0 1344 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2738
timestamp 1745462530
transform 1 0 1296 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2739
timestamp 1745462530
transform 1 0 1288 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2740
timestamp 1745462530
transform 1 0 1280 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2741
timestamp 1745462530
transform 1 0 1272 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2742
timestamp 1745462530
transform 1 0 1264 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2743
timestamp 1745462530
transform 1 0 1216 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2744
timestamp 1745462530
transform 1 0 1208 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2745
timestamp 1745462530
transform 1 0 1200 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2746
timestamp 1745462530
transform 1 0 1192 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2747
timestamp 1745462530
transform 1 0 1144 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2748
timestamp 1745462530
transform 1 0 1136 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2749
timestamp 1745462530
transform 1 0 1112 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2750
timestamp 1745462530
transform 1 0 1080 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2751
timestamp 1745462530
transform 1 0 1072 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2752
timestamp 1745462530
transform 1 0 1064 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2753
timestamp 1745462530
transform 1 0 1056 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2754
timestamp 1745462530
transform 1 0 1024 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2755
timestamp 1745462530
transform 1 0 1016 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2756
timestamp 1745462530
transform 1 0 1008 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2757
timestamp 1745462530
transform 1 0 968 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2758
timestamp 1745462530
transform 1 0 960 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2759
timestamp 1745462530
transform 1 0 952 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2760
timestamp 1745462530
transform 1 0 944 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2761
timestamp 1745462530
transform 1 0 896 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2762
timestamp 1745462530
transform 1 0 888 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2763
timestamp 1745462530
transform 1 0 880 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2764
timestamp 1745462530
transform 1 0 872 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2765
timestamp 1745462530
transform 1 0 824 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2766
timestamp 1745462530
transform 1 0 816 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2767
timestamp 1745462530
transform 1 0 808 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2768
timestamp 1745462530
transform 1 0 760 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2769
timestamp 1745462530
transform 1 0 752 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2770
timestamp 1745462530
transform 1 0 744 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2771
timestamp 1745462530
transform 1 0 736 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2772
timestamp 1745462530
transform 1 0 696 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2773
timestamp 1745462530
transform 1 0 688 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2774
timestamp 1745462530
transform 1 0 680 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2775
timestamp 1745462530
transform 1 0 632 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2776
timestamp 1745462530
transform 1 0 624 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2777
timestamp 1745462530
transform 1 0 616 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2778
timestamp 1745462530
transform 1 0 512 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2779
timestamp 1745462530
transform 1 0 504 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2780
timestamp 1745462530
transform 1 0 464 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2781
timestamp 1745462530
transform 1 0 440 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2782
timestamp 1745462530
transform 1 0 432 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2783
timestamp 1745462530
transform 1 0 328 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2784
timestamp 1745462530
transform 1 0 304 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2785
timestamp 1745462530
transform 1 0 200 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2786
timestamp 1745462530
transform 1 0 176 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2787
timestamp 1745462530
transform 1 0 72 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2788
timestamp 1745462530
transform 1 0 4368 0 1 1770
box -8 -3 16 105
use FILL  FILL_2789
timestamp 1745462530
transform 1 0 4248 0 1 1770
box -8 -3 16 105
use FILL  FILL_2790
timestamp 1745462530
transform 1 0 4200 0 1 1770
box -8 -3 16 105
use FILL  FILL_2791
timestamp 1745462530
transform 1 0 4160 0 1 1770
box -8 -3 16 105
use FILL  FILL_2792
timestamp 1745462530
transform 1 0 4056 0 1 1770
box -8 -3 16 105
use FILL  FILL_2793
timestamp 1745462530
transform 1 0 4048 0 1 1770
box -8 -3 16 105
use FILL  FILL_2794
timestamp 1745462530
transform 1 0 3944 0 1 1770
box -8 -3 16 105
use FILL  FILL_2795
timestamp 1745462530
transform 1 0 3936 0 1 1770
box -8 -3 16 105
use FILL  FILL_2796
timestamp 1745462530
transform 1 0 3912 0 1 1770
box -8 -3 16 105
use FILL  FILL_2797
timestamp 1745462530
transform 1 0 3864 0 1 1770
box -8 -3 16 105
use FILL  FILL_2798
timestamp 1745462530
transform 1 0 3856 0 1 1770
box -8 -3 16 105
use FILL  FILL_2799
timestamp 1745462530
transform 1 0 3808 0 1 1770
box -8 -3 16 105
use FILL  FILL_2800
timestamp 1745462530
transform 1 0 3800 0 1 1770
box -8 -3 16 105
use FILL  FILL_2801
timestamp 1745462530
transform 1 0 3792 0 1 1770
box -8 -3 16 105
use FILL  FILL_2802
timestamp 1745462530
transform 1 0 3744 0 1 1770
box -8 -3 16 105
use FILL  FILL_2803
timestamp 1745462530
transform 1 0 3736 0 1 1770
box -8 -3 16 105
use FILL  FILL_2804
timestamp 1745462530
transform 1 0 3728 0 1 1770
box -8 -3 16 105
use FILL  FILL_2805
timestamp 1745462530
transform 1 0 3720 0 1 1770
box -8 -3 16 105
use FILL  FILL_2806
timestamp 1745462530
transform 1 0 3712 0 1 1770
box -8 -3 16 105
use FILL  FILL_2807
timestamp 1745462530
transform 1 0 3664 0 1 1770
box -8 -3 16 105
use FILL  FILL_2808
timestamp 1745462530
transform 1 0 3656 0 1 1770
box -8 -3 16 105
use FILL  FILL_2809
timestamp 1745462530
transform 1 0 3648 0 1 1770
box -8 -3 16 105
use FILL  FILL_2810
timestamp 1745462530
transform 1 0 3528 0 1 1770
box -8 -3 16 105
use FILL  FILL_2811
timestamp 1745462530
transform 1 0 3520 0 1 1770
box -8 -3 16 105
use FILL  FILL_2812
timestamp 1745462530
transform 1 0 3512 0 1 1770
box -8 -3 16 105
use FILL  FILL_2813
timestamp 1745462530
transform 1 0 3504 0 1 1770
box -8 -3 16 105
use FILL  FILL_2814
timestamp 1745462530
transform 1 0 3456 0 1 1770
box -8 -3 16 105
use FILL  FILL_2815
timestamp 1745462530
transform 1 0 3448 0 1 1770
box -8 -3 16 105
use FILL  FILL_2816
timestamp 1745462530
transform 1 0 3344 0 1 1770
box -8 -3 16 105
use FILL  FILL_2817
timestamp 1745462530
transform 1 0 3320 0 1 1770
box -8 -3 16 105
use FILL  FILL_2818
timestamp 1745462530
transform 1 0 3312 0 1 1770
box -8 -3 16 105
use FILL  FILL_2819
timestamp 1745462530
transform 1 0 3304 0 1 1770
box -8 -3 16 105
use FILL  FILL_2820
timestamp 1745462530
transform 1 0 3256 0 1 1770
box -8 -3 16 105
use FILL  FILL_2821
timestamp 1745462530
transform 1 0 3248 0 1 1770
box -8 -3 16 105
use FILL  FILL_2822
timestamp 1745462530
transform 1 0 3240 0 1 1770
box -8 -3 16 105
use FILL  FILL_2823
timestamp 1745462530
transform 1 0 3232 0 1 1770
box -8 -3 16 105
use FILL  FILL_2824
timestamp 1745462530
transform 1 0 3200 0 1 1770
box -8 -3 16 105
use FILL  FILL_2825
timestamp 1745462530
transform 1 0 3192 0 1 1770
box -8 -3 16 105
use FILL  FILL_2826
timestamp 1745462530
transform 1 0 3160 0 1 1770
box -8 -3 16 105
use FILL  FILL_2827
timestamp 1745462530
transform 1 0 3152 0 1 1770
box -8 -3 16 105
use FILL  FILL_2828
timestamp 1745462530
transform 1 0 3144 0 1 1770
box -8 -3 16 105
use FILL  FILL_2829
timestamp 1745462530
transform 1 0 3040 0 1 1770
box -8 -3 16 105
use FILL  FILL_2830
timestamp 1745462530
transform 1 0 3016 0 1 1770
box -8 -3 16 105
use FILL  FILL_2831
timestamp 1745462530
transform 1 0 3008 0 1 1770
box -8 -3 16 105
use FILL  FILL_2832
timestamp 1745462530
transform 1 0 3000 0 1 1770
box -8 -3 16 105
use FILL  FILL_2833
timestamp 1745462530
transform 1 0 2952 0 1 1770
box -8 -3 16 105
use FILL  FILL_2834
timestamp 1745462530
transform 1 0 2944 0 1 1770
box -8 -3 16 105
use FILL  FILL_2835
timestamp 1745462530
transform 1 0 2936 0 1 1770
box -8 -3 16 105
use FILL  FILL_2836
timestamp 1745462530
transform 1 0 2912 0 1 1770
box -8 -3 16 105
use FILL  FILL_2837
timestamp 1745462530
transform 1 0 2904 0 1 1770
box -8 -3 16 105
use FILL  FILL_2838
timestamp 1745462530
transform 1 0 2896 0 1 1770
box -8 -3 16 105
use FILL  FILL_2839
timestamp 1745462530
transform 1 0 2848 0 1 1770
box -8 -3 16 105
use FILL  FILL_2840
timestamp 1745462530
transform 1 0 2840 0 1 1770
box -8 -3 16 105
use FILL  FILL_2841
timestamp 1745462530
transform 1 0 2832 0 1 1770
box -8 -3 16 105
use FILL  FILL_2842
timestamp 1745462530
transform 1 0 2808 0 1 1770
box -8 -3 16 105
use FILL  FILL_2843
timestamp 1745462530
transform 1 0 2800 0 1 1770
box -8 -3 16 105
use FILL  FILL_2844
timestamp 1745462530
transform 1 0 2752 0 1 1770
box -8 -3 16 105
use FILL  FILL_2845
timestamp 1745462530
transform 1 0 2744 0 1 1770
box -8 -3 16 105
use FILL  FILL_2846
timestamp 1745462530
transform 1 0 2736 0 1 1770
box -8 -3 16 105
use FILL  FILL_2847
timestamp 1745462530
transform 1 0 2728 0 1 1770
box -8 -3 16 105
use FILL  FILL_2848
timestamp 1745462530
transform 1 0 2680 0 1 1770
box -8 -3 16 105
use FILL  FILL_2849
timestamp 1745462530
transform 1 0 2672 0 1 1770
box -8 -3 16 105
use FILL  FILL_2850
timestamp 1745462530
transform 1 0 2664 0 1 1770
box -8 -3 16 105
use FILL  FILL_2851
timestamp 1745462530
transform 1 0 2640 0 1 1770
box -8 -3 16 105
use FILL  FILL_2852
timestamp 1745462530
transform 1 0 2632 0 1 1770
box -8 -3 16 105
use FILL  FILL_2853
timestamp 1745462530
transform 1 0 2624 0 1 1770
box -8 -3 16 105
use FILL  FILL_2854
timestamp 1745462530
transform 1 0 2520 0 1 1770
box -8 -3 16 105
use FILL  FILL_2855
timestamp 1745462530
transform 1 0 2512 0 1 1770
box -8 -3 16 105
use FILL  FILL_2856
timestamp 1745462530
transform 1 0 2504 0 1 1770
box -8 -3 16 105
use FILL  FILL_2857
timestamp 1745462530
transform 1 0 2496 0 1 1770
box -8 -3 16 105
use FILL  FILL_2858
timestamp 1745462530
transform 1 0 2456 0 1 1770
box -8 -3 16 105
use FILL  FILL_2859
timestamp 1745462530
transform 1 0 2448 0 1 1770
box -8 -3 16 105
use FILL  FILL_2860
timestamp 1745462530
transform 1 0 2440 0 1 1770
box -8 -3 16 105
use FILL  FILL_2861
timestamp 1745462530
transform 1 0 2408 0 1 1770
box -8 -3 16 105
use FILL  FILL_2862
timestamp 1745462530
transform 1 0 2400 0 1 1770
box -8 -3 16 105
use FILL  FILL_2863
timestamp 1745462530
transform 1 0 2392 0 1 1770
box -8 -3 16 105
use FILL  FILL_2864
timestamp 1745462530
transform 1 0 2352 0 1 1770
box -8 -3 16 105
use FILL  FILL_2865
timestamp 1745462530
transform 1 0 2344 0 1 1770
box -8 -3 16 105
use FILL  FILL_2866
timestamp 1745462530
transform 1 0 2336 0 1 1770
box -8 -3 16 105
use FILL  FILL_2867
timestamp 1745462530
transform 1 0 2328 0 1 1770
box -8 -3 16 105
use FILL  FILL_2868
timestamp 1745462530
transform 1 0 2280 0 1 1770
box -8 -3 16 105
use FILL  FILL_2869
timestamp 1745462530
transform 1 0 2272 0 1 1770
box -8 -3 16 105
use FILL  FILL_2870
timestamp 1745462530
transform 1 0 2240 0 1 1770
box -8 -3 16 105
use FILL  FILL_2871
timestamp 1745462530
transform 1 0 2232 0 1 1770
box -8 -3 16 105
use FILL  FILL_2872
timestamp 1745462530
transform 1 0 2200 0 1 1770
box -8 -3 16 105
use FILL  FILL_2873
timestamp 1745462530
transform 1 0 2192 0 1 1770
box -8 -3 16 105
use FILL  FILL_2874
timestamp 1745462530
transform 1 0 2184 0 1 1770
box -8 -3 16 105
use FILL  FILL_2875
timestamp 1745462530
transform 1 0 2152 0 1 1770
box -8 -3 16 105
use FILL  FILL_2876
timestamp 1745462530
transform 1 0 2120 0 1 1770
box -8 -3 16 105
use FILL  FILL_2877
timestamp 1745462530
transform 1 0 2112 0 1 1770
box -8 -3 16 105
use FILL  FILL_2878
timestamp 1745462530
transform 1 0 2056 0 1 1770
box -8 -3 16 105
use FILL  FILL_2879
timestamp 1745462530
transform 1 0 2048 0 1 1770
box -8 -3 16 105
use FILL  FILL_2880
timestamp 1745462530
transform 1 0 2040 0 1 1770
box -8 -3 16 105
use FILL  FILL_2881
timestamp 1745462530
transform 1 0 2000 0 1 1770
box -8 -3 16 105
use FILL  FILL_2882
timestamp 1745462530
transform 1 0 1992 0 1 1770
box -8 -3 16 105
use FILL  FILL_2883
timestamp 1745462530
transform 1 0 1984 0 1 1770
box -8 -3 16 105
use FILL  FILL_2884
timestamp 1745462530
transform 1 0 1952 0 1 1770
box -8 -3 16 105
use FILL  FILL_2885
timestamp 1745462530
transform 1 0 1912 0 1 1770
box -8 -3 16 105
use FILL  FILL_2886
timestamp 1745462530
transform 1 0 1904 0 1 1770
box -8 -3 16 105
use FILL  FILL_2887
timestamp 1745462530
transform 1 0 1896 0 1 1770
box -8 -3 16 105
use FILL  FILL_2888
timestamp 1745462530
transform 1 0 1888 0 1 1770
box -8 -3 16 105
use FILL  FILL_2889
timestamp 1745462530
transform 1 0 1856 0 1 1770
box -8 -3 16 105
use FILL  FILL_2890
timestamp 1745462530
transform 1 0 1832 0 1 1770
box -8 -3 16 105
use FILL  FILL_2891
timestamp 1745462530
transform 1 0 1824 0 1 1770
box -8 -3 16 105
use FILL  FILL_2892
timestamp 1745462530
transform 1 0 1816 0 1 1770
box -8 -3 16 105
use FILL  FILL_2893
timestamp 1745462530
transform 1 0 1712 0 1 1770
box -8 -3 16 105
use FILL  FILL_2894
timestamp 1745462530
transform 1 0 1704 0 1 1770
box -8 -3 16 105
use FILL  FILL_2895
timestamp 1745462530
transform 1 0 1696 0 1 1770
box -8 -3 16 105
use FILL  FILL_2896
timestamp 1745462530
transform 1 0 1648 0 1 1770
box -8 -3 16 105
use FILL  FILL_2897
timestamp 1745462530
transform 1 0 1640 0 1 1770
box -8 -3 16 105
use FILL  FILL_2898
timestamp 1745462530
transform 1 0 1632 0 1 1770
box -8 -3 16 105
use FILL  FILL_2899
timestamp 1745462530
transform 1 0 1512 0 1 1770
box -8 -3 16 105
use FILL  FILL_2900
timestamp 1745462530
transform 1 0 1504 0 1 1770
box -8 -3 16 105
use FILL  FILL_2901
timestamp 1745462530
transform 1 0 1496 0 1 1770
box -8 -3 16 105
use FILL  FILL_2902
timestamp 1745462530
transform 1 0 1488 0 1 1770
box -8 -3 16 105
use FILL  FILL_2903
timestamp 1745462530
transform 1 0 1440 0 1 1770
box -8 -3 16 105
use FILL  FILL_2904
timestamp 1745462530
transform 1 0 1432 0 1 1770
box -8 -3 16 105
use FILL  FILL_2905
timestamp 1745462530
transform 1 0 1424 0 1 1770
box -8 -3 16 105
use FILL  FILL_2906
timestamp 1745462530
transform 1 0 1400 0 1 1770
box -8 -3 16 105
use FILL  FILL_2907
timestamp 1745462530
transform 1 0 1392 0 1 1770
box -8 -3 16 105
use FILL  FILL_2908
timestamp 1745462530
transform 1 0 1384 0 1 1770
box -8 -3 16 105
use FILL  FILL_2909
timestamp 1745462530
transform 1 0 1336 0 1 1770
box -8 -3 16 105
use FILL  FILL_2910
timestamp 1745462530
transform 1 0 1328 0 1 1770
box -8 -3 16 105
use FILL  FILL_2911
timestamp 1745462530
transform 1 0 1320 0 1 1770
box -8 -3 16 105
use FILL  FILL_2912
timestamp 1745462530
transform 1 0 1216 0 1 1770
box -8 -3 16 105
use FILL  FILL_2913
timestamp 1745462530
transform 1 0 1192 0 1 1770
box -8 -3 16 105
use FILL  FILL_2914
timestamp 1745462530
transform 1 0 1184 0 1 1770
box -8 -3 16 105
use FILL  FILL_2915
timestamp 1745462530
transform 1 0 1144 0 1 1770
box -8 -3 16 105
use FILL  FILL_2916
timestamp 1745462530
transform 1 0 1136 0 1 1770
box -8 -3 16 105
use FILL  FILL_2917
timestamp 1745462530
transform 1 0 1128 0 1 1770
box -8 -3 16 105
use FILL  FILL_2918
timestamp 1745462530
transform 1 0 1096 0 1 1770
box -8 -3 16 105
use FILL  FILL_2919
timestamp 1745462530
transform 1 0 1088 0 1 1770
box -8 -3 16 105
use FILL  FILL_2920
timestamp 1745462530
transform 1 0 1056 0 1 1770
box -8 -3 16 105
use FILL  FILL_2921
timestamp 1745462530
transform 1 0 1048 0 1 1770
box -8 -3 16 105
use FILL  FILL_2922
timestamp 1745462530
transform 1 0 1008 0 1 1770
box -8 -3 16 105
use FILL  FILL_2923
timestamp 1745462530
transform 1 0 1000 0 1 1770
box -8 -3 16 105
use FILL  FILL_2924
timestamp 1745462530
transform 1 0 992 0 1 1770
box -8 -3 16 105
use FILL  FILL_2925
timestamp 1745462530
transform 1 0 984 0 1 1770
box -8 -3 16 105
use FILL  FILL_2926
timestamp 1745462530
transform 1 0 952 0 1 1770
box -8 -3 16 105
use FILL  FILL_2927
timestamp 1745462530
transform 1 0 944 0 1 1770
box -8 -3 16 105
use FILL  FILL_2928
timestamp 1745462530
transform 1 0 904 0 1 1770
box -8 -3 16 105
use FILL  FILL_2929
timestamp 1745462530
transform 1 0 896 0 1 1770
box -8 -3 16 105
use FILL  FILL_2930
timestamp 1745462530
transform 1 0 888 0 1 1770
box -8 -3 16 105
use FILL  FILL_2931
timestamp 1745462530
transform 1 0 784 0 1 1770
box -8 -3 16 105
use FILL  FILL_2932
timestamp 1745462530
transform 1 0 760 0 1 1770
box -8 -3 16 105
use FILL  FILL_2933
timestamp 1745462530
transform 1 0 752 0 1 1770
box -8 -3 16 105
use FILL  FILL_2934
timestamp 1745462530
transform 1 0 744 0 1 1770
box -8 -3 16 105
use FILL  FILL_2935
timestamp 1745462530
transform 1 0 696 0 1 1770
box -8 -3 16 105
use FILL  FILL_2936
timestamp 1745462530
transform 1 0 688 0 1 1770
box -8 -3 16 105
use FILL  FILL_2937
timestamp 1745462530
transform 1 0 680 0 1 1770
box -8 -3 16 105
use FILL  FILL_2938
timestamp 1745462530
transform 1 0 656 0 1 1770
box -8 -3 16 105
use FILL  FILL_2939
timestamp 1745462530
transform 1 0 648 0 1 1770
box -8 -3 16 105
use FILL  FILL_2940
timestamp 1745462530
transform 1 0 640 0 1 1770
box -8 -3 16 105
use FILL  FILL_2941
timestamp 1745462530
transform 1 0 592 0 1 1770
box -8 -3 16 105
use FILL  FILL_2942
timestamp 1745462530
transform 1 0 584 0 1 1770
box -8 -3 16 105
use FILL  FILL_2943
timestamp 1745462530
transform 1 0 576 0 1 1770
box -8 -3 16 105
use FILL  FILL_2944
timestamp 1745462530
transform 1 0 568 0 1 1770
box -8 -3 16 105
use FILL  FILL_2945
timestamp 1745462530
transform 1 0 464 0 1 1770
box -8 -3 16 105
use FILL  FILL_2946
timestamp 1745462530
transform 1 0 456 0 1 1770
box -8 -3 16 105
use FILL  FILL_2947
timestamp 1745462530
transform 1 0 448 0 1 1770
box -8 -3 16 105
use FILL  FILL_2948
timestamp 1745462530
transform 1 0 400 0 1 1770
box -8 -3 16 105
use FILL  FILL_2949
timestamp 1745462530
transform 1 0 392 0 1 1770
box -8 -3 16 105
use FILL  FILL_2950
timestamp 1745462530
transform 1 0 368 0 1 1770
box -8 -3 16 105
use FILL  FILL_2951
timestamp 1745462530
transform 1 0 320 0 1 1770
box -8 -3 16 105
use FILL  FILL_2952
timestamp 1745462530
transform 1 0 312 0 1 1770
box -8 -3 16 105
use FILL  FILL_2953
timestamp 1745462530
transform 1 0 304 0 1 1770
box -8 -3 16 105
use FILL  FILL_2954
timestamp 1745462530
transform 1 0 256 0 1 1770
box -8 -3 16 105
use FILL  FILL_2955
timestamp 1745462530
transform 1 0 248 0 1 1770
box -8 -3 16 105
use FILL  FILL_2956
timestamp 1745462530
transform 1 0 240 0 1 1770
box -8 -3 16 105
use FILL  FILL_2957
timestamp 1745462530
transform 1 0 216 0 1 1770
box -8 -3 16 105
use FILL  FILL_2958
timestamp 1745462530
transform 1 0 208 0 1 1770
box -8 -3 16 105
use FILL  FILL_2959
timestamp 1745462530
transform 1 0 160 0 1 1770
box -8 -3 16 105
use FILL  FILL_2960
timestamp 1745462530
transform 1 0 152 0 1 1770
box -8 -3 16 105
use FILL  FILL_2961
timestamp 1745462530
transform 1 0 144 0 1 1770
box -8 -3 16 105
use FILL  FILL_2962
timestamp 1745462530
transform 1 0 136 0 1 1770
box -8 -3 16 105
use FILL  FILL_2963
timestamp 1745462530
transform 1 0 128 0 1 1770
box -8 -3 16 105
use FILL  FILL_2964
timestamp 1745462530
transform 1 0 120 0 1 1770
box -8 -3 16 105
use FILL  FILL_2965
timestamp 1745462530
transform 1 0 112 0 1 1770
box -8 -3 16 105
use FILL  FILL_2966
timestamp 1745462530
transform 1 0 104 0 1 1770
box -8 -3 16 105
use FILL  FILL_2967
timestamp 1745462530
transform 1 0 96 0 1 1770
box -8 -3 16 105
use FILL  FILL_2968
timestamp 1745462530
transform 1 0 88 0 1 1770
box -8 -3 16 105
use FILL  FILL_2969
timestamp 1745462530
transform 1 0 80 0 1 1770
box -8 -3 16 105
use FILL  FILL_2970
timestamp 1745462530
transform 1 0 72 0 1 1770
box -8 -3 16 105
use FILL  FILL_2971
timestamp 1745462530
transform 1 0 4272 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2972
timestamp 1745462530
transform 1 0 4264 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2973
timestamp 1745462530
transform 1 0 4088 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2974
timestamp 1745462530
transform 1 0 4040 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2975
timestamp 1745462530
transform 1 0 4032 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2976
timestamp 1745462530
transform 1 0 3928 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2977
timestamp 1745462530
transform 1 0 3904 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2978
timestamp 1745462530
transform 1 0 3856 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2979
timestamp 1745462530
transform 1 0 3832 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2980
timestamp 1745462530
transform 1 0 3760 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2981
timestamp 1745462530
transform 1 0 3752 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2982
timestamp 1745462530
transform 1 0 3744 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2983
timestamp 1745462530
transform 1 0 3696 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2984
timestamp 1745462530
transform 1 0 3688 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2985
timestamp 1745462530
transform 1 0 3584 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2986
timestamp 1745462530
transform 1 0 3544 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2987
timestamp 1745462530
transform 1 0 3536 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2988
timestamp 1745462530
transform 1 0 3488 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2989
timestamp 1745462530
transform 1 0 3480 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2990
timestamp 1745462530
transform 1 0 3472 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2991
timestamp 1745462530
transform 1 0 3440 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2992
timestamp 1745462530
transform 1 0 3400 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2993
timestamp 1745462530
transform 1 0 3392 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2994
timestamp 1745462530
transform 1 0 3384 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2995
timestamp 1745462530
transform 1 0 3376 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2996
timestamp 1745462530
transform 1 0 3328 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2997
timestamp 1745462530
transform 1 0 3320 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2998
timestamp 1745462530
transform 1 0 3312 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2999
timestamp 1745462530
transform 1 0 3264 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3000
timestamp 1745462530
transform 1 0 3240 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3001
timestamp 1745462530
transform 1 0 3232 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3002
timestamp 1745462530
transform 1 0 3184 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3003
timestamp 1745462530
transform 1 0 3176 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3004
timestamp 1745462530
transform 1 0 3168 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3005
timestamp 1745462530
transform 1 0 3120 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3006
timestamp 1745462530
transform 1 0 3112 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3007
timestamp 1745462530
transform 1 0 3104 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3008
timestamp 1745462530
transform 1 0 3064 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3009
timestamp 1745462530
transform 1 0 3032 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3010
timestamp 1745462530
transform 1 0 3024 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3011
timestamp 1745462530
transform 1 0 3016 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3012
timestamp 1745462530
transform 1 0 2968 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3013
timestamp 1745462530
transform 1 0 2960 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3014
timestamp 1745462530
transform 1 0 2952 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3015
timestamp 1745462530
transform 1 0 2904 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3016
timestamp 1745462530
transform 1 0 2896 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3017
timestamp 1745462530
transform 1 0 2888 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3018
timestamp 1745462530
transform 1 0 2840 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3019
timestamp 1745462530
transform 1 0 2832 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3020
timestamp 1745462530
transform 1 0 2808 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3021
timestamp 1745462530
transform 1 0 2800 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3022
timestamp 1745462530
transform 1 0 2752 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3023
timestamp 1745462530
transform 1 0 2744 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3024
timestamp 1745462530
transform 1 0 2688 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3025
timestamp 1745462530
transform 1 0 2648 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3026
timestamp 1745462530
transform 1 0 2640 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3027
timestamp 1745462530
transform 1 0 2632 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3028
timestamp 1745462530
transform 1 0 2592 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3029
timestamp 1745462530
transform 1 0 2584 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3030
timestamp 1745462530
transform 1 0 2552 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3031
timestamp 1745462530
transform 1 0 2520 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3032
timestamp 1745462530
transform 1 0 2512 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3033
timestamp 1745462530
transform 1 0 2472 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3034
timestamp 1745462530
transform 1 0 2464 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3035
timestamp 1745462530
transform 1 0 2456 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3036
timestamp 1745462530
transform 1 0 2416 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3037
timestamp 1745462530
transform 1 0 2384 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3038
timestamp 1745462530
transform 1 0 2376 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3039
timestamp 1745462530
transform 1 0 2336 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3040
timestamp 1745462530
transform 1 0 2328 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3041
timestamp 1745462530
transform 1 0 2320 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3042
timestamp 1745462530
transform 1 0 2280 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3043
timestamp 1745462530
transform 1 0 2248 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3044
timestamp 1745462530
transform 1 0 2240 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3045
timestamp 1745462530
transform 1 0 2184 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3046
timestamp 1745462530
transform 1 0 2104 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3047
timestamp 1745462530
transform 1 0 2096 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3048
timestamp 1745462530
transform 1 0 2088 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3049
timestamp 1745462530
transform 1 0 2040 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3050
timestamp 1745462530
transform 1 0 2032 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3051
timestamp 1745462530
transform 1 0 1976 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3052
timestamp 1745462530
transform 1 0 1944 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3053
timestamp 1745462530
transform 1 0 1936 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3054
timestamp 1745462530
transform 1 0 1928 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3055
timestamp 1745462530
transform 1 0 1888 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3056
timestamp 1745462530
transform 1 0 1880 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3057
timestamp 1745462530
transform 1 0 1824 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3058
timestamp 1745462530
transform 1 0 1816 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3059
timestamp 1745462530
transform 1 0 1808 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3060
timestamp 1745462530
transform 1 0 1776 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3061
timestamp 1745462530
transform 1 0 1744 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3062
timestamp 1745462530
transform 1 0 1736 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3063
timestamp 1745462530
transform 1 0 1728 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3064
timestamp 1745462530
transform 1 0 1672 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3065
timestamp 1745462530
transform 1 0 1640 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3066
timestamp 1745462530
transform 1 0 1608 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3067
timestamp 1745462530
transform 1 0 1600 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3068
timestamp 1745462530
transform 1 0 1568 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3069
timestamp 1745462530
transform 1 0 1560 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3070
timestamp 1745462530
transform 1 0 1552 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3071
timestamp 1745462530
transform 1 0 1544 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3072
timestamp 1745462530
transform 1 0 1504 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3073
timestamp 1745462530
transform 1 0 1496 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3074
timestamp 1745462530
transform 1 0 1488 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3075
timestamp 1745462530
transform 1 0 1480 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3076
timestamp 1745462530
transform 1 0 1432 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3077
timestamp 1745462530
transform 1 0 1424 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3078
timestamp 1745462530
transform 1 0 1320 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3079
timestamp 1745462530
transform 1 0 1288 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3080
timestamp 1745462530
transform 1 0 1280 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3081
timestamp 1745462530
transform 1 0 1272 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3082
timestamp 1745462530
transform 1 0 1232 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3083
timestamp 1745462530
transform 1 0 1224 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3084
timestamp 1745462530
transform 1 0 1216 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3085
timestamp 1745462530
transform 1 0 1208 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3086
timestamp 1745462530
transform 1 0 1160 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3087
timestamp 1745462530
transform 1 0 1152 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3088
timestamp 1745462530
transform 1 0 1144 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3089
timestamp 1745462530
transform 1 0 1136 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3090
timestamp 1745462530
transform 1 0 1128 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3091
timestamp 1745462530
transform 1 0 1080 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3092
timestamp 1745462530
transform 1 0 1072 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3093
timestamp 1745462530
transform 1 0 1064 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3094
timestamp 1745462530
transform 1 0 1032 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3095
timestamp 1745462530
transform 1 0 1024 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3096
timestamp 1745462530
transform 1 0 1016 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3097
timestamp 1745462530
transform 1 0 976 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3098
timestamp 1745462530
transform 1 0 968 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3099
timestamp 1745462530
transform 1 0 960 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3100
timestamp 1745462530
transform 1 0 928 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3101
timestamp 1745462530
transform 1 0 920 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3102
timestamp 1745462530
transform 1 0 912 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3103
timestamp 1745462530
transform 1 0 904 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3104
timestamp 1745462530
transform 1 0 864 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3105
timestamp 1745462530
transform 1 0 856 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3106
timestamp 1745462530
transform 1 0 848 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3107
timestamp 1745462530
transform 1 0 744 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3108
timestamp 1745462530
transform 1 0 736 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3109
timestamp 1745462530
transform 1 0 712 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3110
timestamp 1745462530
transform 1 0 704 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3111
timestamp 1745462530
transform 1 0 696 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3112
timestamp 1745462530
transform 1 0 688 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3113
timestamp 1745462530
transform 1 0 640 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3114
timestamp 1745462530
transform 1 0 632 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3115
timestamp 1745462530
transform 1 0 624 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3116
timestamp 1745462530
transform 1 0 616 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3117
timestamp 1745462530
transform 1 0 608 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3118
timestamp 1745462530
transform 1 0 568 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3119
timestamp 1745462530
transform 1 0 560 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3120
timestamp 1745462530
transform 1 0 552 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3121
timestamp 1745462530
transform 1 0 544 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3122
timestamp 1745462530
transform 1 0 496 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3123
timestamp 1745462530
transform 1 0 488 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3124
timestamp 1745462530
transform 1 0 480 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3125
timestamp 1745462530
transform 1 0 472 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3126
timestamp 1745462530
transform 1 0 408 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3127
timestamp 1745462530
transform 1 0 400 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3128
timestamp 1745462530
transform 1 0 392 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3129
timestamp 1745462530
transform 1 0 288 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3130
timestamp 1745462530
transform 1 0 280 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3131
timestamp 1745462530
transform 1 0 256 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3132
timestamp 1745462530
transform 1 0 248 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3133
timestamp 1745462530
transform 1 0 240 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3134
timestamp 1745462530
transform 1 0 192 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3135
timestamp 1745462530
transform 1 0 184 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3136
timestamp 1745462530
transform 1 0 176 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3137
timestamp 1745462530
transform 1 0 72 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3138
timestamp 1745462530
transform 1 0 4368 0 1 1570
box -8 -3 16 105
use FILL  FILL_3139
timestamp 1745462530
transform 1 0 4344 0 1 1570
box -8 -3 16 105
use FILL  FILL_3140
timestamp 1745462530
transform 1 0 4296 0 1 1570
box -8 -3 16 105
use FILL  FILL_3141
timestamp 1745462530
transform 1 0 4192 0 1 1570
box -8 -3 16 105
use FILL  FILL_3142
timestamp 1745462530
transform 1 0 4144 0 1 1570
box -8 -3 16 105
use FILL  FILL_3143
timestamp 1745462530
transform 1 0 4120 0 1 1570
box -8 -3 16 105
use FILL  FILL_3144
timestamp 1745462530
transform 1 0 4072 0 1 1570
box -8 -3 16 105
use FILL  FILL_3145
timestamp 1745462530
transform 1 0 3968 0 1 1570
box -8 -3 16 105
use FILL  FILL_3146
timestamp 1745462530
transform 1 0 3960 0 1 1570
box -8 -3 16 105
use FILL  FILL_3147
timestamp 1745462530
transform 1 0 3856 0 1 1570
box -8 -3 16 105
use FILL  FILL_3148
timestamp 1745462530
transform 1 0 3792 0 1 1570
box -8 -3 16 105
use FILL  FILL_3149
timestamp 1745462530
transform 1 0 3784 0 1 1570
box -8 -3 16 105
use FILL  FILL_3150
timestamp 1745462530
transform 1 0 3744 0 1 1570
box -8 -3 16 105
use FILL  FILL_3151
timestamp 1745462530
transform 1 0 3696 0 1 1570
box -8 -3 16 105
use FILL  FILL_3152
timestamp 1745462530
transform 1 0 3688 0 1 1570
box -8 -3 16 105
use FILL  FILL_3153
timestamp 1745462530
transform 1 0 3680 0 1 1570
box -8 -3 16 105
use FILL  FILL_3154
timestamp 1745462530
transform 1 0 3632 0 1 1570
box -8 -3 16 105
use FILL  FILL_3155
timestamp 1745462530
transform 1 0 3608 0 1 1570
box -8 -3 16 105
use FILL  FILL_3156
timestamp 1745462530
transform 1 0 3600 0 1 1570
box -8 -3 16 105
use FILL  FILL_3157
timestamp 1745462530
transform 1 0 3552 0 1 1570
box -8 -3 16 105
use FILL  FILL_3158
timestamp 1745462530
transform 1 0 3544 0 1 1570
box -8 -3 16 105
use FILL  FILL_3159
timestamp 1745462530
transform 1 0 3536 0 1 1570
box -8 -3 16 105
use FILL  FILL_3160
timestamp 1745462530
transform 1 0 3432 0 1 1570
box -8 -3 16 105
use FILL  FILL_3161
timestamp 1745462530
transform 1 0 3424 0 1 1570
box -8 -3 16 105
use FILL  FILL_3162
timestamp 1745462530
transform 1 0 3400 0 1 1570
box -8 -3 16 105
use FILL  FILL_3163
timestamp 1745462530
transform 1 0 3392 0 1 1570
box -8 -3 16 105
use FILL  FILL_3164
timestamp 1745462530
transform 1 0 3360 0 1 1570
box -8 -3 16 105
use FILL  FILL_3165
timestamp 1745462530
transform 1 0 3352 0 1 1570
box -8 -3 16 105
use FILL  FILL_3166
timestamp 1745462530
transform 1 0 3344 0 1 1570
box -8 -3 16 105
use FILL  FILL_3167
timestamp 1745462530
transform 1 0 3240 0 1 1570
box -8 -3 16 105
use FILL  FILL_3168
timestamp 1745462530
transform 1 0 3232 0 1 1570
box -8 -3 16 105
use FILL  FILL_3169
timestamp 1745462530
transform 1 0 3184 0 1 1570
box -8 -3 16 105
use FILL  FILL_3170
timestamp 1745462530
transform 1 0 3176 0 1 1570
box -8 -3 16 105
use FILL  FILL_3171
timestamp 1745462530
transform 1 0 3168 0 1 1570
box -8 -3 16 105
use FILL  FILL_3172
timestamp 1745462530
transform 1 0 3160 0 1 1570
box -8 -3 16 105
use FILL  FILL_3173
timestamp 1745462530
transform 1 0 3152 0 1 1570
box -8 -3 16 105
use FILL  FILL_3174
timestamp 1745462530
transform 1 0 3104 0 1 1570
box -8 -3 16 105
use FILL  FILL_3175
timestamp 1745462530
transform 1 0 3096 0 1 1570
box -8 -3 16 105
use FILL  FILL_3176
timestamp 1745462530
transform 1 0 3088 0 1 1570
box -8 -3 16 105
use FILL  FILL_3177
timestamp 1745462530
transform 1 0 3048 0 1 1570
box -8 -3 16 105
use FILL  FILL_3178
timestamp 1745462530
transform 1 0 3040 0 1 1570
box -8 -3 16 105
use FILL  FILL_3179
timestamp 1745462530
transform 1 0 3032 0 1 1570
box -8 -3 16 105
use FILL  FILL_3180
timestamp 1745462530
transform 1 0 2992 0 1 1570
box -8 -3 16 105
use FILL  FILL_3181
timestamp 1745462530
transform 1 0 2984 0 1 1570
box -8 -3 16 105
use FILL  FILL_3182
timestamp 1745462530
transform 1 0 2952 0 1 1570
box -8 -3 16 105
use FILL  FILL_3183
timestamp 1745462530
transform 1 0 2944 0 1 1570
box -8 -3 16 105
use FILL  FILL_3184
timestamp 1745462530
transform 1 0 2936 0 1 1570
box -8 -3 16 105
use FILL  FILL_3185
timestamp 1745462530
transform 1 0 2928 0 1 1570
box -8 -3 16 105
use FILL  FILL_3186
timestamp 1745462530
transform 1 0 2888 0 1 1570
box -8 -3 16 105
use FILL  FILL_3187
timestamp 1745462530
transform 1 0 2880 0 1 1570
box -8 -3 16 105
use FILL  FILL_3188
timestamp 1745462530
transform 1 0 2872 0 1 1570
box -8 -3 16 105
use FILL  FILL_3189
timestamp 1745462530
transform 1 0 2768 0 1 1570
box -8 -3 16 105
use FILL  FILL_3190
timestamp 1745462530
transform 1 0 2760 0 1 1570
box -8 -3 16 105
use FILL  FILL_3191
timestamp 1745462530
transform 1 0 2752 0 1 1570
box -8 -3 16 105
use FILL  FILL_3192
timestamp 1745462530
transform 1 0 2696 0 1 1570
box -8 -3 16 105
use FILL  FILL_3193
timestamp 1745462530
transform 1 0 2688 0 1 1570
box -8 -3 16 105
use FILL  FILL_3194
timestamp 1745462530
transform 1 0 2680 0 1 1570
box -8 -3 16 105
use FILL  FILL_3195
timestamp 1745462530
transform 1 0 2672 0 1 1570
box -8 -3 16 105
use FILL  FILL_3196
timestamp 1745462530
transform 1 0 2640 0 1 1570
box -8 -3 16 105
use FILL  FILL_3197
timestamp 1745462530
transform 1 0 2632 0 1 1570
box -8 -3 16 105
use FILL  FILL_3198
timestamp 1745462530
transform 1 0 2624 0 1 1570
box -8 -3 16 105
use FILL  FILL_3199
timestamp 1745462530
transform 1 0 2592 0 1 1570
box -8 -3 16 105
use FILL  FILL_3200
timestamp 1745462530
transform 1 0 2560 0 1 1570
box -8 -3 16 105
use FILL  FILL_3201
timestamp 1745462530
transform 1 0 2552 0 1 1570
box -8 -3 16 105
use FILL  FILL_3202
timestamp 1745462530
transform 1 0 2544 0 1 1570
box -8 -3 16 105
use FILL  FILL_3203
timestamp 1745462530
transform 1 0 2536 0 1 1570
box -8 -3 16 105
use FILL  FILL_3204
timestamp 1745462530
transform 1 0 2528 0 1 1570
box -8 -3 16 105
use FILL  FILL_3205
timestamp 1745462530
transform 1 0 2488 0 1 1570
box -8 -3 16 105
use FILL  FILL_3206
timestamp 1745462530
transform 1 0 2480 0 1 1570
box -8 -3 16 105
use FILL  FILL_3207
timestamp 1745462530
transform 1 0 2472 0 1 1570
box -8 -3 16 105
use FILL  FILL_3208
timestamp 1745462530
transform 1 0 2464 0 1 1570
box -8 -3 16 105
use FILL  FILL_3209
timestamp 1745462530
transform 1 0 2456 0 1 1570
box -8 -3 16 105
use FILL  FILL_3210
timestamp 1745462530
transform 1 0 2416 0 1 1570
box -8 -3 16 105
use FILL  FILL_3211
timestamp 1745462530
transform 1 0 2408 0 1 1570
box -8 -3 16 105
use FILL  FILL_3212
timestamp 1745462530
transform 1 0 2400 0 1 1570
box -8 -3 16 105
use FILL  FILL_3213
timestamp 1745462530
transform 1 0 2392 0 1 1570
box -8 -3 16 105
use FILL  FILL_3214
timestamp 1745462530
transform 1 0 2352 0 1 1570
box -8 -3 16 105
use FILL  FILL_3215
timestamp 1745462530
transform 1 0 2344 0 1 1570
box -8 -3 16 105
use FILL  FILL_3216
timestamp 1745462530
transform 1 0 2336 0 1 1570
box -8 -3 16 105
use FILL  FILL_3217
timestamp 1745462530
transform 1 0 2304 0 1 1570
box -8 -3 16 105
use FILL  FILL_3218
timestamp 1745462530
transform 1 0 2296 0 1 1570
box -8 -3 16 105
use FILL  FILL_3219
timestamp 1745462530
transform 1 0 2288 0 1 1570
box -8 -3 16 105
use FILL  FILL_3220
timestamp 1745462530
transform 1 0 2248 0 1 1570
box -8 -3 16 105
use FILL  FILL_3221
timestamp 1745462530
transform 1 0 2240 0 1 1570
box -8 -3 16 105
use FILL  FILL_3222
timestamp 1745462530
transform 1 0 2232 0 1 1570
box -8 -3 16 105
use FILL  FILL_3223
timestamp 1745462530
transform 1 0 2224 0 1 1570
box -8 -3 16 105
use FILL  FILL_3224
timestamp 1745462530
transform 1 0 2168 0 1 1570
box -8 -3 16 105
use FILL  FILL_3225
timestamp 1745462530
transform 1 0 2160 0 1 1570
box -8 -3 16 105
use FILL  FILL_3226
timestamp 1745462530
transform 1 0 2152 0 1 1570
box -8 -3 16 105
use FILL  FILL_3227
timestamp 1745462530
transform 1 0 2096 0 1 1570
box -8 -3 16 105
use FILL  FILL_3228
timestamp 1745462530
transform 1 0 2088 0 1 1570
box -8 -3 16 105
use FILL  FILL_3229
timestamp 1745462530
transform 1 0 2080 0 1 1570
box -8 -3 16 105
use FILL  FILL_3230
timestamp 1745462530
transform 1 0 2024 0 1 1570
box -8 -3 16 105
use FILL  FILL_3231
timestamp 1745462530
transform 1 0 2016 0 1 1570
box -8 -3 16 105
use FILL  FILL_3232
timestamp 1745462530
transform 1 0 2008 0 1 1570
box -8 -3 16 105
use FILL  FILL_3233
timestamp 1745462530
transform 1 0 1952 0 1 1570
box -8 -3 16 105
use FILL  FILL_3234
timestamp 1745462530
transform 1 0 1944 0 1 1570
box -8 -3 16 105
use FILL  FILL_3235
timestamp 1745462530
transform 1 0 1936 0 1 1570
box -8 -3 16 105
use FILL  FILL_3236
timestamp 1745462530
transform 1 0 1928 0 1 1570
box -8 -3 16 105
use FILL  FILL_3237
timestamp 1745462530
transform 1 0 1880 0 1 1570
box -8 -3 16 105
use FILL  FILL_3238
timestamp 1745462530
transform 1 0 1872 0 1 1570
box -8 -3 16 105
use FILL  FILL_3239
timestamp 1745462530
transform 1 0 1864 0 1 1570
box -8 -3 16 105
use FILL  FILL_3240
timestamp 1745462530
transform 1 0 1832 0 1 1570
box -8 -3 16 105
use FILL  FILL_3241
timestamp 1745462530
transform 1 0 1824 0 1 1570
box -8 -3 16 105
use FILL  FILL_3242
timestamp 1745462530
transform 1 0 1776 0 1 1570
box -8 -3 16 105
use FILL  FILL_3243
timestamp 1745462530
transform 1 0 1768 0 1 1570
box -8 -3 16 105
use FILL  FILL_3244
timestamp 1745462530
transform 1 0 1760 0 1 1570
box -8 -3 16 105
use FILL  FILL_3245
timestamp 1745462530
transform 1 0 1752 0 1 1570
box -8 -3 16 105
use FILL  FILL_3246
timestamp 1745462530
transform 1 0 1744 0 1 1570
box -8 -3 16 105
use FILL  FILL_3247
timestamp 1745462530
transform 1 0 1704 0 1 1570
box -8 -3 16 105
use FILL  FILL_3248
timestamp 1745462530
transform 1 0 1696 0 1 1570
box -8 -3 16 105
use FILL  FILL_3249
timestamp 1745462530
transform 1 0 1688 0 1 1570
box -8 -3 16 105
use FILL  FILL_3250
timestamp 1745462530
transform 1 0 1680 0 1 1570
box -8 -3 16 105
use FILL  FILL_3251
timestamp 1745462530
transform 1 0 1648 0 1 1570
box -8 -3 16 105
use FILL  FILL_3252
timestamp 1745462530
transform 1 0 1616 0 1 1570
box -8 -3 16 105
use FILL  FILL_3253
timestamp 1745462530
transform 1 0 1608 0 1 1570
box -8 -3 16 105
use FILL  FILL_3254
timestamp 1745462530
transform 1 0 1600 0 1 1570
box -8 -3 16 105
use FILL  FILL_3255
timestamp 1745462530
transform 1 0 1592 0 1 1570
box -8 -3 16 105
use FILL  FILL_3256
timestamp 1745462530
transform 1 0 1544 0 1 1570
box -8 -3 16 105
use FILL  FILL_3257
timestamp 1745462530
transform 1 0 1536 0 1 1570
box -8 -3 16 105
use FILL  FILL_3258
timestamp 1745462530
transform 1 0 1528 0 1 1570
box -8 -3 16 105
use FILL  FILL_3259
timestamp 1745462530
transform 1 0 1520 0 1 1570
box -8 -3 16 105
use FILL  FILL_3260
timestamp 1745462530
transform 1 0 1480 0 1 1570
box -8 -3 16 105
use FILL  FILL_3261
timestamp 1745462530
transform 1 0 1472 0 1 1570
box -8 -3 16 105
use FILL  FILL_3262
timestamp 1745462530
transform 1 0 1464 0 1 1570
box -8 -3 16 105
use FILL  FILL_3263
timestamp 1745462530
transform 1 0 1432 0 1 1570
box -8 -3 16 105
use FILL  FILL_3264
timestamp 1745462530
transform 1 0 1424 0 1 1570
box -8 -3 16 105
use FILL  FILL_3265
timestamp 1745462530
transform 1 0 1392 0 1 1570
box -8 -3 16 105
use FILL  FILL_3266
timestamp 1745462530
transform 1 0 1384 0 1 1570
box -8 -3 16 105
use FILL  FILL_3267
timestamp 1745462530
transform 1 0 1376 0 1 1570
box -8 -3 16 105
use FILL  FILL_3268
timestamp 1745462530
transform 1 0 1368 0 1 1570
box -8 -3 16 105
use FILL  FILL_3269
timestamp 1745462530
transform 1 0 1328 0 1 1570
box -8 -3 16 105
use FILL  FILL_3270
timestamp 1745462530
transform 1 0 1320 0 1 1570
box -8 -3 16 105
use FILL  FILL_3271
timestamp 1745462530
transform 1 0 1312 0 1 1570
box -8 -3 16 105
use FILL  FILL_3272
timestamp 1745462530
transform 1 0 1280 0 1 1570
box -8 -3 16 105
use FILL  FILL_3273
timestamp 1745462530
transform 1 0 1248 0 1 1570
box -8 -3 16 105
use FILL  FILL_3274
timestamp 1745462530
transform 1 0 1240 0 1 1570
box -8 -3 16 105
use FILL  FILL_3275
timestamp 1745462530
transform 1 0 1208 0 1 1570
box -8 -3 16 105
use FILL  FILL_3276
timestamp 1745462530
transform 1 0 1200 0 1 1570
box -8 -3 16 105
use FILL  FILL_3277
timestamp 1745462530
transform 1 0 1192 0 1 1570
box -8 -3 16 105
use FILL  FILL_3278
timestamp 1745462530
transform 1 0 1184 0 1 1570
box -8 -3 16 105
use FILL  FILL_3279
timestamp 1745462530
transform 1 0 1136 0 1 1570
box -8 -3 16 105
use FILL  FILL_3280
timestamp 1745462530
transform 1 0 1128 0 1 1570
box -8 -3 16 105
use FILL  FILL_3281
timestamp 1745462530
transform 1 0 1096 0 1 1570
box -8 -3 16 105
use FILL  FILL_3282
timestamp 1745462530
transform 1 0 1088 0 1 1570
box -8 -3 16 105
use FILL  FILL_3283
timestamp 1745462530
transform 1 0 1080 0 1 1570
box -8 -3 16 105
use FILL  FILL_3284
timestamp 1745462530
transform 1 0 1032 0 1 1570
box -8 -3 16 105
use FILL  FILL_3285
timestamp 1745462530
transform 1 0 1024 0 1 1570
box -8 -3 16 105
use FILL  FILL_3286
timestamp 1745462530
transform 1 0 1016 0 1 1570
box -8 -3 16 105
use FILL  FILL_3287
timestamp 1745462530
transform 1 0 1008 0 1 1570
box -8 -3 16 105
use FILL  FILL_3288
timestamp 1745462530
transform 1 0 1000 0 1 1570
box -8 -3 16 105
use FILL  FILL_3289
timestamp 1745462530
transform 1 0 968 0 1 1570
box -8 -3 16 105
use FILL  FILL_3290
timestamp 1745462530
transform 1 0 960 0 1 1570
box -8 -3 16 105
use FILL  FILL_3291
timestamp 1745462530
transform 1 0 952 0 1 1570
box -8 -3 16 105
use FILL  FILL_3292
timestamp 1745462530
transform 1 0 944 0 1 1570
box -8 -3 16 105
use FILL  FILL_3293
timestamp 1745462530
transform 1 0 904 0 1 1570
box -8 -3 16 105
use FILL  FILL_3294
timestamp 1745462530
transform 1 0 896 0 1 1570
box -8 -3 16 105
use FILL  FILL_3295
timestamp 1745462530
transform 1 0 888 0 1 1570
box -8 -3 16 105
use FILL  FILL_3296
timestamp 1745462530
transform 1 0 880 0 1 1570
box -8 -3 16 105
use FILL  FILL_3297
timestamp 1745462530
transform 1 0 776 0 1 1570
box -8 -3 16 105
use FILL  FILL_3298
timestamp 1745462530
transform 1 0 768 0 1 1570
box -8 -3 16 105
use FILL  FILL_3299
timestamp 1745462530
transform 1 0 760 0 1 1570
box -8 -3 16 105
use FILL  FILL_3300
timestamp 1745462530
transform 1 0 736 0 1 1570
box -8 -3 16 105
use FILL  FILL_3301
timestamp 1745462530
transform 1 0 728 0 1 1570
box -8 -3 16 105
use FILL  FILL_3302
timestamp 1745462530
transform 1 0 720 0 1 1570
box -8 -3 16 105
use FILL  FILL_3303
timestamp 1745462530
transform 1 0 712 0 1 1570
box -8 -3 16 105
use FILL  FILL_3304
timestamp 1745462530
transform 1 0 664 0 1 1570
box -8 -3 16 105
use FILL  FILL_3305
timestamp 1745462530
transform 1 0 656 0 1 1570
box -8 -3 16 105
use FILL  FILL_3306
timestamp 1745462530
transform 1 0 648 0 1 1570
box -8 -3 16 105
use FILL  FILL_3307
timestamp 1745462530
transform 1 0 624 0 1 1570
box -8 -3 16 105
use FILL  FILL_3308
timestamp 1745462530
transform 1 0 616 0 1 1570
box -8 -3 16 105
use FILL  FILL_3309
timestamp 1745462530
transform 1 0 608 0 1 1570
box -8 -3 16 105
use FILL  FILL_3310
timestamp 1745462530
transform 1 0 600 0 1 1570
box -8 -3 16 105
use FILL  FILL_3311
timestamp 1745462530
transform 1 0 552 0 1 1570
box -8 -3 16 105
use FILL  FILL_3312
timestamp 1745462530
transform 1 0 544 0 1 1570
box -8 -3 16 105
use FILL  FILL_3313
timestamp 1745462530
transform 1 0 536 0 1 1570
box -8 -3 16 105
use FILL  FILL_3314
timestamp 1745462530
transform 1 0 528 0 1 1570
box -8 -3 16 105
use FILL  FILL_3315
timestamp 1745462530
transform 1 0 520 0 1 1570
box -8 -3 16 105
use FILL  FILL_3316
timestamp 1745462530
transform 1 0 416 0 1 1570
box -8 -3 16 105
use FILL  FILL_3317
timestamp 1745462530
transform 1 0 408 0 1 1570
box -8 -3 16 105
use FILL  FILL_3318
timestamp 1745462530
transform 1 0 384 0 1 1570
box -8 -3 16 105
use FILL  FILL_3319
timestamp 1745462530
transform 1 0 376 0 1 1570
box -8 -3 16 105
use FILL  FILL_3320
timestamp 1745462530
transform 1 0 328 0 1 1570
box -8 -3 16 105
use FILL  FILL_3321
timestamp 1745462530
transform 1 0 320 0 1 1570
box -8 -3 16 105
use FILL  FILL_3322
timestamp 1745462530
transform 1 0 296 0 1 1570
box -8 -3 16 105
use FILL  FILL_3323
timestamp 1745462530
transform 1 0 288 0 1 1570
box -8 -3 16 105
use FILL  FILL_3324
timestamp 1745462530
transform 1 0 184 0 1 1570
box -8 -3 16 105
use FILL  FILL_3325
timestamp 1745462530
transform 1 0 176 0 1 1570
box -8 -3 16 105
use FILL  FILL_3326
timestamp 1745462530
transform 1 0 168 0 1 1570
box -8 -3 16 105
use FILL  FILL_3327
timestamp 1745462530
transform 1 0 160 0 1 1570
box -8 -3 16 105
use FILL  FILL_3328
timestamp 1745462530
transform 1 0 152 0 1 1570
box -8 -3 16 105
use FILL  FILL_3329
timestamp 1745462530
transform 1 0 144 0 1 1570
box -8 -3 16 105
use FILL  FILL_3330
timestamp 1745462530
transform 1 0 136 0 1 1570
box -8 -3 16 105
use FILL  FILL_3331
timestamp 1745462530
transform 1 0 128 0 1 1570
box -8 -3 16 105
use FILL  FILL_3332
timestamp 1745462530
transform 1 0 120 0 1 1570
box -8 -3 16 105
use FILL  FILL_3333
timestamp 1745462530
transform 1 0 112 0 1 1570
box -8 -3 16 105
use FILL  FILL_3334
timestamp 1745462530
transform 1 0 104 0 1 1570
box -8 -3 16 105
use FILL  FILL_3335
timestamp 1745462530
transform 1 0 96 0 1 1570
box -8 -3 16 105
use FILL  FILL_3336
timestamp 1745462530
transform 1 0 88 0 1 1570
box -8 -3 16 105
use FILL  FILL_3337
timestamp 1745462530
transform 1 0 80 0 1 1570
box -8 -3 16 105
use FILL  FILL_3338
timestamp 1745462530
transform 1 0 72 0 1 1570
box -8 -3 16 105
use FILL  FILL_3339
timestamp 1745462530
transform 1 0 4256 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3340
timestamp 1745462530
transform 1 0 4248 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3341
timestamp 1745462530
transform 1 0 4200 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3342
timestamp 1745462530
transform 1 0 4096 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3343
timestamp 1745462530
transform 1 0 4048 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3344
timestamp 1745462530
transform 1 0 4024 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3345
timestamp 1745462530
transform 1 0 4016 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3346
timestamp 1745462530
transform 1 0 3968 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3347
timestamp 1745462530
transform 1 0 3960 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3348
timestamp 1745462530
transform 1 0 3952 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3349
timestamp 1745462530
transform 1 0 3912 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3350
timestamp 1745462530
transform 1 0 3904 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3351
timestamp 1745462530
transform 1 0 3856 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3352
timestamp 1745462530
transform 1 0 3848 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3353
timestamp 1745462530
transform 1 0 3840 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3354
timestamp 1745462530
transform 1 0 3808 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3355
timestamp 1745462530
transform 1 0 3800 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3356
timestamp 1745462530
transform 1 0 3760 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3357
timestamp 1745462530
transform 1 0 3752 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3358
timestamp 1745462530
transform 1 0 3744 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3359
timestamp 1745462530
transform 1 0 3736 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3360
timestamp 1745462530
transform 1 0 3680 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3361
timestamp 1745462530
transform 1 0 3672 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3362
timestamp 1745462530
transform 1 0 3664 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3363
timestamp 1745462530
transform 1 0 3656 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3364
timestamp 1745462530
transform 1 0 3608 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3365
timestamp 1745462530
transform 1 0 3600 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3366
timestamp 1745462530
transform 1 0 3592 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3367
timestamp 1745462530
transform 1 0 3584 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3368
timestamp 1745462530
transform 1 0 3576 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3369
timestamp 1745462530
transform 1 0 3568 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3370
timestamp 1745462530
transform 1 0 3536 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3371
timestamp 1745462530
transform 1 0 3528 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3372
timestamp 1745462530
transform 1 0 3520 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3373
timestamp 1745462530
transform 1 0 3512 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3374
timestamp 1745462530
transform 1 0 3504 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3375
timestamp 1745462530
transform 1 0 3456 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3376
timestamp 1745462530
transform 1 0 3448 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3377
timestamp 1745462530
transform 1 0 3440 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3378
timestamp 1745462530
transform 1 0 3432 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3379
timestamp 1745462530
transform 1 0 3424 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3380
timestamp 1745462530
transform 1 0 3376 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3381
timestamp 1745462530
transform 1 0 3368 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3382
timestamp 1745462530
transform 1 0 3360 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3383
timestamp 1745462530
transform 1 0 3352 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3384
timestamp 1745462530
transform 1 0 3344 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3385
timestamp 1745462530
transform 1 0 3296 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3386
timestamp 1745462530
transform 1 0 3288 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3387
timestamp 1745462530
transform 1 0 3280 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3388
timestamp 1745462530
transform 1 0 3272 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3389
timestamp 1745462530
transform 1 0 3264 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3390
timestamp 1745462530
transform 1 0 3224 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3391
timestamp 1745462530
transform 1 0 3216 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3392
timestamp 1745462530
transform 1 0 3208 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3393
timestamp 1745462530
transform 1 0 3200 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3394
timestamp 1745462530
transform 1 0 3192 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3395
timestamp 1745462530
transform 1 0 3152 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3396
timestamp 1745462530
transform 1 0 3144 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3397
timestamp 1745462530
transform 1 0 3136 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3398
timestamp 1745462530
transform 1 0 3128 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3399
timestamp 1745462530
transform 1 0 3120 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3400
timestamp 1745462530
transform 1 0 3072 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3401
timestamp 1745462530
transform 1 0 3064 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3402
timestamp 1745462530
transform 1 0 3056 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3403
timestamp 1745462530
transform 1 0 3048 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3404
timestamp 1745462530
transform 1 0 3040 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3405
timestamp 1745462530
transform 1 0 2992 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3406
timestamp 1745462530
transform 1 0 2984 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3407
timestamp 1745462530
transform 1 0 2976 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3408
timestamp 1745462530
transform 1 0 2968 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3409
timestamp 1745462530
transform 1 0 2936 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3410
timestamp 1745462530
transform 1 0 2928 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3411
timestamp 1745462530
transform 1 0 2920 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3412
timestamp 1745462530
transform 1 0 2912 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3413
timestamp 1745462530
transform 1 0 2856 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3414
timestamp 1745462530
transform 1 0 2848 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3415
timestamp 1745462530
transform 1 0 2840 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3416
timestamp 1745462530
transform 1 0 2832 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3417
timestamp 1745462530
transform 1 0 2784 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3418
timestamp 1745462530
transform 1 0 2776 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3419
timestamp 1745462530
transform 1 0 2768 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3420
timestamp 1745462530
transform 1 0 2760 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3421
timestamp 1745462530
transform 1 0 2656 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3422
timestamp 1745462530
transform 1 0 2648 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3423
timestamp 1745462530
transform 1 0 2640 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3424
timestamp 1745462530
transform 1 0 2608 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3425
timestamp 1745462530
transform 1 0 2576 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3426
timestamp 1745462530
transform 1 0 2544 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3427
timestamp 1745462530
transform 1 0 2536 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3428
timestamp 1745462530
transform 1 0 2504 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3429
timestamp 1745462530
transform 1 0 2496 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3430
timestamp 1745462530
transform 1 0 2488 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3431
timestamp 1745462530
transform 1 0 2480 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3432
timestamp 1745462530
transform 1 0 2440 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3433
timestamp 1745462530
transform 1 0 2432 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3434
timestamp 1745462530
transform 1 0 2424 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3435
timestamp 1745462530
transform 1 0 2320 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3436
timestamp 1745462530
transform 1 0 2312 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3437
timestamp 1745462530
transform 1 0 2304 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3438
timestamp 1745462530
transform 1 0 2256 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3439
timestamp 1745462530
transform 1 0 2248 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3440
timestamp 1745462530
transform 1 0 2240 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3441
timestamp 1745462530
transform 1 0 2232 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3442
timestamp 1745462530
transform 1 0 2176 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3443
timestamp 1745462530
transform 1 0 2168 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3444
timestamp 1745462530
transform 1 0 2112 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3445
timestamp 1745462530
transform 1 0 2104 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3446
timestamp 1745462530
transform 1 0 2000 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3447
timestamp 1745462530
transform 1 0 1992 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3448
timestamp 1745462530
transform 1 0 1936 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3449
timestamp 1745462530
transform 1 0 1928 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3450
timestamp 1745462530
transform 1 0 1920 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3451
timestamp 1745462530
transform 1 0 1880 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3452
timestamp 1745462530
transform 1 0 1872 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3453
timestamp 1745462530
transform 1 0 1864 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3454
timestamp 1745462530
transform 1 0 1832 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3455
timestamp 1745462530
transform 1 0 1824 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3456
timestamp 1745462530
transform 1 0 1816 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3457
timestamp 1745462530
transform 1 0 1784 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3458
timestamp 1745462530
transform 1 0 1752 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3459
timestamp 1745462530
transform 1 0 1744 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3460
timestamp 1745462530
transform 1 0 1712 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3461
timestamp 1745462530
transform 1 0 1704 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3462
timestamp 1745462530
transform 1 0 1696 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3463
timestamp 1745462530
transform 1 0 1664 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3464
timestamp 1745462530
transform 1 0 1560 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3465
timestamp 1745462530
transform 1 0 1552 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3466
timestamp 1745462530
transform 1 0 1544 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3467
timestamp 1745462530
transform 1 0 1536 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3468
timestamp 1745462530
transform 1 0 1496 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3469
timestamp 1745462530
transform 1 0 1488 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3470
timestamp 1745462530
transform 1 0 1480 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3471
timestamp 1745462530
transform 1 0 1472 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3472
timestamp 1745462530
transform 1 0 1440 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3473
timestamp 1745462530
transform 1 0 1432 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3474
timestamp 1745462530
transform 1 0 1424 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3475
timestamp 1745462530
transform 1 0 1416 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3476
timestamp 1745462530
transform 1 0 1368 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3477
timestamp 1745462530
transform 1 0 1360 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3478
timestamp 1745462530
transform 1 0 1352 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3479
timestamp 1745462530
transform 1 0 1296 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3480
timestamp 1745462530
transform 1 0 1264 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3481
timestamp 1745462530
transform 1 0 1256 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3482
timestamp 1745462530
transform 1 0 1248 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3483
timestamp 1745462530
transform 1 0 1208 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3484
timestamp 1745462530
transform 1 0 1200 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3485
timestamp 1745462530
transform 1 0 1192 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3486
timestamp 1745462530
transform 1 0 1184 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3487
timestamp 1745462530
transform 1 0 1176 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3488
timestamp 1745462530
transform 1 0 1144 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3489
timestamp 1745462530
transform 1 0 1136 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3490
timestamp 1745462530
transform 1 0 1128 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3491
timestamp 1745462530
transform 1 0 1096 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3492
timestamp 1745462530
transform 1 0 1088 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3493
timestamp 1745462530
transform 1 0 1080 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3494
timestamp 1745462530
transform 1 0 1040 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3495
timestamp 1745462530
transform 1 0 1032 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3496
timestamp 1745462530
transform 1 0 1024 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3497
timestamp 1745462530
transform 1 0 992 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3498
timestamp 1745462530
transform 1 0 984 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3499
timestamp 1745462530
transform 1 0 976 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3500
timestamp 1745462530
transform 1 0 936 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3501
timestamp 1745462530
transform 1 0 928 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3502
timestamp 1745462530
transform 1 0 896 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3503
timestamp 1745462530
transform 1 0 888 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3504
timestamp 1745462530
transform 1 0 784 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3505
timestamp 1745462530
transform 1 0 776 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3506
timestamp 1745462530
transform 1 0 752 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3507
timestamp 1745462530
transform 1 0 648 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3508
timestamp 1745462530
transform 1 0 640 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3509
timestamp 1745462530
transform 1 0 632 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3510
timestamp 1745462530
transform 1 0 528 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3511
timestamp 1745462530
transform 1 0 520 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3512
timestamp 1745462530
transform 1 0 512 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3513
timestamp 1745462530
transform 1 0 464 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3514
timestamp 1745462530
transform 1 0 456 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3515
timestamp 1745462530
transform 1 0 448 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3516
timestamp 1745462530
transform 1 0 400 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3517
timestamp 1745462530
transform 1 0 392 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3518
timestamp 1745462530
transform 1 0 384 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3519
timestamp 1745462530
transform 1 0 336 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3520
timestamp 1745462530
transform 1 0 328 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3521
timestamp 1745462530
transform 1 0 320 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3522
timestamp 1745462530
transform 1 0 272 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3523
timestamp 1745462530
transform 1 0 264 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3524
timestamp 1745462530
transform 1 0 256 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3525
timestamp 1745462530
transform 1 0 248 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3526
timestamp 1745462530
transform 1 0 200 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3527
timestamp 1745462530
transform 1 0 176 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3528
timestamp 1745462530
transform 1 0 72 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3529
timestamp 1745462530
transform 1 0 4368 0 1 1370
box -8 -3 16 105
use FILL  FILL_3530
timestamp 1745462530
transform 1 0 4264 0 1 1370
box -8 -3 16 105
use FILL  FILL_3531
timestamp 1745462530
transform 1 0 4240 0 1 1370
box -8 -3 16 105
use FILL  FILL_3532
timestamp 1745462530
transform 1 0 4192 0 1 1370
box -8 -3 16 105
use FILL  FILL_3533
timestamp 1745462530
transform 1 0 4184 0 1 1370
box -8 -3 16 105
use FILL  FILL_3534
timestamp 1745462530
transform 1 0 4176 0 1 1370
box -8 -3 16 105
use FILL  FILL_3535
timestamp 1745462530
transform 1 0 4128 0 1 1370
box -8 -3 16 105
use FILL  FILL_3536
timestamp 1745462530
transform 1 0 4120 0 1 1370
box -8 -3 16 105
use FILL  FILL_3537
timestamp 1745462530
transform 1 0 4112 0 1 1370
box -8 -3 16 105
use FILL  FILL_3538
timestamp 1745462530
transform 1 0 4064 0 1 1370
box -8 -3 16 105
use FILL  FILL_3539
timestamp 1745462530
transform 1 0 4040 0 1 1370
box -8 -3 16 105
use FILL  FILL_3540
timestamp 1745462530
transform 1 0 4032 0 1 1370
box -8 -3 16 105
use FILL  FILL_3541
timestamp 1745462530
transform 1 0 3928 0 1 1370
box -8 -3 16 105
use FILL  FILL_3542
timestamp 1745462530
transform 1 0 3920 0 1 1370
box -8 -3 16 105
use FILL  FILL_3543
timestamp 1745462530
transform 1 0 3912 0 1 1370
box -8 -3 16 105
use FILL  FILL_3544
timestamp 1745462530
transform 1 0 3864 0 1 1370
box -8 -3 16 105
use FILL  FILL_3545
timestamp 1745462530
transform 1 0 3856 0 1 1370
box -8 -3 16 105
use FILL  FILL_3546
timestamp 1745462530
transform 1 0 3832 0 1 1370
box -8 -3 16 105
use FILL  FILL_3547
timestamp 1745462530
transform 1 0 3784 0 1 1370
box -8 -3 16 105
use FILL  FILL_3548
timestamp 1745462530
transform 1 0 3776 0 1 1370
box -8 -3 16 105
use FILL  FILL_3549
timestamp 1745462530
transform 1 0 3728 0 1 1370
box -8 -3 16 105
use FILL  FILL_3550
timestamp 1745462530
transform 1 0 3720 0 1 1370
box -8 -3 16 105
use FILL  FILL_3551
timestamp 1745462530
transform 1 0 3712 0 1 1370
box -8 -3 16 105
use FILL  FILL_3552
timestamp 1745462530
transform 1 0 3704 0 1 1370
box -8 -3 16 105
use FILL  FILL_3553
timestamp 1745462530
transform 1 0 3656 0 1 1370
box -8 -3 16 105
use FILL  FILL_3554
timestamp 1745462530
transform 1 0 3648 0 1 1370
box -8 -3 16 105
use FILL  FILL_3555
timestamp 1745462530
transform 1 0 3624 0 1 1370
box -8 -3 16 105
use FILL  FILL_3556
timestamp 1745462530
transform 1 0 3616 0 1 1370
box -8 -3 16 105
use FILL  FILL_3557
timestamp 1745462530
transform 1 0 3608 0 1 1370
box -8 -3 16 105
use FILL  FILL_3558
timestamp 1745462530
transform 1 0 3560 0 1 1370
box -8 -3 16 105
use FILL  FILL_3559
timestamp 1745462530
transform 1 0 3552 0 1 1370
box -8 -3 16 105
use FILL  FILL_3560
timestamp 1745462530
transform 1 0 3544 0 1 1370
box -8 -3 16 105
use FILL  FILL_3561
timestamp 1745462530
transform 1 0 3536 0 1 1370
box -8 -3 16 105
use FILL  FILL_3562
timestamp 1745462530
transform 1 0 3488 0 1 1370
box -8 -3 16 105
use FILL  FILL_3563
timestamp 1745462530
transform 1 0 3480 0 1 1370
box -8 -3 16 105
use FILL  FILL_3564
timestamp 1745462530
transform 1 0 3456 0 1 1370
box -8 -3 16 105
use FILL  FILL_3565
timestamp 1745462530
transform 1 0 3448 0 1 1370
box -8 -3 16 105
use FILL  FILL_3566
timestamp 1745462530
transform 1 0 3440 0 1 1370
box -8 -3 16 105
use FILL  FILL_3567
timestamp 1745462530
transform 1 0 3392 0 1 1370
box -8 -3 16 105
use FILL  FILL_3568
timestamp 1745462530
transform 1 0 3384 0 1 1370
box -8 -3 16 105
use FILL  FILL_3569
timestamp 1745462530
transform 1 0 3376 0 1 1370
box -8 -3 16 105
use FILL  FILL_3570
timestamp 1745462530
transform 1 0 3368 0 1 1370
box -8 -3 16 105
use FILL  FILL_3571
timestamp 1745462530
transform 1 0 3336 0 1 1370
box -8 -3 16 105
use FILL  FILL_3572
timestamp 1745462530
transform 1 0 3328 0 1 1370
box -8 -3 16 105
use FILL  FILL_3573
timestamp 1745462530
transform 1 0 3296 0 1 1370
box -8 -3 16 105
use FILL  FILL_3574
timestamp 1745462530
transform 1 0 3288 0 1 1370
box -8 -3 16 105
use FILL  FILL_3575
timestamp 1745462530
transform 1 0 3280 0 1 1370
box -8 -3 16 105
use FILL  FILL_3576
timestamp 1745462530
transform 1 0 3248 0 1 1370
box -8 -3 16 105
use FILL  FILL_3577
timestamp 1745462530
transform 1 0 3240 0 1 1370
box -8 -3 16 105
use FILL  FILL_3578
timestamp 1745462530
transform 1 0 3232 0 1 1370
box -8 -3 16 105
use FILL  FILL_3579
timestamp 1745462530
transform 1 0 3184 0 1 1370
box -8 -3 16 105
use FILL  FILL_3580
timestamp 1745462530
transform 1 0 3176 0 1 1370
box -8 -3 16 105
use FILL  FILL_3581
timestamp 1745462530
transform 1 0 3168 0 1 1370
box -8 -3 16 105
use FILL  FILL_3582
timestamp 1745462530
transform 1 0 3160 0 1 1370
box -8 -3 16 105
use FILL  FILL_3583
timestamp 1745462530
transform 1 0 3128 0 1 1370
box -8 -3 16 105
use FILL  FILL_3584
timestamp 1745462530
transform 1 0 3096 0 1 1370
box -8 -3 16 105
use FILL  FILL_3585
timestamp 1745462530
transform 1 0 3088 0 1 1370
box -8 -3 16 105
use FILL  FILL_3586
timestamp 1745462530
transform 1 0 3080 0 1 1370
box -8 -3 16 105
use FILL  FILL_3587
timestamp 1745462530
transform 1 0 3072 0 1 1370
box -8 -3 16 105
use FILL  FILL_3588
timestamp 1745462530
transform 1 0 3024 0 1 1370
box -8 -3 16 105
use FILL  FILL_3589
timestamp 1745462530
transform 1 0 3016 0 1 1370
box -8 -3 16 105
use FILL  FILL_3590
timestamp 1745462530
transform 1 0 3008 0 1 1370
box -8 -3 16 105
use FILL  FILL_3591
timestamp 1745462530
transform 1 0 2904 0 1 1370
box -8 -3 16 105
use FILL  FILL_3592
timestamp 1745462530
transform 1 0 2880 0 1 1370
box -8 -3 16 105
use FILL  FILL_3593
timestamp 1745462530
transform 1 0 2872 0 1 1370
box -8 -3 16 105
use FILL  FILL_3594
timestamp 1745462530
transform 1 0 2824 0 1 1370
box -8 -3 16 105
use FILL  FILL_3595
timestamp 1745462530
transform 1 0 2816 0 1 1370
box -8 -3 16 105
use FILL  FILL_3596
timestamp 1745462530
transform 1 0 2808 0 1 1370
box -8 -3 16 105
use FILL  FILL_3597
timestamp 1745462530
transform 1 0 2800 0 1 1370
box -8 -3 16 105
use FILL  FILL_3598
timestamp 1745462530
transform 1 0 2768 0 1 1370
box -8 -3 16 105
use FILL  FILL_3599
timestamp 1745462530
transform 1 0 2760 0 1 1370
box -8 -3 16 105
use FILL  FILL_3600
timestamp 1745462530
transform 1 0 2720 0 1 1370
box -8 -3 16 105
use FILL  FILL_3601
timestamp 1745462530
transform 1 0 2712 0 1 1370
box -8 -3 16 105
use FILL  FILL_3602
timestamp 1745462530
transform 1 0 2704 0 1 1370
box -8 -3 16 105
use FILL  FILL_3603
timestamp 1745462530
transform 1 0 2680 0 1 1370
box -8 -3 16 105
use FILL  FILL_3604
timestamp 1745462530
transform 1 0 2672 0 1 1370
box -8 -3 16 105
use FILL  FILL_3605
timestamp 1745462530
transform 1 0 2664 0 1 1370
box -8 -3 16 105
use FILL  FILL_3606
timestamp 1745462530
transform 1 0 2616 0 1 1370
box -8 -3 16 105
use FILL  FILL_3607
timestamp 1745462530
transform 1 0 2608 0 1 1370
box -8 -3 16 105
use FILL  FILL_3608
timestamp 1745462530
transform 1 0 2600 0 1 1370
box -8 -3 16 105
use FILL  FILL_3609
timestamp 1745462530
transform 1 0 2544 0 1 1370
box -8 -3 16 105
use FILL  FILL_3610
timestamp 1745462530
transform 1 0 2536 0 1 1370
box -8 -3 16 105
use FILL  FILL_3611
timestamp 1745462530
transform 1 0 2528 0 1 1370
box -8 -3 16 105
use FILL  FILL_3612
timestamp 1745462530
transform 1 0 2480 0 1 1370
box -8 -3 16 105
use FILL  FILL_3613
timestamp 1745462530
transform 1 0 2472 0 1 1370
box -8 -3 16 105
use FILL  FILL_3614
timestamp 1745462530
transform 1 0 2464 0 1 1370
box -8 -3 16 105
use FILL  FILL_3615
timestamp 1745462530
transform 1 0 2440 0 1 1370
box -8 -3 16 105
use FILL  FILL_3616
timestamp 1745462530
transform 1 0 2432 0 1 1370
box -8 -3 16 105
use FILL  FILL_3617
timestamp 1745462530
transform 1 0 2424 0 1 1370
box -8 -3 16 105
use FILL  FILL_3618
timestamp 1745462530
transform 1 0 2376 0 1 1370
box -8 -3 16 105
use FILL  FILL_3619
timestamp 1745462530
transform 1 0 2368 0 1 1370
box -8 -3 16 105
use FILL  FILL_3620
timestamp 1745462530
transform 1 0 2360 0 1 1370
box -8 -3 16 105
use FILL  FILL_3621
timestamp 1745462530
transform 1 0 2352 0 1 1370
box -8 -3 16 105
use FILL  FILL_3622
timestamp 1745462530
transform 1 0 2312 0 1 1370
box -8 -3 16 105
use FILL  FILL_3623
timestamp 1745462530
transform 1 0 2304 0 1 1370
box -8 -3 16 105
use FILL  FILL_3624
timestamp 1745462530
transform 1 0 2296 0 1 1370
box -8 -3 16 105
use FILL  FILL_3625
timestamp 1745462530
transform 1 0 2288 0 1 1370
box -8 -3 16 105
use FILL  FILL_3626
timestamp 1745462530
transform 1 0 2256 0 1 1370
box -8 -3 16 105
use FILL  FILL_3627
timestamp 1745462530
transform 1 0 2248 0 1 1370
box -8 -3 16 105
use FILL  FILL_3628
timestamp 1745462530
transform 1 0 2240 0 1 1370
box -8 -3 16 105
use FILL  FILL_3629
timestamp 1745462530
transform 1 0 2208 0 1 1370
box -8 -3 16 105
use FILL  FILL_3630
timestamp 1745462530
transform 1 0 2200 0 1 1370
box -8 -3 16 105
use FILL  FILL_3631
timestamp 1745462530
transform 1 0 2168 0 1 1370
box -8 -3 16 105
use FILL  FILL_3632
timestamp 1745462530
transform 1 0 2160 0 1 1370
box -8 -3 16 105
use FILL  FILL_3633
timestamp 1745462530
transform 1 0 2128 0 1 1370
box -8 -3 16 105
use FILL  FILL_3634
timestamp 1745462530
transform 1 0 2120 0 1 1370
box -8 -3 16 105
use FILL  FILL_3635
timestamp 1745462530
transform 1 0 2088 0 1 1370
box -8 -3 16 105
use FILL  FILL_3636
timestamp 1745462530
transform 1 0 2080 0 1 1370
box -8 -3 16 105
use FILL  FILL_3637
timestamp 1745462530
transform 1 0 2072 0 1 1370
box -8 -3 16 105
use FILL  FILL_3638
timestamp 1745462530
transform 1 0 2064 0 1 1370
box -8 -3 16 105
use FILL  FILL_3639
timestamp 1745462530
transform 1 0 2056 0 1 1370
box -8 -3 16 105
use FILL  FILL_3640
timestamp 1745462530
transform 1 0 2008 0 1 1370
box -8 -3 16 105
use FILL  FILL_3641
timestamp 1745462530
transform 1 0 2000 0 1 1370
box -8 -3 16 105
use FILL  FILL_3642
timestamp 1745462530
transform 1 0 1976 0 1 1370
box -8 -3 16 105
use FILL  FILL_3643
timestamp 1745462530
transform 1 0 1968 0 1 1370
box -8 -3 16 105
use FILL  FILL_3644
timestamp 1745462530
transform 1 0 1960 0 1 1370
box -8 -3 16 105
use FILL  FILL_3645
timestamp 1745462530
transform 1 0 1912 0 1 1370
box -8 -3 16 105
use FILL  FILL_3646
timestamp 1745462530
transform 1 0 1904 0 1 1370
box -8 -3 16 105
use FILL  FILL_3647
timestamp 1745462530
transform 1 0 1880 0 1 1370
box -8 -3 16 105
use FILL  FILL_3648
timestamp 1745462530
transform 1 0 1872 0 1 1370
box -8 -3 16 105
use FILL  FILL_3649
timestamp 1745462530
transform 1 0 1864 0 1 1370
box -8 -3 16 105
use FILL  FILL_3650
timestamp 1745462530
transform 1 0 1816 0 1 1370
box -8 -3 16 105
use FILL  FILL_3651
timestamp 1745462530
transform 1 0 1808 0 1 1370
box -8 -3 16 105
use FILL  FILL_3652
timestamp 1745462530
transform 1 0 1760 0 1 1370
box -8 -3 16 105
use FILL  FILL_3653
timestamp 1745462530
transform 1 0 1752 0 1 1370
box -8 -3 16 105
use FILL  FILL_3654
timestamp 1745462530
transform 1 0 1744 0 1 1370
box -8 -3 16 105
use FILL  FILL_3655
timestamp 1745462530
transform 1 0 1704 0 1 1370
box -8 -3 16 105
use FILL  FILL_3656
timestamp 1745462530
transform 1 0 1696 0 1 1370
box -8 -3 16 105
use FILL  FILL_3657
timestamp 1745462530
transform 1 0 1688 0 1 1370
box -8 -3 16 105
use FILL  FILL_3658
timestamp 1745462530
transform 1 0 1640 0 1 1370
box -8 -3 16 105
use FILL  FILL_3659
timestamp 1745462530
transform 1 0 1632 0 1 1370
box -8 -3 16 105
use FILL  FILL_3660
timestamp 1745462530
transform 1 0 1624 0 1 1370
box -8 -3 16 105
use FILL  FILL_3661
timestamp 1745462530
transform 1 0 1616 0 1 1370
box -8 -3 16 105
use FILL  FILL_3662
timestamp 1745462530
transform 1 0 1568 0 1 1370
box -8 -3 16 105
use FILL  FILL_3663
timestamp 1745462530
transform 1 0 1560 0 1 1370
box -8 -3 16 105
use FILL  FILL_3664
timestamp 1745462530
transform 1 0 1552 0 1 1370
box -8 -3 16 105
use FILL  FILL_3665
timestamp 1745462530
transform 1 0 1504 0 1 1370
box -8 -3 16 105
use FILL  FILL_3666
timestamp 1745462530
transform 1 0 1496 0 1 1370
box -8 -3 16 105
use FILL  FILL_3667
timestamp 1745462530
transform 1 0 1488 0 1 1370
box -8 -3 16 105
use FILL  FILL_3668
timestamp 1745462530
transform 1 0 1464 0 1 1370
box -8 -3 16 105
use FILL  FILL_3669
timestamp 1745462530
transform 1 0 1360 0 1 1370
box -8 -3 16 105
use FILL  FILL_3670
timestamp 1745462530
transform 1 0 1352 0 1 1370
box -8 -3 16 105
use FILL  FILL_3671
timestamp 1745462530
transform 1 0 1296 0 1 1370
box -8 -3 16 105
use FILL  FILL_3672
timestamp 1745462530
transform 1 0 1288 0 1 1370
box -8 -3 16 105
use FILL  FILL_3673
timestamp 1745462530
transform 1 0 1280 0 1 1370
box -8 -3 16 105
use FILL  FILL_3674
timestamp 1745462530
transform 1 0 1240 0 1 1370
box -8 -3 16 105
use FILL  FILL_3675
timestamp 1745462530
transform 1 0 1232 0 1 1370
box -8 -3 16 105
use FILL  FILL_3676
timestamp 1745462530
transform 1 0 1224 0 1 1370
box -8 -3 16 105
use FILL  FILL_3677
timestamp 1745462530
transform 1 0 1216 0 1 1370
box -8 -3 16 105
use FILL  FILL_3678
timestamp 1745462530
transform 1 0 1184 0 1 1370
box -8 -3 16 105
use FILL  FILL_3679
timestamp 1745462530
transform 1 0 1176 0 1 1370
box -8 -3 16 105
use FILL  FILL_3680
timestamp 1745462530
transform 1 0 1144 0 1 1370
box -8 -3 16 105
use FILL  FILL_3681
timestamp 1745462530
transform 1 0 1136 0 1 1370
box -8 -3 16 105
use FILL  FILL_3682
timestamp 1745462530
transform 1 0 1096 0 1 1370
box -8 -3 16 105
use FILL  FILL_3683
timestamp 1745462530
transform 1 0 1088 0 1 1370
box -8 -3 16 105
use FILL  FILL_3684
timestamp 1745462530
transform 1 0 1080 0 1 1370
box -8 -3 16 105
use FILL  FILL_3685
timestamp 1745462530
transform 1 0 1048 0 1 1370
box -8 -3 16 105
use FILL  FILL_3686
timestamp 1745462530
transform 1 0 1008 0 1 1370
box -8 -3 16 105
use FILL  FILL_3687
timestamp 1745462530
transform 1 0 1000 0 1 1370
box -8 -3 16 105
use FILL  FILL_3688
timestamp 1745462530
transform 1 0 992 0 1 1370
box -8 -3 16 105
use FILL  FILL_3689
timestamp 1745462530
transform 1 0 960 0 1 1370
box -8 -3 16 105
use FILL  FILL_3690
timestamp 1745462530
transform 1 0 952 0 1 1370
box -8 -3 16 105
use FILL  FILL_3691
timestamp 1745462530
transform 1 0 912 0 1 1370
box -8 -3 16 105
use FILL  FILL_3692
timestamp 1745462530
transform 1 0 888 0 1 1370
box -8 -3 16 105
use FILL  FILL_3693
timestamp 1745462530
transform 1 0 880 0 1 1370
box -8 -3 16 105
use FILL  FILL_3694
timestamp 1745462530
transform 1 0 872 0 1 1370
box -8 -3 16 105
use FILL  FILL_3695
timestamp 1745462530
transform 1 0 824 0 1 1370
box -8 -3 16 105
use FILL  FILL_3696
timestamp 1745462530
transform 1 0 816 0 1 1370
box -8 -3 16 105
use FILL  FILL_3697
timestamp 1745462530
transform 1 0 792 0 1 1370
box -8 -3 16 105
use FILL  FILL_3698
timestamp 1745462530
transform 1 0 744 0 1 1370
box -8 -3 16 105
use FILL  FILL_3699
timestamp 1745462530
transform 1 0 736 0 1 1370
box -8 -3 16 105
use FILL  FILL_3700
timestamp 1745462530
transform 1 0 728 0 1 1370
box -8 -3 16 105
use FILL  FILL_3701
timestamp 1745462530
transform 1 0 680 0 1 1370
box -8 -3 16 105
use FILL  FILL_3702
timestamp 1745462530
transform 1 0 672 0 1 1370
box -8 -3 16 105
use FILL  FILL_3703
timestamp 1745462530
transform 1 0 552 0 1 1370
box -8 -3 16 105
use FILL  FILL_3704
timestamp 1745462530
transform 1 0 544 0 1 1370
box -8 -3 16 105
use FILL  FILL_3705
timestamp 1745462530
transform 1 0 312 0 1 1370
box -8 -3 16 105
use FILL  FILL_3706
timestamp 1745462530
transform 1 0 192 0 1 1370
box -8 -3 16 105
use FILL  FILL_3707
timestamp 1745462530
transform 1 0 72 0 1 1370
box -8 -3 16 105
use FILL  FILL_3708
timestamp 1745462530
transform 1 0 4368 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3709
timestamp 1745462530
transform 1 0 4264 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3710
timestamp 1745462530
transform 1 0 4240 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3711
timestamp 1745462530
transform 1 0 4192 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3712
timestamp 1745462530
transform 1 0 4184 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3713
timestamp 1745462530
transform 1 0 4160 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3714
timestamp 1745462530
transform 1 0 4056 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3715
timestamp 1745462530
transform 1 0 4048 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3716
timestamp 1745462530
transform 1 0 4040 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3717
timestamp 1745462530
transform 1 0 4008 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3718
timestamp 1745462530
transform 1 0 4000 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3719
timestamp 1745462530
transform 1 0 3968 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3720
timestamp 1745462530
transform 1 0 3960 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3721
timestamp 1745462530
transform 1 0 3952 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3722
timestamp 1745462530
transform 1 0 3912 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3723
timestamp 1745462530
transform 1 0 3904 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3724
timestamp 1745462530
transform 1 0 3896 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3725
timestamp 1745462530
transform 1 0 3856 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3726
timestamp 1745462530
transform 1 0 3848 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3727
timestamp 1745462530
transform 1 0 3840 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3728
timestamp 1745462530
transform 1 0 3736 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3729
timestamp 1745462530
transform 1 0 3728 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3730
timestamp 1745462530
transform 1 0 3720 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3731
timestamp 1745462530
transform 1 0 3712 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3732
timestamp 1745462530
transform 1 0 3608 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3733
timestamp 1745462530
transform 1 0 3600 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3734
timestamp 1745462530
transform 1 0 3592 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3735
timestamp 1745462530
transform 1 0 3488 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3736
timestamp 1745462530
transform 1 0 3480 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3737
timestamp 1745462530
transform 1 0 3472 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3738
timestamp 1745462530
transform 1 0 3432 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3739
timestamp 1745462530
transform 1 0 3424 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3740
timestamp 1745462530
transform 1 0 3416 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3741
timestamp 1745462530
transform 1 0 3408 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3742
timestamp 1745462530
transform 1 0 3376 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3743
timestamp 1745462530
transform 1 0 3368 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3744
timestamp 1745462530
transform 1 0 3328 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3745
timestamp 1745462530
transform 1 0 3320 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3746
timestamp 1745462530
transform 1 0 3312 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3747
timestamp 1745462530
transform 1 0 3304 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3748
timestamp 1745462530
transform 1 0 3272 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3749
timestamp 1745462530
transform 1 0 3264 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3750
timestamp 1745462530
transform 1 0 3240 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3751
timestamp 1745462530
transform 1 0 3232 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3752
timestamp 1745462530
transform 1 0 3200 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3753
timestamp 1745462530
transform 1 0 3192 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3754
timestamp 1745462530
transform 1 0 3184 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3755
timestamp 1745462530
transform 1 0 3176 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3756
timestamp 1745462530
transform 1 0 3144 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3757
timestamp 1745462530
transform 1 0 3136 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3758
timestamp 1745462530
transform 1 0 3128 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3759
timestamp 1745462530
transform 1 0 3088 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3760
timestamp 1745462530
transform 1 0 3080 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3761
timestamp 1745462530
transform 1 0 3072 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3762
timestamp 1745462530
transform 1 0 3040 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3763
timestamp 1745462530
transform 1 0 3032 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3764
timestamp 1745462530
transform 1 0 2992 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3765
timestamp 1745462530
transform 1 0 2984 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3766
timestamp 1745462530
transform 1 0 2976 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3767
timestamp 1745462530
transform 1 0 2872 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3768
timestamp 1745462530
transform 1 0 2848 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3769
timestamp 1745462530
transform 1 0 2840 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3770
timestamp 1745462530
transform 1 0 2832 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3771
timestamp 1745462530
transform 1 0 2784 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3772
timestamp 1745462530
transform 1 0 2776 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3773
timestamp 1745462530
transform 1 0 2768 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3774
timestamp 1745462530
transform 1 0 2760 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3775
timestamp 1745462530
transform 1 0 2720 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3776
timestamp 1745462530
transform 1 0 2712 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3777
timestamp 1745462530
transform 1 0 2704 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3778
timestamp 1745462530
transform 1 0 2656 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3779
timestamp 1745462530
transform 1 0 2648 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3780
timestamp 1745462530
transform 1 0 2640 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3781
timestamp 1745462530
transform 1 0 2632 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3782
timestamp 1745462530
transform 1 0 2584 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3783
timestamp 1745462530
transform 1 0 2576 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3784
timestamp 1745462530
transform 1 0 2552 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3785
timestamp 1745462530
transform 1 0 2544 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3786
timestamp 1745462530
transform 1 0 2504 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3787
timestamp 1745462530
transform 1 0 2496 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3788
timestamp 1745462530
transform 1 0 2488 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3789
timestamp 1745462530
transform 1 0 2456 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3790
timestamp 1745462530
transform 1 0 2448 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3791
timestamp 1745462530
transform 1 0 2416 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3792
timestamp 1745462530
transform 1 0 2408 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3793
timestamp 1745462530
transform 1 0 2400 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3794
timestamp 1745462530
transform 1 0 2352 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3795
timestamp 1745462530
transform 1 0 2344 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3796
timestamp 1745462530
transform 1 0 2336 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3797
timestamp 1745462530
transform 1 0 2312 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3798
timestamp 1745462530
transform 1 0 2208 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3799
timestamp 1745462530
transform 1 0 2128 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3800
timestamp 1745462530
transform 1 0 2120 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3801
timestamp 1745462530
transform 1 0 2112 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3802
timestamp 1745462530
transform 1 0 2072 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3803
timestamp 1745462530
transform 1 0 2064 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3804
timestamp 1745462530
transform 1 0 2040 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3805
timestamp 1745462530
transform 1 0 2032 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3806
timestamp 1745462530
transform 1 0 2024 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3807
timestamp 1745462530
transform 1 0 1976 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3808
timestamp 1745462530
transform 1 0 1968 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3809
timestamp 1745462530
transform 1 0 1960 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3810
timestamp 1745462530
transform 1 0 1952 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3811
timestamp 1745462530
transform 1 0 1848 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3812
timestamp 1745462530
transform 1 0 1840 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3813
timestamp 1745462530
transform 1 0 1808 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3814
timestamp 1745462530
transform 1 0 1800 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3815
timestamp 1745462530
transform 1 0 1696 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3816
timestamp 1745462530
transform 1 0 1688 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3817
timestamp 1745462530
transform 1 0 1680 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3818
timestamp 1745462530
transform 1 0 1656 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3819
timestamp 1745462530
transform 1 0 1648 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3820
timestamp 1745462530
transform 1 0 1640 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3821
timestamp 1745462530
transform 1 0 1616 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3822
timestamp 1745462530
transform 1 0 1584 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3823
timestamp 1745462530
transform 1 0 1576 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3824
timestamp 1745462530
transform 1 0 1568 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3825
timestamp 1745462530
transform 1 0 1560 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3826
timestamp 1745462530
transform 1 0 1520 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3827
timestamp 1745462530
transform 1 0 1512 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3828
timestamp 1745462530
transform 1 0 1504 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3829
timestamp 1745462530
transform 1 0 1496 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3830
timestamp 1745462530
transform 1 0 1448 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3831
timestamp 1745462530
transform 1 0 1440 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3832
timestamp 1745462530
transform 1 0 1432 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3833
timestamp 1745462530
transform 1 0 1424 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3834
timestamp 1745462530
transform 1 0 1400 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3835
timestamp 1745462530
transform 1 0 1296 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3836
timestamp 1745462530
transform 1 0 1288 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3837
timestamp 1745462530
transform 1 0 1240 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3838
timestamp 1745462530
transform 1 0 1232 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3839
timestamp 1745462530
transform 1 0 1224 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3840
timestamp 1745462530
transform 1 0 1192 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3841
timestamp 1745462530
transform 1 0 1184 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3842
timestamp 1745462530
transform 1 0 1144 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3843
timestamp 1745462530
transform 1 0 1136 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3844
timestamp 1745462530
transform 1 0 1104 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3845
timestamp 1745462530
transform 1 0 1000 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3846
timestamp 1745462530
transform 1 0 976 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3847
timestamp 1745462530
transform 1 0 928 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3848
timestamp 1745462530
transform 1 0 920 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3849
timestamp 1745462530
transform 1 0 912 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3850
timestamp 1745462530
transform 1 0 888 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3851
timestamp 1745462530
transform 1 0 840 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3852
timestamp 1745462530
transform 1 0 832 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3853
timestamp 1745462530
transform 1 0 728 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3854
timestamp 1745462530
transform 1 0 720 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3855
timestamp 1745462530
transform 1 0 712 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3856
timestamp 1745462530
transform 1 0 664 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3857
timestamp 1745462530
transform 1 0 656 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3858
timestamp 1745462530
transform 1 0 632 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3859
timestamp 1745462530
transform 1 0 528 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3860
timestamp 1745462530
transform 1 0 464 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3861
timestamp 1745462530
transform 1 0 456 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3862
timestamp 1745462530
transform 1 0 352 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3863
timestamp 1745462530
transform 1 0 248 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3864
timestamp 1745462530
transform 1 0 240 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3865
timestamp 1745462530
transform 1 0 176 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3866
timestamp 1745462530
transform 1 0 72 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3867
timestamp 1745462530
transform 1 0 4272 0 1 1170
box -8 -3 16 105
use FILL  FILL_3868
timestamp 1745462530
transform 1 0 3976 0 1 1170
box -8 -3 16 105
use FILL  FILL_3869
timestamp 1745462530
transform 1 0 3952 0 1 1170
box -8 -3 16 105
use FILL  FILL_3870
timestamp 1745462530
transform 1 0 3904 0 1 1170
box -8 -3 16 105
use FILL  FILL_3871
timestamp 1745462530
transform 1 0 3856 0 1 1170
box -8 -3 16 105
use FILL  FILL_3872
timestamp 1745462530
transform 1 0 3832 0 1 1170
box -8 -3 16 105
use FILL  FILL_3873
timestamp 1745462530
transform 1 0 3808 0 1 1170
box -8 -3 16 105
use FILL  FILL_3874
timestamp 1745462530
transform 1 0 3760 0 1 1170
box -8 -3 16 105
use FILL  FILL_3875
timestamp 1745462530
transform 1 0 3752 0 1 1170
box -8 -3 16 105
use FILL  FILL_3876
timestamp 1745462530
transform 1 0 3704 0 1 1170
box -8 -3 16 105
use FILL  FILL_3877
timestamp 1745462530
transform 1 0 3696 0 1 1170
box -8 -3 16 105
use FILL  FILL_3878
timestamp 1745462530
transform 1 0 3656 0 1 1170
box -8 -3 16 105
use FILL  FILL_3879
timestamp 1745462530
transform 1 0 3648 0 1 1170
box -8 -3 16 105
use FILL  FILL_3880
timestamp 1745462530
transform 1 0 3640 0 1 1170
box -8 -3 16 105
use FILL  FILL_3881
timestamp 1745462530
transform 1 0 3576 0 1 1170
box -8 -3 16 105
use FILL  FILL_3882
timestamp 1745462530
transform 1 0 3568 0 1 1170
box -8 -3 16 105
use FILL  FILL_3883
timestamp 1745462530
transform 1 0 3528 0 1 1170
box -8 -3 16 105
use FILL  FILL_3884
timestamp 1745462530
transform 1 0 3496 0 1 1170
box -8 -3 16 105
use FILL  FILL_3885
timestamp 1745462530
transform 1 0 3488 0 1 1170
box -8 -3 16 105
use FILL  FILL_3886
timestamp 1745462530
transform 1 0 3480 0 1 1170
box -8 -3 16 105
use FILL  FILL_3887
timestamp 1745462530
transform 1 0 3432 0 1 1170
box -8 -3 16 105
use FILL  FILL_3888
timestamp 1745462530
transform 1 0 3408 0 1 1170
box -8 -3 16 105
use FILL  FILL_3889
timestamp 1745462530
transform 1 0 3400 0 1 1170
box -8 -3 16 105
use FILL  FILL_3890
timestamp 1745462530
transform 1 0 3352 0 1 1170
box -8 -3 16 105
use FILL  FILL_3891
timestamp 1745462530
transform 1 0 3344 0 1 1170
box -8 -3 16 105
use FILL  FILL_3892
timestamp 1745462530
transform 1 0 3320 0 1 1170
box -8 -3 16 105
use FILL  FILL_3893
timestamp 1745462530
transform 1 0 3216 0 1 1170
box -8 -3 16 105
use FILL  FILL_3894
timestamp 1745462530
transform 1 0 3208 0 1 1170
box -8 -3 16 105
use FILL  FILL_3895
timestamp 1745462530
transform 1 0 3176 0 1 1170
box -8 -3 16 105
use FILL  FILL_3896
timestamp 1745462530
transform 1 0 3168 0 1 1170
box -8 -3 16 105
use FILL  FILL_3897
timestamp 1745462530
transform 1 0 3136 0 1 1170
box -8 -3 16 105
use FILL  FILL_3898
timestamp 1745462530
transform 1 0 3128 0 1 1170
box -8 -3 16 105
use FILL  FILL_3899
timestamp 1745462530
transform 1 0 3088 0 1 1170
box -8 -3 16 105
use FILL  FILL_3900
timestamp 1745462530
transform 1 0 3080 0 1 1170
box -8 -3 16 105
use FILL  FILL_3901
timestamp 1745462530
transform 1 0 2976 0 1 1170
box -8 -3 16 105
use FILL  FILL_3902
timestamp 1745462530
transform 1 0 2968 0 1 1170
box -8 -3 16 105
use FILL  FILL_3903
timestamp 1745462530
transform 1 0 2960 0 1 1170
box -8 -3 16 105
use FILL  FILL_3904
timestamp 1745462530
transform 1 0 2912 0 1 1170
box -8 -3 16 105
use FILL  FILL_3905
timestamp 1745462530
transform 1 0 2904 0 1 1170
box -8 -3 16 105
use FILL  FILL_3906
timestamp 1745462530
transform 1 0 2880 0 1 1170
box -8 -3 16 105
use FILL  FILL_3907
timestamp 1745462530
transform 1 0 2832 0 1 1170
box -8 -3 16 105
use FILL  FILL_3908
timestamp 1745462530
transform 1 0 2824 0 1 1170
box -8 -3 16 105
use FILL  FILL_3909
timestamp 1745462530
transform 1 0 2816 0 1 1170
box -8 -3 16 105
use FILL  FILL_3910
timestamp 1745462530
transform 1 0 2768 0 1 1170
box -8 -3 16 105
use FILL  FILL_3911
timestamp 1745462530
transform 1 0 2760 0 1 1170
box -8 -3 16 105
use FILL  FILL_3912
timestamp 1745462530
transform 1 0 2752 0 1 1170
box -8 -3 16 105
use FILL  FILL_3913
timestamp 1745462530
transform 1 0 2648 0 1 1170
box -8 -3 16 105
use FILL  FILL_3914
timestamp 1745462530
transform 1 0 2544 0 1 1170
box -8 -3 16 105
use FILL  FILL_3915
timestamp 1745462530
transform 1 0 2536 0 1 1170
box -8 -3 16 105
use FILL  FILL_3916
timestamp 1745462530
transform 1 0 2488 0 1 1170
box -8 -3 16 105
use FILL  FILL_3917
timestamp 1745462530
transform 1 0 2480 0 1 1170
box -8 -3 16 105
use FILL  FILL_3918
timestamp 1745462530
transform 1 0 2472 0 1 1170
box -8 -3 16 105
use FILL  FILL_3919
timestamp 1745462530
transform 1 0 2424 0 1 1170
box -8 -3 16 105
use FILL  FILL_3920
timestamp 1745462530
transform 1 0 2416 0 1 1170
box -8 -3 16 105
use FILL  FILL_3921
timestamp 1745462530
transform 1 0 2312 0 1 1170
box -8 -3 16 105
use FILL  FILL_3922
timestamp 1745462530
transform 1 0 2304 0 1 1170
box -8 -3 16 105
use FILL  FILL_3923
timestamp 1745462530
transform 1 0 2272 0 1 1170
box -8 -3 16 105
use FILL  FILL_3924
timestamp 1745462530
transform 1 0 2168 0 1 1170
box -8 -3 16 105
use FILL  FILL_3925
timestamp 1745462530
transform 1 0 2160 0 1 1170
box -8 -3 16 105
use FILL  FILL_3926
timestamp 1745462530
transform 1 0 2056 0 1 1170
box -8 -3 16 105
use FILL  FILL_3927
timestamp 1745462530
transform 1 0 2032 0 1 1170
box -8 -3 16 105
use FILL  FILL_3928
timestamp 1745462530
transform 1 0 2024 0 1 1170
box -8 -3 16 105
use FILL  FILL_3929
timestamp 1745462530
transform 1 0 1976 0 1 1170
box -8 -3 16 105
use FILL  FILL_3930
timestamp 1745462530
transform 1 0 1968 0 1 1170
box -8 -3 16 105
use FILL  FILL_3931
timestamp 1745462530
transform 1 0 1960 0 1 1170
box -8 -3 16 105
use FILL  FILL_3932
timestamp 1745462530
transform 1 0 1936 0 1 1170
box -8 -3 16 105
use FILL  FILL_3933
timestamp 1745462530
transform 1 0 1928 0 1 1170
box -8 -3 16 105
use FILL  FILL_3934
timestamp 1745462530
transform 1 0 1880 0 1 1170
box -8 -3 16 105
use FILL  FILL_3935
timestamp 1745462530
transform 1 0 1872 0 1 1170
box -8 -3 16 105
use FILL  FILL_3936
timestamp 1745462530
transform 1 0 1864 0 1 1170
box -8 -3 16 105
use FILL  FILL_3937
timestamp 1745462530
transform 1 0 1816 0 1 1170
box -8 -3 16 105
use FILL  FILL_3938
timestamp 1745462530
transform 1 0 1808 0 1 1170
box -8 -3 16 105
use FILL  FILL_3939
timestamp 1745462530
transform 1 0 1688 0 1 1170
box -8 -3 16 105
use FILL  FILL_3940
timestamp 1745462530
transform 1 0 1680 0 1 1170
box -8 -3 16 105
use FILL  FILL_3941
timestamp 1745462530
transform 1 0 1632 0 1 1170
box -8 -3 16 105
use FILL  FILL_3942
timestamp 1745462530
transform 1 0 1624 0 1 1170
box -8 -3 16 105
use FILL  FILL_3943
timestamp 1745462530
transform 1 0 1616 0 1 1170
box -8 -3 16 105
use FILL  FILL_3944
timestamp 1745462530
transform 1 0 1568 0 1 1170
box -8 -3 16 105
use FILL  FILL_3945
timestamp 1745462530
transform 1 0 1560 0 1 1170
box -8 -3 16 105
use FILL  FILL_3946
timestamp 1745462530
transform 1 0 1552 0 1 1170
box -8 -3 16 105
use FILL  FILL_3947
timestamp 1745462530
transform 1 0 1528 0 1 1170
box -8 -3 16 105
use FILL  FILL_3948
timestamp 1745462530
transform 1 0 1520 0 1 1170
box -8 -3 16 105
use FILL  FILL_3949
timestamp 1745462530
transform 1 0 1472 0 1 1170
box -8 -3 16 105
use FILL  FILL_3950
timestamp 1745462530
transform 1 0 1464 0 1 1170
box -8 -3 16 105
use FILL  FILL_3951
timestamp 1745462530
transform 1 0 1456 0 1 1170
box -8 -3 16 105
use FILL  FILL_3952
timestamp 1745462530
transform 1 0 1448 0 1 1170
box -8 -3 16 105
use FILL  FILL_3953
timestamp 1745462530
transform 1 0 1440 0 1 1170
box -8 -3 16 105
use FILL  FILL_3954
timestamp 1745462530
transform 1 0 1392 0 1 1170
box -8 -3 16 105
use FILL  FILL_3955
timestamp 1745462530
transform 1 0 1384 0 1 1170
box -8 -3 16 105
use FILL  FILL_3956
timestamp 1745462530
transform 1 0 1376 0 1 1170
box -8 -3 16 105
use FILL  FILL_3957
timestamp 1745462530
transform 1 0 1368 0 1 1170
box -8 -3 16 105
use FILL  FILL_3958
timestamp 1745462530
transform 1 0 1360 0 1 1170
box -8 -3 16 105
use FILL  FILL_3959
timestamp 1745462530
transform 1 0 1336 0 1 1170
box -8 -3 16 105
use FILL  FILL_3960
timestamp 1745462530
transform 1 0 1328 0 1 1170
box -8 -3 16 105
use FILL  FILL_3961
timestamp 1745462530
transform 1 0 1320 0 1 1170
box -8 -3 16 105
use FILL  FILL_3962
timestamp 1745462530
transform 1 0 1272 0 1 1170
box -8 -3 16 105
use FILL  FILL_3963
timestamp 1745462530
transform 1 0 1264 0 1 1170
box -8 -3 16 105
use FILL  FILL_3964
timestamp 1745462530
transform 1 0 1256 0 1 1170
box -8 -3 16 105
use FILL  FILL_3965
timestamp 1745462530
transform 1 0 1248 0 1 1170
box -8 -3 16 105
use FILL  FILL_3966
timestamp 1745462530
transform 1 0 1240 0 1 1170
box -8 -3 16 105
use FILL  FILL_3967
timestamp 1745462530
transform 1 0 1208 0 1 1170
box -8 -3 16 105
use FILL  FILL_3968
timestamp 1745462530
transform 1 0 1200 0 1 1170
box -8 -3 16 105
use FILL  FILL_3969
timestamp 1745462530
transform 1 0 1192 0 1 1170
box -8 -3 16 105
use FILL  FILL_3970
timestamp 1745462530
transform 1 0 1184 0 1 1170
box -8 -3 16 105
use FILL  FILL_3971
timestamp 1745462530
transform 1 0 1152 0 1 1170
box -8 -3 16 105
use FILL  FILL_3972
timestamp 1745462530
transform 1 0 1144 0 1 1170
box -8 -3 16 105
use FILL  FILL_3973
timestamp 1745462530
transform 1 0 1136 0 1 1170
box -8 -3 16 105
use FILL  FILL_3974
timestamp 1745462530
transform 1 0 1104 0 1 1170
box -8 -3 16 105
use FILL  FILL_3975
timestamp 1745462530
transform 1 0 1096 0 1 1170
box -8 -3 16 105
use FILL  FILL_3976
timestamp 1745462530
transform 1 0 1088 0 1 1170
box -8 -3 16 105
use FILL  FILL_3977
timestamp 1745462530
transform 1 0 1080 0 1 1170
box -8 -3 16 105
use FILL  FILL_3978
timestamp 1745462530
transform 1 0 1040 0 1 1170
box -8 -3 16 105
use FILL  FILL_3979
timestamp 1745462530
transform 1 0 1032 0 1 1170
box -8 -3 16 105
use FILL  FILL_3980
timestamp 1745462530
transform 1 0 1024 0 1 1170
box -8 -3 16 105
use FILL  FILL_3981
timestamp 1745462530
transform 1 0 1016 0 1 1170
box -8 -3 16 105
use FILL  FILL_3982
timestamp 1745462530
transform 1 0 968 0 1 1170
box -8 -3 16 105
use FILL  FILL_3983
timestamp 1745462530
transform 1 0 960 0 1 1170
box -8 -3 16 105
use FILL  FILL_3984
timestamp 1745462530
transform 1 0 952 0 1 1170
box -8 -3 16 105
use FILL  FILL_3985
timestamp 1745462530
transform 1 0 920 0 1 1170
box -8 -3 16 105
use FILL  FILL_3986
timestamp 1745462530
transform 1 0 912 0 1 1170
box -8 -3 16 105
use FILL  FILL_3987
timestamp 1745462530
transform 1 0 864 0 1 1170
box -8 -3 16 105
use FILL  FILL_3988
timestamp 1745462530
transform 1 0 856 0 1 1170
box -8 -3 16 105
use FILL  FILL_3989
timestamp 1745462530
transform 1 0 848 0 1 1170
box -8 -3 16 105
use FILL  FILL_3990
timestamp 1745462530
transform 1 0 840 0 1 1170
box -8 -3 16 105
use FILL  FILL_3991
timestamp 1745462530
transform 1 0 792 0 1 1170
box -8 -3 16 105
use FILL  FILL_3992
timestamp 1745462530
transform 1 0 784 0 1 1170
box -8 -3 16 105
use FILL  FILL_3993
timestamp 1745462530
transform 1 0 776 0 1 1170
box -8 -3 16 105
use FILL  FILL_3994
timestamp 1745462530
transform 1 0 672 0 1 1170
box -8 -3 16 105
use FILL  FILL_3995
timestamp 1745462530
transform 1 0 664 0 1 1170
box -8 -3 16 105
use FILL  FILL_3996
timestamp 1745462530
transform 1 0 656 0 1 1170
box -8 -3 16 105
use FILL  FILL_3997
timestamp 1745462530
transform 1 0 608 0 1 1170
box -8 -3 16 105
use FILL  FILL_3998
timestamp 1745462530
transform 1 0 600 0 1 1170
box -8 -3 16 105
use FILL  FILL_3999
timestamp 1745462530
transform 1 0 592 0 1 1170
box -8 -3 16 105
use FILL  FILL_4000
timestamp 1745462530
transform 1 0 560 0 1 1170
box -8 -3 16 105
use FILL  FILL_4001
timestamp 1745462530
transform 1 0 552 0 1 1170
box -8 -3 16 105
use FILL  FILL_4002
timestamp 1745462530
transform 1 0 544 0 1 1170
box -8 -3 16 105
use FILL  FILL_4003
timestamp 1745462530
transform 1 0 496 0 1 1170
box -8 -3 16 105
use FILL  FILL_4004
timestamp 1745462530
transform 1 0 488 0 1 1170
box -8 -3 16 105
use FILL  FILL_4005
timestamp 1745462530
transform 1 0 480 0 1 1170
box -8 -3 16 105
use FILL  FILL_4006
timestamp 1745462530
transform 1 0 472 0 1 1170
box -8 -3 16 105
use FILL  FILL_4007
timestamp 1745462530
transform 1 0 448 0 1 1170
box -8 -3 16 105
use FILL  FILL_4008
timestamp 1745462530
transform 1 0 440 0 1 1170
box -8 -3 16 105
use FILL  FILL_4009
timestamp 1745462530
transform 1 0 392 0 1 1170
box -8 -3 16 105
use FILL  FILL_4010
timestamp 1745462530
transform 1 0 384 0 1 1170
box -8 -3 16 105
use FILL  FILL_4011
timestamp 1745462530
transform 1 0 376 0 1 1170
box -8 -3 16 105
use FILL  FILL_4012
timestamp 1745462530
transform 1 0 352 0 1 1170
box -8 -3 16 105
use FILL  FILL_4013
timestamp 1745462530
transform 1 0 344 0 1 1170
box -8 -3 16 105
use FILL  FILL_4014
timestamp 1745462530
transform 1 0 296 0 1 1170
box -8 -3 16 105
use FILL  FILL_4015
timestamp 1745462530
transform 1 0 288 0 1 1170
box -8 -3 16 105
use FILL  FILL_4016
timestamp 1745462530
transform 1 0 280 0 1 1170
box -8 -3 16 105
use FILL  FILL_4017
timestamp 1745462530
transform 1 0 272 0 1 1170
box -8 -3 16 105
use FILL  FILL_4018
timestamp 1745462530
transform 1 0 264 0 1 1170
box -8 -3 16 105
use FILL  FILL_4019
timestamp 1745462530
transform 1 0 240 0 1 1170
box -8 -3 16 105
use FILL  FILL_4020
timestamp 1745462530
transform 1 0 232 0 1 1170
box -8 -3 16 105
use FILL  FILL_4021
timestamp 1745462530
transform 1 0 224 0 1 1170
box -8 -3 16 105
use FILL  FILL_4022
timestamp 1745462530
transform 1 0 216 0 1 1170
box -8 -3 16 105
use FILL  FILL_4023
timestamp 1745462530
transform 1 0 208 0 1 1170
box -8 -3 16 105
use FILL  FILL_4024
timestamp 1745462530
transform 1 0 200 0 1 1170
box -8 -3 16 105
use FILL  FILL_4025
timestamp 1745462530
transform 1 0 96 0 1 1170
box -8 -3 16 105
use FILL  FILL_4026
timestamp 1745462530
transform 1 0 88 0 1 1170
box -8 -3 16 105
use FILL  FILL_4027
timestamp 1745462530
transform 1 0 80 0 1 1170
box -8 -3 16 105
use FILL  FILL_4028
timestamp 1745462530
transform 1 0 72 0 1 1170
box -8 -3 16 105
use FILL  FILL_4029
timestamp 1745462530
transform 1 0 4368 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4030
timestamp 1745462530
transform 1 0 4168 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4031
timestamp 1745462530
transform 1 0 4160 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4032
timestamp 1745462530
transform 1 0 4096 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4033
timestamp 1745462530
transform 1 0 4088 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4034
timestamp 1745462530
transform 1 0 4032 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4035
timestamp 1745462530
transform 1 0 4024 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4036
timestamp 1745462530
transform 1 0 4016 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4037
timestamp 1745462530
transform 1 0 3968 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4038
timestamp 1745462530
transform 1 0 3920 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4039
timestamp 1745462530
transform 1 0 3912 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4040
timestamp 1745462530
transform 1 0 3904 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4041
timestamp 1745462530
transform 1 0 3856 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4042
timestamp 1745462530
transform 1 0 3848 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4043
timestamp 1745462530
transform 1 0 3800 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4044
timestamp 1745462530
transform 1 0 3792 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4045
timestamp 1745462530
transform 1 0 3688 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4046
timestamp 1745462530
transform 1 0 3680 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4047
timestamp 1745462530
transform 1 0 3576 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4048
timestamp 1745462530
transform 1 0 3568 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4049
timestamp 1745462530
transform 1 0 3464 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4050
timestamp 1745462530
transform 1 0 3424 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4051
timestamp 1745462530
transform 1 0 3416 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4052
timestamp 1745462530
transform 1 0 3408 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4053
timestamp 1745462530
transform 1 0 3368 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4054
timestamp 1745462530
transform 1 0 3336 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4055
timestamp 1745462530
transform 1 0 3328 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4056
timestamp 1745462530
transform 1 0 3320 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4057
timestamp 1745462530
transform 1 0 3272 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4058
timestamp 1745462530
transform 1 0 3264 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4059
timestamp 1745462530
transform 1 0 3232 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4060
timestamp 1745462530
transform 1 0 3200 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4061
timestamp 1745462530
transform 1 0 3192 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4062
timestamp 1745462530
transform 1 0 3120 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4063
timestamp 1745462530
transform 1 0 3112 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4064
timestamp 1745462530
transform 1 0 3104 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4065
timestamp 1745462530
transform 1 0 3032 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4066
timestamp 1745462530
transform 1 0 3024 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4067
timestamp 1745462530
transform 1 0 2976 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4068
timestamp 1745462530
transform 1 0 2816 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4069
timestamp 1745462530
transform 1 0 2808 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4070
timestamp 1745462530
transform 1 0 2776 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4071
timestamp 1745462530
transform 1 0 2728 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4072
timestamp 1745462530
transform 1 0 2704 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4073
timestamp 1745462530
transform 1 0 2656 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4074
timestamp 1745462530
transform 1 0 2632 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4075
timestamp 1745462530
transform 1 0 2584 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4076
timestamp 1745462530
transform 1 0 2576 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4077
timestamp 1745462530
transform 1 0 2512 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4078
timestamp 1745462530
transform 1 0 2504 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4079
timestamp 1745462530
transform 1 0 2472 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4080
timestamp 1745462530
transform 1 0 2464 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4081
timestamp 1745462530
transform 1 0 2432 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4082
timestamp 1745462530
transform 1 0 2424 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4083
timestamp 1745462530
transform 1 0 2400 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4084
timestamp 1745462530
transform 1 0 2392 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4085
timestamp 1745462530
transform 1 0 2344 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4086
timestamp 1745462530
transform 1 0 2336 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4087
timestamp 1745462530
transform 1 0 2328 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4088
timestamp 1745462530
transform 1 0 2280 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4089
timestamp 1745462530
transform 1 0 2272 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4090
timestamp 1745462530
transform 1 0 2264 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4091
timestamp 1745462530
transform 1 0 2240 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4092
timestamp 1745462530
transform 1 0 2136 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4093
timestamp 1745462530
transform 1 0 2112 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4094
timestamp 1745462530
transform 1 0 2104 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4095
timestamp 1745462530
transform 1 0 2096 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4096
timestamp 1745462530
transform 1 0 2048 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4097
timestamp 1745462530
transform 1 0 2040 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4098
timestamp 1745462530
transform 1 0 2032 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4099
timestamp 1745462530
transform 1 0 1984 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4100
timestamp 1745462530
transform 1 0 1976 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4101
timestamp 1745462530
transform 1 0 1872 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4102
timestamp 1745462530
transform 1 0 1864 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4103
timestamp 1745462530
transform 1 0 1856 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4104
timestamp 1745462530
transform 1 0 1808 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4105
timestamp 1745462530
transform 1 0 1800 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4106
timestamp 1745462530
transform 1 0 1768 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4107
timestamp 1745462530
transform 1 0 1760 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4108
timestamp 1745462530
transform 1 0 1752 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4109
timestamp 1745462530
transform 1 0 1704 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4110
timestamp 1745462530
transform 1 0 1696 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4111
timestamp 1745462530
transform 1 0 1688 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4112
timestamp 1745462530
transform 1 0 1680 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4113
timestamp 1745462530
transform 1 0 1648 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4114
timestamp 1745462530
transform 1 0 1640 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4115
timestamp 1745462530
transform 1 0 1536 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4116
timestamp 1745462530
transform 1 0 1528 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4117
timestamp 1745462530
transform 1 0 1496 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4118
timestamp 1745462530
transform 1 0 1488 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4119
timestamp 1745462530
transform 1 0 1480 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4120
timestamp 1745462530
transform 1 0 1440 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4121
timestamp 1745462530
transform 1 0 1432 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4122
timestamp 1745462530
transform 1 0 1424 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4123
timestamp 1745462530
transform 1 0 1416 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4124
timestamp 1745462530
transform 1 0 1384 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4125
timestamp 1745462530
transform 1 0 1376 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4126
timestamp 1745462530
transform 1 0 1272 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4127
timestamp 1745462530
transform 1 0 1264 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4128
timestamp 1745462530
transform 1 0 1256 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4129
timestamp 1745462530
transform 1 0 1216 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4130
timestamp 1745462530
transform 1 0 1208 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4131
timestamp 1745462530
transform 1 0 1200 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4132
timestamp 1745462530
transform 1 0 1168 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4133
timestamp 1745462530
transform 1 0 1136 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4134
timestamp 1745462530
transform 1 0 1128 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4135
timestamp 1745462530
transform 1 0 1120 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4136
timestamp 1745462530
transform 1 0 1072 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4137
timestamp 1745462530
transform 1 0 1064 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4138
timestamp 1745462530
transform 1 0 1056 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4139
timestamp 1745462530
transform 1 0 1048 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4140
timestamp 1745462530
transform 1 0 1016 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4141
timestamp 1745462530
transform 1 0 1008 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4142
timestamp 1745462530
transform 1 0 968 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4143
timestamp 1745462530
transform 1 0 960 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4144
timestamp 1745462530
transform 1 0 928 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4145
timestamp 1745462530
transform 1 0 920 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4146
timestamp 1745462530
transform 1 0 912 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4147
timestamp 1745462530
transform 1 0 864 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4148
timestamp 1745462530
transform 1 0 856 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4149
timestamp 1745462530
transform 1 0 848 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4150
timestamp 1745462530
transform 1 0 800 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4151
timestamp 1745462530
transform 1 0 792 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4152
timestamp 1745462530
transform 1 0 784 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4153
timestamp 1745462530
transform 1 0 776 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4154
timestamp 1745462530
transform 1 0 728 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4155
timestamp 1745462530
transform 1 0 720 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4156
timestamp 1745462530
transform 1 0 712 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4157
timestamp 1745462530
transform 1 0 664 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4158
timestamp 1745462530
transform 1 0 656 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4159
timestamp 1745462530
transform 1 0 648 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4160
timestamp 1745462530
transform 1 0 616 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4161
timestamp 1745462530
transform 1 0 608 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4162
timestamp 1745462530
transform 1 0 600 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4163
timestamp 1745462530
transform 1 0 552 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4164
timestamp 1745462530
transform 1 0 544 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4165
timestamp 1745462530
transform 1 0 536 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4166
timestamp 1745462530
transform 1 0 432 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4167
timestamp 1745462530
transform 1 0 424 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4168
timestamp 1745462530
transform 1 0 360 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4169
timestamp 1745462530
transform 1 0 352 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4170
timestamp 1745462530
transform 1 0 344 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4171
timestamp 1745462530
transform 1 0 240 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4172
timestamp 1745462530
transform 1 0 232 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4173
timestamp 1745462530
transform 1 0 224 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4174
timestamp 1745462530
transform 1 0 176 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4175
timestamp 1745462530
transform 1 0 168 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4176
timestamp 1745462530
transform 1 0 160 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4177
timestamp 1745462530
transform 1 0 136 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4178
timestamp 1745462530
transform 1 0 128 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4179
timestamp 1745462530
transform 1 0 120 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4180
timestamp 1745462530
transform 1 0 112 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4181
timestamp 1745462530
transform 1 0 104 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4182
timestamp 1745462530
transform 1 0 96 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4183
timestamp 1745462530
transform 1 0 88 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4184
timestamp 1745462530
transform 1 0 80 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4185
timestamp 1745462530
transform 1 0 72 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4186
timestamp 1745462530
transform 1 0 4352 0 1 970
box -8 -3 16 105
use FILL  FILL_4187
timestamp 1745462530
transform 1 0 4344 0 1 970
box -8 -3 16 105
use FILL  FILL_4188
timestamp 1745462530
transform 1 0 4336 0 1 970
box -8 -3 16 105
use FILL  FILL_4189
timestamp 1745462530
transform 1 0 4288 0 1 970
box -8 -3 16 105
use FILL  FILL_4190
timestamp 1745462530
transform 1 0 4280 0 1 970
box -8 -3 16 105
use FILL  FILL_4191
timestamp 1745462530
transform 1 0 4272 0 1 970
box -8 -3 16 105
use FILL  FILL_4192
timestamp 1745462530
transform 1 0 4248 0 1 970
box -8 -3 16 105
use FILL  FILL_4193
timestamp 1745462530
transform 1 0 4200 0 1 970
box -8 -3 16 105
use FILL  FILL_4194
timestamp 1745462530
transform 1 0 4192 0 1 970
box -8 -3 16 105
use FILL  FILL_4195
timestamp 1745462530
transform 1 0 4184 0 1 970
box -8 -3 16 105
use FILL  FILL_4196
timestamp 1745462530
transform 1 0 4136 0 1 970
box -8 -3 16 105
use FILL  FILL_4197
timestamp 1745462530
transform 1 0 4096 0 1 970
box -8 -3 16 105
use FILL  FILL_4198
timestamp 1745462530
transform 1 0 4088 0 1 970
box -8 -3 16 105
use FILL  FILL_4199
timestamp 1745462530
transform 1 0 4080 0 1 970
box -8 -3 16 105
use FILL  FILL_4200
timestamp 1745462530
transform 1 0 4032 0 1 970
box -8 -3 16 105
use FILL  FILL_4201
timestamp 1745462530
transform 1 0 4024 0 1 970
box -8 -3 16 105
use FILL  FILL_4202
timestamp 1745462530
transform 1 0 4016 0 1 970
box -8 -3 16 105
use FILL  FILL_4203
timestamp 1745462530
transform 1 0 3968 0 1 970
box -8 -3 16 105
use FILL  FILL_4204
timestamp 1745462530
transform 1 0 3960 0 1 970
box -8 -3 16 105
use FILL  FILL_4205
timestamp 1745462530
transform 1 0 3952 0 1 970
box -8 -3 16 105
use FILL  FILL_4206
timestamp 1745462530
transform 1 0 3904 0 1 970
box -8 -3 16 105
use FILL  FILL_4207
timestamp 1745462530
transform 1 0 3896 0 1 970
box -8 -3 16 105
use FILL  FILL_4208
timestamp 1745462530
transform 1 0 3888 0 1 970
box -8 -3 16 105
use FILL  FILL_4209
timestamp 1745462530
transform 1 0 3848 0 1 970
box -8 -3 16 105
use FILL  FILL_4210
timestamp 1745462530
transform 1 0 3840 0 1 970
box -8 -3 16 105
use FILL  FILL_4211
timestamp 1745462530
transform 1 0 3832 0 1 970
box -8 -3 16 105
use FILL  FILL_4212
timestamp 1745462530
transform 1 0 3784 0 1 970
box -8 -3 16 105
use FILL  FILL_4213
timestamp 1745462530
transform 1 0 3776 0 1 970
box -8 -3 16 105
use FILL  FILL_4214
timestamp 1745462530
transform 1 0 3768 0 1 970
box -8 -3 16 105
use FILL  FILL_4215
timestamp 1745462530
transform 1 0 3720 0 1 970
box -8 -3 16 105
use FILL  FILL_4216
timestamp 1745462530
transform 1 0 3712 0 1 970
box -8 -3 16 105
use FILL  FILL_4217
timestamp 1745462530
transform 1 0 3704 0 1 970
box -8 -3 16 105
use FILL  FILL_4218
timestamp 1745462530
transform 1 0 3656 0 1 970
box -8 -3 16 105
use FILL  FILL_4219
timestamp 1745462530
transform 1 0 3648 0 1 970
box -8 -3 16 105
use FILL  FILL_4220
timestamp 1745462530
transform 1 0 3640 0 1 970
box -8 -3 16 105
use FILL  FILL_4221
timestamp 1745462530
transform 1 0 3592 0 1 970
box -8 -3 16 105
use FILL  FILL_4222
timestamp 1745462530
transform 1 0 3584 0 1 970
box -8 -3 16 105
use FILL  FILL_4223
timestamp 1745462530
transform 1 0 3576 0 1 970
box -8 -3 16 105
use FILL  FILL_4224
timestamp 1745462530
transform 1 0 3568 0 1 970
box -8 -3 16 105
use FILL  FILL_4225
timestamp 1745462530
transform 1 0 3520 0 1 970
box -8 -3 16 105
use FILL  FILL_4226
timestamp 1745462530
transform 1 0 3512 0 1 970
box -8 -3 16 105
use FILL  FILL_4227
timestamp 1745462530
transform 1 0 3488 0 1 970
box -8 -3 16 105
use FILL  FILL_4228
timestamp 1745462530
transform 1 0 3480 0 1 970
box -8 -3 16 105
use FILL  FILL_4229
timestamp 1745462530
transform 1 0 3432 0 1 970
box -8 -3 16 105
use FILL  FILL_4230
timestamp 1745462530
transform 1 0 3424 0 1 970
box -8 -3 16 105
use FILL  FILL_4231
timestamp 1745462530
transform 1 0 3416 0 1 970
box -8 -3 16 105
use FILL  FILL_4232
timestamp 1745462530
transform 1 0 3368 0 1 970
box -8 -3 16 105
use FILL  FILL_4233
timestamp 1745462530
transform 1 0 3360 0 1 970
box -8 -3 16 105
use FILL  FILL_4234
timestamp 1745462530
transform 1 0 3352 0 1 970
box -8 -3 16 105
use FILL  FILL_4235
timestamp 1745462530
transform 1 0 3304 0 1 970
box -8 -3 16 105
use FILL  FILL_4236
timestamp 1745462530
transform 1 0 3280 0 1 970
box -8 -3 16 105
use FILL  FILL_4237
timestamp 1745462530
transform 1 0 3272 0 1 970
box -8 -3 16 105
use FILL  FILL_4238
timestamp 1745462530
transform 1 0 3232 0 1 970
box -8 -3 16 105
use FILL  FILL_4239
timestamp 1745462530
transform 1 0 3224 0 1 970
box -8 -3 16 105
use FILL  FILL_4240
timestamp 1745462530
transform 1 0 3192 0 1 970
box -8 -3 16 105
use FILL  FILL_4241
timestamp 1745462530
transform 1 0 3184 0 1 970
box -8 -3 16 105
use FILL  FILL_4242
timestamp 1745462530
transform 1 0 3144 0 1 970
box -8 -3 16 105
use FILL  FILL_4243
timestamp 1745462530
transform 1 0 3136 0 1 970
box -8 -3 16 105
use FILL  FILL_4244
timestamp 1745462530
transform 1 0 3088 0 1 970
box -8 -3 16 105
use FILL  FILL_4245
timestamp 1745462530
transform 1 0 3080 0 1 970
box -8 -3 16 105
use FILL  FILL_4246
timestamp 1745462530
transform 1 0 3072 0 1 970
box -8 -3 16 105
use FILL  FILL_4247
timestamp 1745462530
transform 1 0 3024 0 1 970
box -8 -3 16 105
use FILL  FILL_4248
timestamp 1745462530
transform 1 0 3016 0 1 970
box -8 -3 16 105
use FILL  FILL_4249
timestamp 1745462530
transform 1 0 3008 0 1 970
box -8 -3 16 105
use FILL  FILL_4250
timestamp 1745462530
transform 1 0 2968 0 1 970
box -8 -3 16 105
use FILL  FILL_4251
timestamp 1745462530
transform 1 0 2944 0 1 970
box -8 -3 16 105
use FILL  FILL_4252
timestamp 1745462530
transform 1 0 2936 0 1 970
box -8 -3 16 105
use FILL  FILL_4253
timestamp 1745462530
transform 1 0 2888 0 1 970
box -8 -3 16 105
use FILL  FILL_4254
timestamp 1745462530
transform 1 0 2880 0 1 970
box -8 -3 16 105
use FILL  FILL_4255
timestamp 1745462530
transform 1 0 2872 0 1 970
box -8 -3 16 105
use FILL  FILL_4256
timestamp 1745462530
transform 1 0 2832 0 1 970
box -8 -3 16 105
use FILL  FILL_4257
timestamp 1745462530
transform 1 0 2824 0 1 970
box -8 -3 16 105
use FILL  FILL_4258
timestamp 1745462530
transform 1 0 2784 0 1 970
box -8 -3 16 105
use FILL  FILL_4259
timestamp 1745462530
transform 1 0 2776 0 1 970
box -8 -3 16 105
use FILL  FILL_4260
timestamp 1745462530
transform 1 0 2752 0 1 970
box -8 -3 16 105
use FILL  FILL_4261
timestamp 1745462530
transform 1 0 2720 0 1 970
box -8 -3 16 105
use FILL  FILL_4262
timestamp 1745462530
transform 1 0 2712 0 1 970
box -8 -3 16 105
use FILL  FILL_4263
timestamp 1745462530
transform 1 0 2704 0 1 970
box -8 -3 16 105
use FILL  FILL_4264
timestamp 1745462530
transform 1 0 2672 0 1 970
box -8 -3 16 105
use FILL  FILL_4265
timestamp 1745462530
transform 1 0 2664 0 1 970
box -8 -3 16 105
use FILL  FILL_4266
timestamp 1745462530
transform 1 0 2656 0 1 970
box -8 -3 16 105
use FILL  FILL_4267
timestamp 1745462530
transform 1 0 2552 0 1 970
box -8 -3 16 105
use FILL  FILL_4268
timestamp 1745462530
transform 1 0 2544 0 1 970
box -8 -3 16 105
use FILL  FILL_4269
timestamp 1745462530
transform 1 0 2536 0 1 970
box -8 -3 16 105
use FILL  FILL_4270
timestamp 1745462530
transform 1 0 2488 0 1 970
box -8 -3 16 105
use FILL  FILL_4271
timestamp 1745462530
transform 1 0 2480 0 1 970
box -8 -3 16 105
use FILL  FILL_4272
timestamp 1745462530
transform 1 0 2472 0 1 970
box -8 -3 16 105
use FILL  FILL_4273
timestamp 1745462530
transform 1 0 2464 0 1 970
box -8 -3 16 105
use FILL  FILL_4274
timestamp 1745462530
transform 1 0 2416 0 1 970
box -8 -3 16 105
use FILL  FILL_4275
timestamp 1745462530
transform 1 0 2408 0 1 970
box -8 -3 16 105
use FILL  FILL_4276
timestamp 1745462530
transform 1 0 2400 0 1 970
box -8 -3 16 105
use FILL  FILL_4277
timestamp 1745462530
transform 1 0 2352 0 1 970
box -8 -3 16 105
use FILL  FILL_4278
timestamp 1745462530
transform 1 0 2344 0 1 970
box -8 -3 16 105
use FILL  FILL_4279
timestamp 1745462530
transform 1 0 2336 0 1 970
box -8 -3 16 105
use FILL  FILL_4280
timestamp 1745462530
transform 1 0 2328 0 1 970
box -8 -3 16 105
use FILL  FILL_4281
timestamp 1745462530
transform 1 0 2288 0 1 970
box -8 -3 16 105
use FILL  FILL_4282
timestamp 1745462530
transform 1 0 2280 0 1 970
box -8 -3 16 105
use FILL  FILL_4283
timestamp 1745462530
transform 1 0 2248 0 1 970
box -8 -3 16 105
use FILL  FILL_4284
timestamp 1745462530
transform 1 0 2240 0 1 970
box -8 -3 16 105
use FILL  FILL_4285
timestamp 1745462530
transform 1 0 2232 0 1 970
box -8 -3 16 105
use FILL  FILL_4286
timestamp 1745462530
transform 1 0 2184 0 1 970
box -8 -3 16 105
use FILL  FILL_4287
timestamp 1745462530
transform 1 0 2176 0 1 970
box -8 -3 16 105
use FILL  FILL_4288
timestamp 1745462530
transform 1 0 2168 0 1 970
box -8 -3 16 105
use FILL  FILL_4289
timestamp 1745462530
transform 1 0 2160 0 1 970
box -8 -3 16 105
use FILL  FILL_4290
timestamp 1745462530
transform 1 0 2112 0 1 970
box -8 -3 16 105
use FILL  FILL_4291
timestamp 1745462530
transform 1 0 2104 0 1 970
box -8 -3 16 105
use FILL  FILL_4292
timestamp 1745462530
transform 1 0 2072 0 1 970
box -8 -3 16 105
use FILL  FILL_4293
timestamp 1745462530
transform 1 0 2064 0 1 970
box -8 -3 16 105
use FILL  FILL_4294
timestamp 1745462530
transform 1 0 2056 0 1 970
box -8 -3 16 105
use FILL  FILL_4295
timestamp 1745462530
transform 1 0 2008 0 1 970
box -8 -3 16 105
use FILL  FILL_4296
timestamp 1745462530
transform 1 0 1984 0 1 970
box -8 -3 16 105
use FILL  FILL_4297
timestamp 1745462530
transform 1 0 1880 0 1 970
box -8 -3 16 105
use FILL  FILL_4298
timestamp 1745462530
transform 1 0 1832 0 1 970
box -8 -3 16 105
use FILL  FILL_4299
timestamp 1745462530
transform 1 0 1824 0 1 970
box -8 -3 16 105
use FILL  FILL_4300
timestamp 1745462530
transform 1 0 1816 0 1 970
box -8 -3 16 105
use FILL  FILL_4301
timestamp 1745462530
transform 1 0 1752 0 1 970
box -8 -3 16 105
use FILL  FILL_4302
timestamp 1745462530
transform 1 0 1744 0 1 970
box -8 -3 16 105
use FILL  FILL_4303
timestamp 1745462530
transform 1 0 1736 0 1 970
box -8 -3 16 105
use FILL  FILL_4304
timestamp 1745462530
transform 1 0 1688 0 1 970
box -8 -3 16 105
use FILL  FILL_4305
timestamp 1745462530
transform 1 0 1680 0 1 970
box -8 -3 16 105
use FILL  FILL_4306
timestamp 1745462530
transform 1 0 1640 0 1 970
box -8 -3 16 105
use FILL  FILL_4307
timestamp 1745462530
transform 1 0 1608 0 1 970
box -8 -3 16 105
use FILL  FILL_4308
timestamp 1745462530
transform 1 0 1576 0 1 970
box -8 -3 16 105
use FILL  FILL_4309
timestamp 1745462530
transform 1 0 1568 0 1 970
box -8 -3 16 105
use FILL  FILL_4310
timestamp 1745462530
transform 1 0 1560 0 1 970
box -8 -3 16 105
use FILL  FILL_4311
timestamp 1745462530
transform 1 0 1512 0 1 970
box -8 -3 16 105
use FILL  FILL_4312
timestamp 1745462530
transform 1 0 1504 0 1 970
box -8 -3 16 105
use FILL  FILL_4313
timestamp 1745462530
transform 1 0 1496 0 1 970
box -8 -3 16 105
use FILL  FILL_4314
timestamp 1745462530
transform 1 0 1456 0 1 970
box -8 -3 16 105
use FILL  FILL_4315
timestamp 1745462530
transform 1 0 1448 0 1 970
box -8 -3 16 105
use FILL  FILL_4316
timestamp 1745462530
transform 1 0 1400 0 1 970
box -8 -3 16 105
use FILL  FILL_4317
timestamp 1745462530
transform 1 0 1392 0 1 970
box -8 -3 16 105
use FILL  FILL_4318
timestamp 1745462530
transform 1 0 1384 0 1 970
box -8 -3 16 105
use FILL  FILL_4319
timestamp 1745462530
transform 1 0 1264 0 1 970
box -8 -3 16 105
use FILL  FILL_4320
timestamp 1745462530
transform 1 0 1256 0 1 970
box -8 -3 16 105
use FILL  FILL_4321
timestamp 1745462530
transform 1 0 1208 0 1 970
box -8 -3 16 105
use FILL  FILL_4322
timestamp 1745462530
transform 1 0 1200 0 1 970
box -8 -3 16 105
use FILL  FILL_4323
timestamp 1745462530
transform 1 0 1192 0 1 970
box -8 -3 16 105
use FILL  FILL_4324
timestamp 1745462530
transform 1 0 1144 0 1 970
box -8 -3 16 105
use FILL  FILL_4325
timestamp 1745462530
transform 1 0 1136 0 1 970
box -8 -3 16 105
use FILL  FILL_4326
timestamp 1745462530
transform 1 0 1128 0 1 970
box -8 -3 16 105
use FILL  FILL_4327
timestamp 1745462530
transform 1 0 1088 0 1 970
box -8 -3 16 105
use FILL  FILL_4328
timestamp 1745462530
transform 1 0 1056 0 1 970
box -8 -3 16 105
use FILL  FILL_4329
timestamp 1745462530
transform 1 0 1048 0 1 970
box -8 -3 16 105
use FILL  FILL_4330
timestamp 1745462530
transform 1 0 1000 0 1 970
box -8 -3 16 105
use FILL  FILL_4331
timestamp 1745462530
transform 1 0 992 0 1 970
box -8 -3 16 105
use FILL  FILL_4332
timestamp 1745462530
transform 1 0 984 0 1 970
box -8 -3 16 105
use FILL  FILL_4333
timestamp 1745462530
transform 1 0 952 0 1 970
box -8 -3 16 105
use FILL  FILL_4334
timestamp 1745462530
transform 1 0 912 0 1 970
box -8 -3 16 105
use FILL  FILL_4335
timestamp 1745462530
transform 1 0 904 0 1 970
box -8 -3 16 105
use FILL  FILL_4336
timestamp 1745462530
transform 1 0 856 0 1 970
box -8 -3 16 105
use FILL  FILL_4337
timestamp 1745462530
transform 1 0 848 0 1 970
box -8 -3 16 105
use FILL  FILL_4338
timestamp 1745462530
transform 1 0 840 0 1 970
box -8 -3 16 105
use FILL  FILL_4339
timestamp 1745462530
transform 1 0 776 0 1 970
box -8 -3 16 105
use FILL  FILL_4340
timestamp 1745462530
transform 1 0 768 0 1 970
box -8 -3 16 105
use FILL  FILL_4341
timestamp 1745462530
transform 1 0 760 0 1 970
box -8 -3 16 105
use FILL  FILL_4342
timestamp 1745462530
transform 1 0 752 0 1 970
box -8 -3 16 105
use FILL  FILL_4343
timestamp 1745462530
transform 1 0 704 0 1 970
box -8 -3 16 105
use FILL  FILL_4344
timestamp 1745462530
transform 1 0 696 0 1 970
box -8 -3 16 105
use FILL  FILL_4345
timestamp 1745462530
transform 1 0 656 0 1 970
box -8 -3 16 105
use FILL  FILL_4346
timestamp 1745462530
transform 1 0 624 0 1 970
box -8 -3 16 105
use FILL  FILL_4347
timestamp 1745462530
transform 1 0 616 0 1 970
box -8 -3 16 105
use FILL  FILL_4348
timestamp 1745462530
transform 1 0 608 0 1 970
box -8 -3 16 105
use FILL  FILL_4349
timestamp 1745462530
transform 1 0 560 0 1 970
box -8 -3 16 105
use FILL  FILL_4350
timestamp 1745462530
transform 1 0 552 0 1 970
box -8 -3 16 105
use FILL  FILL_4351
timestamp 1745462530
transform 1 0 448 0 1 970
box -8 -3 16 105
use FILL  FILL_4352
timestamp 1745462530
transform 1 0 440 0 1 970
box -8 -3 16 105
use FILL  FILL_4353
timestamp 1745462530
transform 1 0 400 0 1 970
box -8 -3 16 105
use FILL  FILL_4354
timestamp 1745462530
transform 1 0 352 0 1 970
box -8 -3 16 105
use FILL  FILL_4355
timestamp 1745462530
transform 1 0 344 0 1 970
box -8 -3 16 105
use FILL  FILL_4356
timestamp 1745462530
transform 1 0 312 0 1 970
box -8 -3 16 105
use FILL  FILL_4357
timestamp 1745462530
transform 1 0 264 0 1 970
box -8 -3 16 105
use FILL  FILL_4358
timestamp 1745462530
transform 1 0 256 0 1 970
box -8 -3 16 105
use FILL  FILL_4359
timestamp 1745462530
transform 1 0 248 0 1 970
box -8 -3 16 105
use FILL  FILL_4360
timestamp 1745462530
transform 1 0 184 0 1 970
box -8 -3 16 105
use FILL  FILL_4361
timestamp 1745462530
transform 1 0 176 0 1 970
box -8 -3 16 105
use FILL  FILL_4362
timestamp 1745462530
transform 1 0 72 0 1 970
box -8 -3 16 105
use FILL  FILL_4363
timestamp 1745462530
transform 1 0 4272 0 -1 970
box -8 -3 16 105
use FILL  FILL_4364
timestamp 1745462530
transform 1 0 4224 0 -1 970
box -8 -3 16 105
use FILL  FILL_4365
timestamp 1745462530
transform 1 0 4216 0 -1 970
box -8 -3 16 105
use FILL  FILL_4366
timestamp 1745462530
transform 1 0 4208 0 -1 970
box -8 -3 16 105
use FILL  FILL_4367
timestamp 1745462530
transform 1 0 4072 0 -1 970
box -8 -3 16 105
use FILL  FILL_4368
timestamp 1745462530
transform 1 0 4064 0 -1 970
box -8 -3 16 105
use FILL  FILL_4369
timestamp 1745462530
transform 1 0 4024 0 -1 970
box -8 -3 16 105
use FILL  FILL_4370
timestamp 1745462530
transform 1 0 4016 0 -1 970
box -8 -3 16 105
use FILL  FILL_4371
timestamp 1745462530
transform 1 0 4008 0 -1 970
box -8 -3 16 105
use FILL  FILL_4372
timestamp 1745462530
transform 1 0 3968 0 -1 970
box -8 -3 16 105
use FILL  FILL_4373
timestamp 1745462530
transform 1 0 3960 0 -1 970
box -8 -3 16 105
use FILL  FILL_4374
timestamp 1745462530
transform 1 0 3952 0 -1 970
box -8 -3 16 105
use FILL  FILL_4375
timestamp 1745462530
transform 1 0 3904 0 -1 970
box -8 -3 16 105
use FILL  FILL_4376
timestamp 1745462530
transform 1 0 3896 0 -1 970
box -8 -3 16 105
use FILL  FILL_4377
timestamp 1745462530
transform 1 0 3888 0 -1 970
box -8 -3 16 105
use FILL  FILL_4378
timestamp 1745462530
transform 1 0 3848 0 -1 970
box -8 -3 16 105
use FILL  FILL_4379
timestamp 1745462530
transform 1 0 3840 0 -1 970
box -8 -3 16 105
use FILL  FILL_4380
timestamp 1745462530
transform 1 0 3736 0 -1 970
box -8 -3 16 105
use FILL  FILL_4381
timestamp 1745462530
transform 1 0 3728 0 -1 970
box -8 -3 16 105
use FILL  FILL_4382
timestamp 1745462530
transform 1 0 3696 0 -1 970
box -8 -3 16 105
use FILL  FILL_4383
timestamp 1745462530
transform 1 0 3688 0 -1 970
box -8 -3 16 105
use FILL  FILL_4384
timestamp 1745462530
transform 1 0 3680 0 -1 970
box -8 -3 16 105
use FILL  FILL_4385
timestamp 1745462530
transform 1 0 3632 0 -1 970
box -8 -3 16 105
use FILL  FILL_4386
timestamp 1745462530
transform 1 0 3624 0 -1 970
box -8 -3 16 105
use FILL  FILL_4387
timestamp 1745462530
transform 1 0 3616 0 -1 970
box -8 -3 16 105
use FILL  FILL_4388
timestamp 1745462530
transform 1 0 3568 0 -1 970
box -8 -3 16 105
use FILL  FILL_4389
timestamp 1745462530
transform 1 0 3560 0 -1 970
box -8 -3 16 105
use FILL  FILL_4390
timestamp 1745462530
transform 1 0 3528 0 -1 970
box -8 -3 16 105
use FILL  FILL_4391
timestamp 1745462530
transform 1 0 3520 0 -1 970
box -8 -3 16 105
use FILL  FILL_4392
timestamp 1745462530
transform 1 0 3416 0 -1 970
box -8 -3 16 105
use FILL  FILL_4393
timestamp 1745462530
transform 1 0 3408 0 -1 970
box -8 -3 16 105
use FILL  FILL_4394
timestamp 1745462530
transform 1 0 3400 0 -1 970
box -8 -3 16 105
use FILL  FILL_4395
timestamp 1745462530
transform 1 0 3352 0 -1 970
box -8 -3 16 105
use FILL  FILL_4396
timestamp 1745462530
transform 1 0 3344 0 -1 970
box -8 -3 16 105
use FILL  FILL_4397
timestamp 1745462530
transform 1 0 3240 0 -1 970
box -8 -3 16 105
use FILL  FILL_4398
timestamp 1745462530
transform 1 0 3232 0 -1 970
box -8 -3 16 105
use FILL  FILL_4399
timestamp 1745462530
transform 1 0 3224 0 -1 970
box -8 -3 16 105
use FILL  FILL_4400
timestamp 1745462530
transform 1 0 3192 0 -1 970
box -8 -3 16 105
use FILL  FILL_4401
timestamp 1745462530
transform 1 0 3160 0 -1 970
box -8 -3 16 105
use FILL  FILL_4402
timestamp 1745462530
transform 1 0 3152 0 -1 970
box -8 -3 16 105
use FILL  FILL_4403
timestamp 1745462530
transform 1 0 3144 0 -1 970
box -8 -3 16 105
use FILL  FILL_4404
timestamp 1745462530
transform 1 0 3104 0 -1 970
box -8 -3 16 105
use FILL  FILL_4405
timestamp 1745462530
transform 1 0 3096 0 -1 970
box -8 -3 16 105
use FILL  FILL_4406
timestamp 1745462530
transform 1 0 3048 0 -1 970
box -8 -3 16 105
use FILL  FILL_4407
timestamp 1745462530
transform 1 0 3040 0 -1 970
box -8 -3 16 105
use FILL  FILL_4408
timestamp 1745462530
transform 1 0 2936 0 -1 970
box -8 -3 16 105
use FILL  FILL_4409
timestamp 1745462530
transform 1 0 2928 0 -1 970
box -8 -3 16 105
use FILL  FILL_4410
timestamp 1745462530
transform 1 0 2880 0 -1 970
box -8 -3 16 105
use FILL  FILL_4411
timestamp 1745462530
transform 1 0 2872 0 -1 970
box -8 -3 16 105
use FILL  FILL_4412
timestamp 1745462530
transform 1 0 2832 0 -1 970
box -8 -3 16 105
use FILL  FILL_4413
timestamp 1745462530
transform 1 0 2824 0 -1 970
box -8 -3 16 105
use FILL  FILL_4414
timestamp 1745462530
transform 1 0 2776 0 -1 970
box -8 -3 16 105
use FILL  FILL_4415
timestamp 1745462530
transform 1 0 2768 0 -1 970
box -8 -3 16 105
use FILL  FILL_4416
timestamp 1745462530
transform 1 0 2704 0 -1 970
box -8 -3 16 105
use FILL  FILL_4417
timestamp 1745462530
transform 1 0 2696 0 -1 970
box -8 -3 16 105
use FILL  FILL_4418
timestamp 1745462530
transform 1 0 2592 0 -1 970
box -8 -3 16 105
use FILL  FILL_4419
timestamp 1745462530
transform 1 0 2584 0 -1 970
box -8 -3 16 105
use FILL  FILL_4420
timestamp 1745462530
transform 1 0 2536 0 -1 970
box -8 -3 16 105
use FILL  FILL_4421
timestamp 1745462530
transform 1 0 2512 0 -1 970
box -8 -3 16 105
use FILL  FILL_4422
timestamp 1745462530
transform 1 0 2504 0 -1 970
box -8 -3 16 105
use FILL  FILL_4423
timestamp 1745462530
transform 1 0 2456 0 -1 970
box -8 -3 16 105
use FILL  FILL_4424
timestamp 1745462530
transform 1 0 2448 0 -1 970
box -8 -3 16 105
use FILL  FILL_4425
timestamp 1745462530
transform 1 0 2392 0 -1 970
box -8 -3 16 105
use FILL  FILL_4426
timestamp 1745462530
transform 1 0 2384 0 -1 970
box -8 -3 16 105
use FILL  FILL_4427
timestamp 1745462530
transform 1 0 2376 0 -1 970
box -8 -3 16 105
use FILL  FILL_4428
timestamp 1745462530
transform 1 0 2328 0 -1 970
box -8 -3 16 105
use FILL  FILL_4429
timestamp 1745462530
transform 1 0 2320 0 -1 970
box -8 -3 16 105
use FILL  FILL_4430
timestamp 1745462530
transform 1 0 2312 0 -1 970
box -8 -3 16 105
use FILL  FILL_4431
timestamp 1745462530
transform 1 0 2264 0 -1 970
box -8 -3 16 105
use FILL  FILL_4432
timestamp 1745462530
transform 1 0 2256 0 -1 970
box -8 -3 16 105
use FILL  FILL_4433
timestamp 1745462530
transform 1 0 2152 0 -1 970
box -8 -3 16 105
use FILL  FILL_4434
timestamp 1745462530
transform 1 0 2144 0 -1 970
box -8 -3 16 105
use FILL  FILL_4435
timestamp 1745462530
transform 1 0 2040 0 -1 970
box -8 -3 16 105
use FILL  FILL_4436
timestamp 1745462530
transform 1 0 2032 0 -1 970
box -8 -3 16 105
use FILL  FILL_4437
timestamp 1745462530
transform 1 0 1984 0 -1 970
box -8 -3 16 105
use FILL  FILL_4438
timestamp 1745462530
transform 1 0 1976 0 -1 970
box -8 -3 16 105
use FILL  FILL_4439
timestamp 1745462530
transform 1 0 1936 0 -1 970
box -8 -3 16 105
use FILL  FILL_4440
timestamp 1745462530
transform 1 0 1928 0 -1 970
box -8 -3 16 105
use FILL  FILL_4441
timestamp 1745462530
transform 1 0 1880 0 -1 970
box -8 -3 16 105
use FILL  FILL_4442
timestamp 1745462530
transform 1 0 1872 0 -1 970
box -8 -3 16 105
use FILL  FILL_4443
timestamp 1745462530
transform 1 0 1832 0 -1 970
box -8 -3 16 105
use FILL  FILL_4444
timestamp 1745462530
transform 1 0 1728 0 -1 970
box -8 -3 16 105
use FILL  FILL_4445
timestamp 1745462530
transform 1 0 1696 0 -1 970
box -8 -3 16 105
use FILL  FILL_4446
timestamp 1745462530
transform 1 0 1688 0 -1 970
box -8 -3 16 105
use FILL  FILL_4447
timestamp 1745462530
transform 1 0 1640 0 -1 970
box -8 -3 16 105
use FILL  FILL_4448
timestamp 1745462530
transform 1 0 1632 0 -1 970
box -8 -3 16 105
use FILL  FILL_4449
timestamp 1745462530
transform 1 0 1624 0 -1 970
box -8 -3 16 105
use FILL  FILL_4450
timestamp 1745462530
transform 1 0 1576 0 -1 970
box -8 -3 16 105
use FILL  FILL_4451
timestamp 1745462530
transform 1 0 1568 0 -1 970
box -8 -3 16 105
use FILL  FILL_4452
timestamp 1745462530
transform 1 0 1544 0 -1 970
box -8 -3 16 105
use FILL  FILL_4453
timestamp 1745462530
transform 1 0 1512 0 -1 970
box -8 -3 16 105
use FILL  FILL_4454
timestamp 1745462530
transform 1 0 1504 0 -1 970
box -8 -3 16 105
use FILL  FILL_4455
timestamp 1745462530
transform 1 0 1464 0 -1 970
box -8 -3 16 105
use FILL  FILL_4456
timestamp 1745462530
transform 1 0 1456 0 -1 970
box -8 -3 16 105
use FILL  FILL_4457
timestamp 1745462530
transform 1 0 1448 0 -1 970
box -8 -3 16 105
use FILL  FILL_4458
timestamp 1745462530
transform 1 0 1400 0 -1 970
box -8 -3 16 105
use FILL  FILL_4459
timestamp 1745462530
transform 1 0 1392 0 -1 970
box -8 -3 16 105
use FILL  FILL_4460
timestamp 1745462530
transform 1 0 1384 0 -1 970
box -8 -3 16 105
use FILL  FILL_4461
timestamp 1745462530
transform 1 0 1264 0 -1 970
box -8 -3 16 105
use FILL  FILL_4462
timestamp 1745462530
transform 1 0 1256 0 -1 970
box -8 -3 16 105
use FILL  FILL_4463
timestamp 1745462530
transform 1 0 1208 0 -1 970
box -8 -3 16 105
use FILL  FILL_4464
timestamp 1745462530
transform 1 0 1200 0 -1 970
box -8 -3 16 105
use FILL  FILL_4465
timestamp 1745462530
transform 1 0 1192 0 -1 970
box -8 -3 16 105
use FILL  FILL_4466
timestamp 1745462530
transform 1 0 1152 0 -1 970
box -8 -3 16 105
use FILL  FILL_4467
timestamp 1745462530
transform 1 0 1144 0 -1 970
box -8 -3 16 105
use FILL  FILL_4468
timestamp 1745462530
transform 1 0 1112 0 -1 970
box -8 -3 16 105
use FILL  FILL_4469
timestamp 1745462530
transform 1 0 1104 0 -1 970
box -8 -3 16 105
use FILL  FILL_4470
timestamp 1745462530
transform 1 0 1064 0 -1 970
box -8 -3 16 105
use FILL  FILL_4471
timestamp 1745462530
transform 1 0 1056 0 -1 970
box -8 -3 16 105
use FILL  FILL_4472
timestamp 1745462530
transform 1 0 1048 0 -1 970
box -8 -3 16 105
use FILL  FILL_4473
timestamp 1745462530
transform 1 0 1000 0 -1 970
box -8 -3 16 105
use FILL  FILL_4474
timestamp 1745462530
transform 1 0 992 0 -1 970
box -8 -3 16 105
use FILL  FILL_4475
timestamp 1745462530
transform 1 0 984 0 -1 970
box -8 -3 16 105
use FILL  FILL_4476
timestamp 1745462530
transform 1 0 936 0 -1 970
box -8 -3 16 105
use FILL  FILL_4477
timestamp 1745462530
transform 1 0 928 0 -1 970
box -8 -3 16 105
use FILL  FILL_4478
timestamp 1745462530
transform 1 0 920 0 -1 970
box -8 -3 16 105
use FILL  FILL_4479
timestamp 1745462530
transform 1 0 872 0 -1 970
box -8 -3 16 105
use FILL  FILL_4480
timestamp 1745462530
transform 1 0 864 0 -1 970
box -8 -3 16 105
use FILL  FILL_4481
timestamp 1745462530
transform 1 0 824 0 -1 970
box -8 -3 16 105
use FILL  FILL_4482
timestamp 1745462530
transform 1 0 816 0 -1 970
box -8 -3 16 105
use FILL  FILL_4483
timestamp 1745462530
transform 1 0 776 0 -1 970
box -8 -3 16 105
use FILL  FILL_4484
timestamp 1745462530
transform 1 0 768 0 -1 970
box -8 -3 16 105
use FILL  FILL_4485
timestamp 1745462530
transform 1 0 728 0 -1 970
box -8 -3 16 105
use FILL  FILL_4486
timestamp 1745462530
transform 1 0 720 0 -1 970
box -8 -3 16 105
use FILL  FILL_4487
timestamp 1745462530
transform 1 0 712 0 -1 970
box -8 -3 16 105
use FILL  FILL_4488
timestamp 1745462530
transform 1 0 664 0 -1 970
box -8 -3 16 105
use FILL  FILL_4489
timestamp 1745462530
transform 1 0 656 0 -1 970
box -8 -3 16 105
use FILL  FILL_4490
timestamp 1745462530
transform 1 0 648 0 -1 970
box -8 -3 16 105
use FILL  FILL_4491
timestamp 1745462530
transform 1 0 600 0 -1 970
box -8 -3 16 105
use FILL  FILL_4492
timestamp 1745462530
transform 1 0 592 0 -1 970
box -8 -3 16 105
use FILL  FILL_4493
timestamp 1745462530
transform 1 0 584 0 -1 970
box -8 -3 16 105
use FILL  FILL_4494
timestamp 1745462530
transform 1 0 536 0 -1 970
box -8 -3 16 105
use FILL  FILL_4495
timestamp 1745462530
transform 1 0 504 0 -1 970
box -8 -3 16 105
use FILL  FILL_4496
timestamp 1745462530
transform 1 0 496 0 -1 970
box -8 -3 16 105
use FILL  FILL_4497
timestamp 1745462530
transform 1 0 448 0 -1 970
box -8 -3 16 105
use FILL  FILL_4498
timestamp 1745462530
transform 1 0 440 0 -1 970
box -8 -3 16 105
use FILL  FILL_4499
timestamp 1745462530
transform 1 0 408 0 -1 970
box -8 -3 16 105
use FILL  FILL_4500
timestamp 1745462530
transform 1 0 360 0 -1 970
box -8 -3 16 105
use FILL  FILL_4501
timestamp 1745462530
transform 1 0 352 0 -1 970
box -8 -3 16 105
use FILL  FILL_4502
timestamp 1745462530
transform 1 0 304 0 -1 970
box -8 -3 16 105
use FILL  FILL_4503
timestamp 1745462530
transform 1 0 280 0 -1 970
box -8 -3 16 105
use FILL  FILL_4504
timestamp 1745462530
transform 1 0 272 0 -1 970
box -8 -3 16 105
use FILL  FILL_4505
timestamp 1745462530
transform 1 0 224 0 -1 970
box -8 -3 16 105
use FILL  FILL_4506
timestamp 1745462530
transform 1 0 200 0 -1 970
box -8 -3 16 105
use FILL  FILL_4507
timestamp 1745462530
transform 1 0 192 0 -1 970
box -8 -3 16 105
use FILL  FILL_4508
timestamp 1745462530
transform 1 0 184 0 -1 970
box -8 -3 16 105
use FILL  FILL_4509
timestamp 1745462530
transform 1 0 80 0 -1 970
box -8 -3 16 105
use FILL  FILL_4510
timestamp 1745462530
transform 1 0 72 0 -1 970
box -8 -3 16 105
use FILL  FILL_4511
timestamp 1745462530
transform 1 0 4368 0 1 770
box -8 -3 16 105
use FILL  FILL_4512
timestamp 1745462530
transform 1 0 4264 0 1 770
box -8 -3 16 105
use FILL  FILL_4513
timestamp 1745462530
transform 1 0 4256 0 1 770
box -8 -3 16 105
use FILL  FILL_4514
timestamp 1745462530
transform 1 0 4208 0 1 770
box -8 -3 16 105
use FILL  FILL_4515
timestamp 1745462530
transform 1 0 4184 0 1 770
box -8 -3 16 105
use FILL  FILL_4516
timestamp 1745462530
transform 1 0 4176 0 1 770
box -8 -3 16 105
use FILL  FILL_4517
timestamp 1745462530
transform 1 0 4128 0 1 770
box -8 -3 16 105
use FILL  FILL_4518
timestamp 1745462530
transform 1 0 4120 0 1 770
box -8 -3 16 105
use FILL  FILL_4519
timestamp 1745462530
transform 1 0 4096 0 1 770
box -8 -3 16 105
use FILL  FILL_4520
timestamp 1745462530
transform 1 0 4088 0 1 770
box -8 -3 16 105
use FILL  FILL_4521
timestamp 1745462530
transform 1 0 4040 0 1 770
box -8 -3 16 105
use FILL  FILL_4522
timestamp 1745462530
transform 1 0 4032 0 1 770
box -8 -3 16 105
use FILL  FILL_4523
timestamp 1745462530
transform 1 0 4024 0 1 770
box -8 -3 16 105
use FILL  FILL_4524
timestamp 1745462530
transform 1 0 4000 0 1 770
box -8 -3 16 105
use FILL  FILL_4525
timestamp 1745462530
transform 1 0 3992 0 1 770
box -8 -3 16 105
use FILL  FILL_4526
timestamp 1745462530
transform 1 0 3984 0 1 770
box -8 -3 16 105
use FILL  FILL_4527
timestamp 1745462530
transform 1 0 3936 0 1 770
box -8 -3 16 105
use FILL  FILL_4528
timestamp 1745462530
transform 1 0 3928 0 1 770
box -8 -3 16 105
use FILL  FILL_4529
timestamp 1745462530
transform 1 0 3904 0 1 770
box -8 -3 16 105
use FILL  FILL_4530
timestamp 1745462530
transform 1 0 3896 0 1 770
box -8 -3 16 105
use FILL  FILL_4531
timestamp 1745462530
transform 1 0 3848 0 1 770
box -8 -3 16 105
use FILL  FILL_4532
timestamp 1745462530
transform 1 0 3840 0 1 770
box -8 -3 16 105
use FILL  FILL_4533
timestamp 1745462530
transform 1 0 3792 0 1 770
box -8 -3 16 105
use FILL  FILL_4534
timestamp 1745462530
transform 1 0 3784 0 1 770
box -8 -3 16 105
use FILL  FILL_4535
timestamp 1745462530
transform 1 0 3776 0 1 770
box -8 -3 16 105
use FILL  FILL_4536
timestamp 1745462530
transform 1 0 3736 0 1 770
box -8 -3 16 105
use FILL  FILL_4537
timestamp 1745462530
transform 1 0 3728 0 1 770
box -8 -3 16 105
use FILL  FILL_4538
timestamp 1745462530
transform 1 0 3680 0 1 770
box -8 -3 16 105
use FILL  FILL_4539
timestamp 1745462530
transform 1 0 3672 0 1 770
box -8 -3 16 105
use FILL  FILL_4540
timestamp 1745462530
transform 1 0 3664 0 1 770
box -8 -3 16 105
use FILL  FILL_4541
timestamp 1745462530
transform 1 0 3616 0 1 770
box -8 -3 16 105
use FILL  FILL_4542
timestamp 1745462530
transform 1 0 3608 0 1 770
box -8 -3 16 105
use FILL  FILL_4543
timestamp 1745462530
transform 1 0 3568 0 1 770
box -8 -3 16 105
use FILL  FILL_4544
timestamp 1745462530
transform 1 0 3536 0 1 770
box -8 -3 16 105
use FILL  FILL_4545
timestamp 1745462530
transform 1 0 3528 0 1 770
box -8 -3 16 105
use FILL  FILL_4546
timestamp 1745462530
transform 1 0 3520 0 1 770
box -8 -3 16 105
use FILL  FILL_4547
timestamp 1745462530
transform 1 0 3472 0 1 770
box -8 -3 16 105
use FILL  FILL_4548
timestamp 1745462530
transform 1 0 3464 0 1 770
box -8 -3 16 105
use FILL  FILL_4549
timestamp 1745462530
transform 1 0 3424 0 1 770
box -8 -3 16 105
use FILL  FILL_4550
timestamp 1745462530
transform 1 0 3416 0 1 770
box -8 -3 16 105
use FILL  FILL_4551
timestamp 1745462530
transform 1 0 3408 0 1 770
box -8 -3 16 105
use FILL  FILL_4552
timestamp 1745462530
transform 1 0 3368 0 1 770
box -8 -3 16 105
use FILL  FILL_4553
timestamp 1745462530
transform 1 0 3360 0 1 770
box -8 -3 16 105
use FILL  FILL_4554
timestamp 1745462530
transform 1 0 3312 0 1 770
box -8 -3 16 105
use FILL  FILL_4555
timestamp 1745462530
transform 1 0 3304 0 1 770
box -8 -3 16 105
use FILL  FILL_4556
timestamp 1745462530
transform 1 0 3264 0 1 770
box -8 -3 16 105
use FILL  FILL_4557
timestamp 1745462530
transform 1 0 3232 0 1 770
box -8 -3 16 105
use FILL  FILL_4558
timestamp 1745462530
transform 1 0 3224 0 1 770
box -8 -3 16 105
use FILL  FILL_4559
timestamp 1745462530
transform 1 0 3176 0 1 770
box -8 -3 16 105
use FILL  FILL_4560
timestamp 1745462530
transform 1 0 3168 0 1 770
box -8 -3 16 105
use FILL  FILL_4561
timestamp 1745462530
transform 1 0 3136 0 1 770
box -8 -3 16 105
use FILL  FILL_4562
timestamp 1745462530
transform 1 0 3088 0 1 770
box -8 -3 16 105
use FILL  FILL_4563
timestamp 1745462530
transform 1 0 3080 0 1 770
box -8 -3 16 105
use FILL  FILL_4564
timestamp 1745462530
transform 1 0 3032 0 1 770
box -8 -3 16 105
use FILL  FILL_4565
timestamp 1745462530
transform 1 0 2992 0 1 770
box -8 -3 16 105
use FILL  FILL_4566
timestamp 1745462530
transform 1 0 2872 0 1 770
box -8 -3 16 105
use FILL  FILL_4567
timestamp 1745462530
transform 1 0 2864 0 1 770
box -8 -3 16 105
use FILL  FILL_4568
timestamp 1745462530
transform 1 0 2816 0 1 770
box -8 -3 16 105
use FILL  FILL_4569
timestamp 1745462530
transform 1 0 2808 0 1 770
box -8 -3 16 105
use FILL  FILL_4570
timestamp 1745462530
transform 1 0 2768 0 1 770
box -8 -3 16 105
use FILL  FILL_4571
timestamp 1745462530
transform 1 0 2664 0 1 770
box -8 -3 16 105
use FILL  FILL_4572
timestamp 1745462530
transform 1 0 2616 0 1 770
box -8 -3 16 105
use FILL  FILL_4573
timestamp 1745462530
transform 1 0 2544 0 1 770
box -8 -3 16 105
use FILL  FILL_4574
timestamp 1745462530
transform 1 0 2536 0 1 770
box -8 -3 16 105
use FILL  FILL_4575
timestamp 1745462530
transform 1 0 2488 0 1 770
box -8 -3 16 105
use FILL  FILL_4576
timestamp 1745462530
transform 1 0 2480 0 1 770
box -8 -3 16 105
use FILL  FILL_4577
timestamp 1745462530
transform 1 0 2440 0 1 770
box -8 -3 16 105
use FILL  FILL_4578
timestamp 1745462530
transform 1 0 2432 0 1 770
box -8 -3 16 105
use FILL  FILL_4579
timestamp 1745462530
transform 1 0 2424 0 1 770
box -8 -3 16 105
use FILL  FILL_4580
timestamp 1745462530
transform 1 0 2376 0 1 770
box -8 -3 16 105
use FILL  FILL_4581
timestamp 1745462530
transform 1 0 2368 0 1 770
box -8 -3 16 105
use FILL  FILL_4582
timestamp 1745462530
transform 1 0 2360 0 1 770
box -8 -3 16 105
use FILL  FILL_4583
timestamp 1745462530
transform 1 0 2312 0 1 770
box -8 -3 16 105
use FILL  FILL_4584
timestamp 1745462530
transform 1 0 2288 0 1 770
box -8 -3 16 105
use FILL  FILL_4585
timestamp 1745462530
transform 1 0 2280 0 1 770
box -8 -3 16 105
use FILL  FILL_4586
timestamp 1745462530
transform 1 0 2240 0 1 770
box -8 -3 16 105
use FILL  FILL_4587
timestamp 1745462530
transform 1 0 2136 0 1 770
box -8 -3 16 105
use FILL  FILL_4588
timestamp 1745462530
transform 1 0 2128 0 1 770
box -8 -3 16 105
use FILL  FILL_4589
timestamp 1745462530
transform 1 0 2080 0 1 770
box -8 -3 16 105
use FILL  FILL_4590
timestamp 1745462530
transform 1 0 2072 0 1 770
box -8 -3 16 105
use FILL  FILL_4591
timestamp 1745462530
transform 1 0 2032 0 1 770
box -8 -3 16 105
use FILL  FILL_4592
timestamp 1745462530
transform 1 0 2024 0 1 770
box -8 -3 16 105
use FILL  FILL_4593
timestamp 1745462530
transform 1 0 1984 0 1 770
box -8 -3 16 105
use FILL  FILL_4594
timestamp 1745462530
transform 1 0 1936 0 1 770
box -8 -3 16 105
use FILL  FILL_4595
timestamp 1745462530
transform 1 0 1928 0 1 770
box -8 -3 16 105
use FILL  FILL_4596
timestamp 1745462530
transform 1 0 1800 0 1 770
box -8 -3 16 105
use FILL  FILL_4597
timestamp 1745462530
transform 1 0 1760 0 1 770
box -8 -3 16 105
use FILL  FILL_4598
timestamp 1745462530
transform 1 0 1656 0 1 770
box -8 -3 16 105
use FILL  FILL_4599
timestamp 1745462530
transform 1 0 1616 0 1 770
box -8 -3 16 105
use FILL  FILL_4600
timestamp 1745462530
transform 1 0 1608 0 1 770
box -8 -3 16 105
use FILL  FILL_4601
timestamp 1745462530
transform 1 0 1504 0 1 770
box -8 -3 16 105
use FILL  FILL_4602
timestamp 1745462530
transform 1 0 1456 0 1 770
box -8 -3 16 105
use FILL  FILL_4603
timestamp 1745462530
transform 1 0 1448 0 1 770
box -8 -3 16 105
use FILL  FILL_4604
timestamp 1745462530
transform 1 0 1440 0 1 770
box -8 -3 16 105
use FILL  FILL_4605
timestamp 1745462530
transform 1 0 1392 0 1 770
box -8 -3 16 105
use FILL  FILL_4606
timestamp 1745462530
transform 1 0 1384 0 1 770
box -8 -3 16 105
use FILL  FILL_4607
timestamp 1745462530
transform 1 0 1376 0 1 770
box -8 -3 16 105
use FILL  FILL_4608
timestamp 1745462530
transform 1 0 1272 0 1 770
box -8 -3 16 105
use FILL  FILL_4609
timestamp 1745462530
transform 1 0 1168 0 1 770
box -8 -3 16 105
use FILL  FILL_4610
timestamp 1745462530
transform 1 0 1160 0 1 770
box -8 -3 16 105
use FILL  FILL_4611
timestamp 1745462530
transform 1 0 1152 0 1 770
box -8 -3 16 105
use FILL  FILL_4612
timestamp 1745462530
transform 1 0 1104 0 1 770
box -8 -3 16 105
use FILL  FILL_4613
timestamp 1745462530
transform 1 0 1096 0 1 770
box -8 -3 16 105
use FILL  FILL_4614
timestamp 1745462530
transform 1 0 1088 0 1 770
box -8 -3 16 105
use FILL  FILL_4615
timestamp 1745462530
transform 1 0 1048 0 1 770
box -8 -3 16 105
use FILL  FILL_4616
timestamp 1745462530
transform 1 0 1040 0 1 770
box -8 -3 16 105
use FILL  FILL_4617
timestamp 1745462530
transform 1 0 992 0 1 770
box -8 -3 16 105
use FILL  FILL_4618
timestamp 1745462530
transform 1 0 984 0 1 770
box -8 -3 16 105
use FILL  FILL_4619
timestamp 1745462530
transform 1 0 976 0 1 770
box -8 -3 16 105
use FILL  FILL_4620
timestamp 1745462530
transform 1 0 952 0 1 770
box -8 -3 16 105
use FILL  FILL_4621
timestamp 1745462530
transform 1 0 904 0 1 770
box -8 -3 16 105
use FILL  FILL_4622
timestamp 1745462530
transform 1 0 896 0 1 770
box -8 -3 16 105
use FILL  FILL_4623
timestamp 1745462530
transform 1 0 888 0 1 770
box -8 -3 16 105
use FILL  FILL_4624
timestamp 1745462530
transform 1 0 880 0 1 770
box -8 -3 16 105
use FILL  FILL_4625
timestamp 1745462530
transform 1 0 840 0 1 770
box -8 -3 16 105
use FILL  FILL_4626
timestamp 1745462530
transform 1 0 832 0 1 770
box -8 -3 16 105
use FILL  FILL_4627
timestamp 1745462530
transform 1 0 824 0 1 770
box -8 -3 16 105
use FILL  FILL_4628
timestamp 1745462530
transform 1 0 776 0 1 770
box -8 -3 16 105
use FILL  FILL_4629
timestamp 1745462530
transform 1 0 768 0 1 770
box -8 -3 16 105
use FILL  FILL_4630
timestamp 1745462530
transform 1 0 760 0 1 770
box -8 -3 16 105
use FILL  FILL_4631
timestamp 1745462530
transform 1 0 720 0 1 770
box -8 -3 16 105
use FILL  FILL_4632
timestamp 1745462530
transform 1 0 712 0 1 770
box -8 -3 16 105
use FILL  FILL_4633
timestamp 1745462530
transform 1 0 672 0 1 770
box -8 -3 16 105
use FILL  FILL_4634
timestamp 1745462530
transform 1 0 664 0 1 770
box -8 -3 16 105
use FILL  FILL_4635
timestamp 1745462530
transform 1 0 656 0 1 770
box -8 -3 16 105
use FILL  FILL_4636
timestamp 1745462530
transform 1 0 616 0 1 770
box -8 -3 16 105
use FILL  FILL_4637
timestamp 1745462530
transform 1 0 608 0 1 770
box -8 -3 16 105
use FILL  FILL_4638
timestamp 1745462530
transform 1 0 560 0 1 770
box -8 -3 16 105
use FILL  FILL_4639
timestamp 1745462530
transform 1 0 552 0 1 770
box -8 -3 16 105
use FILL  FILL_4640
timestamp 1745462530
transform 1 0 544 0 1 770
box -8 -3 16 105
use FILL  FILL_4641
timestamp 1745462530
transform 1 0 472 0 1 770
box -8 -3 16 105
use FILL  FILL_4642
timestamp 1745462530
transform 1 0 464 0 1 770
box -8 -3 16 105
use FILL  FILL_4643
timestamp 1745462530
transform 1 0 408 0 1 770
box -8 -3 16 105
use FILL  FILL_4644
timestamp 1745462530
transform 1 0 400 0 1 770
box -8 -3 16 105
use FILL  FILL_4645
timestamp 1745462530
transform 1 0 352 0 1 770
box -8 -3 16 105
use FILL  FILL_4646
timestamp 1745462530
transform 1 0 248 0 1 770
box -8 -3 16 105
use FILL  FILL_4647
timestamp 1745462530
transform 1 0 184 0 1 770
box -8 -3 16 105
use FILL  FILL_4648
timestamp 1745462530
transform 1 0 176 0 1 770
box -8 -3 16 105
use FILL  FILL_4649
timestamp 1745462530
transform 1 0 72 0 1 770
box -8 -3 16 105
use FILL  FILL_4650
timestamp 1745462530
transform 1 0 4368 0 -1 770
box -8 -3 16 105
use FILL  FILL_4651
timestamp 1745462530
transform 1 0 4264 0 -1 770
box -8 -3 16 105
use FILL  FILL_4652
timestamp 1745462530
transform 1 0 4256 0 -1 770
box -8 -3 16 105
use FILL  FILL_4653
timestamp 1745462530
transform 1 0 4232 0 -1 770
box -8 -3 16 105
use FILL  FILL_4654
timestamp 1745462530
transform 1 0 4224 0 -1 770
box -8 -3 16 105
use FILL  FILL_4655
timestamp 1745462530
transform 1 0 4216 0 -1 770
box -8 -3 16 105
use FILL  FILL_4656
timestamp 1745462530
transform 1 0 4112 0 -1 770
box -8 -3 16 105
use FILL  FILL_4657
timestamp 1745462530
transform 1 0 4088 0 -1 770
box -8 -3 16 105
use FILL  FILL_4658
timestamp 1745462530
transform 1 0 4080 0 -1 770
box -8 -3 16 105
use FILL  FILL_4659
timestamp 1745462530
transform 1 0 4072 0 -1 770
box -8 -3 16 105
use FILL  FILL_4660
timestamp 1745462530
transform 1 0 3968 0 -1 770
box -8 -3 16 105
use FILL  FILL_4661
timestamp 1745462530
transform 1 0 3960 0 -1 770
box -8 -3 16 105
use FILL  FILL_4662
timestamp 1745462530
transform 1 0 3952 0 -1 770
box -8 -3 16 105
use FILL  FILL_4663
timestamp 1745462530
transform 1 0 3944 0 -1 770
box -8 -3 16 105
use FILL  FILL_4664
timestamp 1745462530
transform 1 0 3840 0 -1 770
box -8 -3 16 105
use FILL  FILL_4665
timestamp 1745462530
transform 1 0 3832 0 -1 770
box -8 -3 16 105
use FILL  FILL_4666
timestamp 1745462530
transform 1 0 3824 0 -1 770
box -8 -3 16 105
use FILL  FILL_4667
timestamp 1745462530
transform 1 0 3816 0 -1 770
box -8 -3 16 105
use FILL  FILL_4668
timestamp 1745462530
transform 1 0 3792 0 -1 770
box -8 -3 16 105
use FILL  FILL_4669
timestamp 1745462530
transform 1 0 3784 0 -1 770
box -8 -3 16 105
use FILL  FILL_4670
timestamp 1745462530
transform 1 0 3776 0 -1 770
box -8 -3 16 105
use FILL  FILL_4671
timestamp 1745462530
transform 1 0 3736 0 -1 770
box -8 -3 16 105
use FILL  FILL_4672
timestamp 1745462530
transform 1 0 3728 0 -1 770
box -8 -3 16 105
use FILL  FILL_4673
timestamp 1745462530
transform 1 0 3720 0 -1 770
box -8 -3 16 105
use FILL  FILL_4674
timestamp 1745462530
transform 1 0 3712 0 -1 770
box -8 -3 16 105
use FILL  FILL_4675
timestamp 1745462530
transform 1 0 3664 0 -1 770
box -8 -3 16 105
use FILL  FILL_4676
timestamp 1745462530
transform 1 0 3656 0 -1 770
box -8 -3 16 105
use FILL  FILL_4677
timestamp 1745462530
transform 1 0 3648 0 -1 770
box -8 -3 16 105
use FILL  FILL_4678
timestamp 1745462530
transform 1 0 3640 0 -1 770
box -8 -3 16 105
use FILL  FILL_4679
timestamp 1745462530
transform 1 0 3600 0 -1 770
box -8 -3 16 105
use FILL  FILL_4680
timestamp 1745462530
transform 1 0 3592 0 -1 770
box -8 -3 16 105
use FILL  FILL_4681
timestamp 1745462530
transform 1 0 3584 0 -1 770
box -8 -3 16 105
use FILL  FILL_4682
timestamp 1745462530
transform 1 0 3560 0 -1 770
box -8 -3 16 105
use FILL  FILL_4683
timestamp 1745462530
transform 1 0 3552 0 -1 770
box -8 -3 16 105
use FILL  FILL_4684
timestamp 1745462530
transform 1 0 3448 0 -1 770
box -8 -3 16 105
use FILL  FILL_4685
timestamp 1745462530
transform 1 0 3440 0 -1 770
box -8 -3 16 105
use FILL  FILL_4686
timestamp 1745462530
transform 1 0 3432 0 -1 770
box -8 -3 16 105
use FILL  FILL_4687
timestamp 1745462530
transform 1 0 3328 0 -1 770
box -8 -3 16 105
use FILL  FILL_4688
timestamp 1745462530
transform 1 0 3320 0 -1 770
box -8 -3 16 105
use FILL  FILL_4689
timestamp 1745462530
transform 1 0 3312 0 -1 770
box -8 -3 16 105
use FILL  FILL_4690
timestamp 1745462530
transform 1 0 3272 0 -1 770
box -8 -3 16 105
use FILL  FILL_4691
timestamp 1745462530
transform 1 0 3264 0 -1 770
box -8 -3 16 105
use FILL  FILL_4692
timestamp 1745462530
transform 1 0 3240 0 -1 770
box -8 -3 16 105
use FILL  FILL_4693
timestamp 1745462530
transform 1 0 3232 0 -1 770
box -8 -3 16 105
use FILL  FILL_4694
timestamp 1745462530
transform 1 0 3128 0 -1 770
box -8 -3 16 105
use FILL  FILL_4695
timestamp 1745462530
transform 1 0 3104 0 -1 770
box -8 -3 16 105
use FILL  FILL_4696
timestamp 1745462530
transform 1 0 3056 0 -1 770
box -8 -3 16 105
use FILL  FILL_4697
timestamp 1745462530
transform 1 0 3048 0 -1 770
box -8 -3 16 105
use FILL  FILL_4698
timestamp 1745462530
transform 1 0 3040 0 -1 770
box -8 -3 16 105
use FILL  FILL_4699
timestamp 1745462530
transform 1 0 3000 0 -1 770
box -8 -3 16 105
use FILL  FILL_4700
timestamp 1745462530
transform 1 0 2968 0 -1 770
box -8 -3 16 105
use FILL  FILL_4701
timestamp 1745462530
transform 1 0 2960 0 -1 770
box -8 -3 16 105
use FILL  FILL_4702
timestamp 1745462530
transform 1 0 2912 0 -1 770
box -8 -3 16 105
use FILL  FILL_4703
timestamp 1745462530
transform 1 0 2904 0 -1 770
box -8 -3 16 105
use FILL  FILL_4704
timestamp 1745462530
transform 1 0 2800 0 -1 770
box -8 -3 16 105
use FILL  FILL_4705
timestamp 1745462530
transform 1 0 2776 0 -1 770
box -8 -3 16 105
use FILL  FILL_4706
timestamp 1745462530
transform 1 0 2728 0 -1 770
box -8 -3 16 105
use FILL  FILL_4707
timestamp 1745462530
transform 1 0 2720 0 -1 770
box -8 -3 16 105
use FILL  FILL_4708
timestamp 1745462530
transform 1 0 2696 0 -1 770
box -8 -3 16 105
use FILL  FILL_4709
timestamp 1745462530
transform 1 0 2648 0 -1 770
box -8 -3 16 105
use FILL  FILL_4710
timestamp 1745462530
transform 1 0 2640 0 -1 770
box -8 -3 16 105
use FILL  FILL_4711
timestamp 1745462530
transform 1 0 2632 0 -1 770
box -8 -3 16 105
use FILL  FILL_4712
timestamp 1745462530
transform 1 0 2592 0 -1 770
box -8 -3 16 105
use FILL  FILL_4713
timestamp 1745462530
transform 1 0 2560 0 -1 770
box -8 -3 16 105
use FILL  FILL_4714
timestamp 1745462530
transform 1 0 2552 0 -1 770
box -8 -3 16 105
use FILL  FILL_4715
timestamp 1745462530
transform 1 0 2512 0 -1 770
box -8 -3 16 105
use FILL  FILL_4716
timestamp 1745462530
transform 1 0 2504 0 -1 770
box -8 -3 16 105
use FILL  FILL_4717
timestamp 1745462530
transform 1 0 2496 0 -1 770
box -8 -3 16 105
use FILL  FILL_4718
timestamp 1745462530
transform 1 0 2448 0 -1 770
box -8 -3 16 105
use FILL  FILL_4719
timestamp 1745462530
transform 1 0 2424 0 -1 770
box -8 -3 16 105
use FILL  FILL_4720
timestamp 1745462530
transform 1 0 2320 0 -1 770
box -8 -3 16 105
use FILL  FILL_4721
timestamp 1745462530
transform 1 0 2312 0 -1 770
box -8 -3 16 105
use FILL  FILL_4722
timestamp 1745462530
transform 1 0 2264 0 -1 770
box -8 -3 16 105
use FILL  FILL_4723
timestamp 1745462530
transform 1 0 2256 0 -1 770
box -8 -3 16 105
use FILL  FILL_4724
timestamp 1745462530
transform 1 0 2232 0 -1 770
box -8 -3 16 105
use FILL  FILL_4725
timestamp 1745462530
transform 1 0 2224 0 -1 770
box -8 -3 16 105
use FILL  FILL_4726
timestamp 1745462530
transform 1 0 2176 0 -1 770
box -8 -3 16 105
use FILL  FILL_4727
timestamp 1745462530
transform 1 0 2168 0 -1 770
box -8 -3 16 105
use FILL  FILL_4728
timestamp 1745462530
transform 1 0 2064 0 -1 770
box -8 -3 16 105
use FILL  FILL_4729
timestamp 1745462530
transform 1 0 2056 0 -1 770
box -8 -3 16 105
use FILL  FILL_4730
timestamp 1745462530
transform 1 0 1952 0 -1 770
box -8 -3 16 105
use FILL  FILL_4731
timestamp 1745462530
transform 1 0 1928 0 -1 770
box -8 -3 16 105
use FILL  FILL_4732
timestamp 1745462530
transform 1 0 1920 0 -1 770
box -8 -3 16 105
use FILL  FILL_4733
timestamp 1745462530
transform 1 0 1872 0 -1 770
box -8 -3 16 105
use FILL  FILL_4734
timestamp 1745462530
transform 1 0 1864 0 -1 770
box -8 -3 16 105
use FILL  FILL_4735
timestamp 1745462530
transform 1 0 1856 0 -1 770
box -8 -3 16 105
use FILL  FILL_4736
timestamp 1745462530
transform 1 0 1808 0 -1 770
box -8 -3 16 105
use FILL  FILL_4737
timestamp 1745462530
transform 1 0 1800 0 -1 770
box -8 -3 16 105
use FILL  FILL_4738
timestamp 1745462530
transform 1 0 1776 0 -1 770
box -8 -3 16 105
use FILL  FILL_4739
timestamp 1745462530
transform 1 0 1768 0 -1 770
box -8 -3 16 105
use FILL  FILL_4740
timestamp 1745462530
transform 1 0 1760 0 -1 770
box -8 -3 16 105
use FILL  FILL_4741
timestamp 1745462530
transform 1 0 1712 0 -1 770
box -8 -3 16 105
use FILL  FILL_4742
timestamp 1745462530
transform 1 0 1704 0 -1 770
box -8 -3 16 105
use FILL  FILL_4743
timestamp 1745462530
transform 1 0 1680 0 -1 770
box -8 -3 16 105
use FILL  FILL_4744
timestamp 1745462530
transform 1 0 1672 0 -1 770
box -8 -3 16 105
use FILL  FILL_4745
timestamp 1745462530
transform 1 0 1640 0 -1 770
box -8 -3 16 105
use FILL  FILL_4746
timestamp 1745462530
transform 1 0 1632 0 -1 770
box -8 -3 16 105
use FILL  FILL_4747
timestamp 1745462530
transform 1 0 1608 0 -1 770
box -8 -3 16 105
use FILL  FILL_4748
timestamp 1745462530
transform 1 0 1600 0 -1 770
box -8 -3 16 105
use FILL  FILL_4749
timestamp 1745462530
transform 1 0 1568 0 -1 770
box -8 -3 16 105
use FILL  FILL_4750
timestamp 1745462530
transform 1 0 1544 0 -1 770
box -8 -3 16 105
use FILL  FILL_4751
timestamp 1745462530
transform 1 0 1536 0 -1 770
box -8 -3 16 105
use FILL  FILL_4752
timestamp 1745462530
transform 1 0 1528 0 -1 770
box -8 -3 16 105
use FILL  FILL_4753
timestamp 1745462530
transform 1 0 1488 0 -1 770
box -8 -3 16 105
use FILL  FILL_4754
timestamp 1745462530
transform 1 0 1480 0 -1 770
box -8 -3 16 105
use FILL  FILL_4755
timestamp 1745462530
transform 1 0 1456 0 -1 770
box -8 -3 16 105
use FILL  FILL_4756
timestamp 1745462530
transform 1 0 1448 0 -1 770
box -8 -3 16 105
use FILL  FILL_4757
timestamp 1745462530
transform 1 0 1400 0 -1 770
box -8 -3 16 105
use FILL  FILL_4758
timestamp 1745462530
transform 1 0 1392 0 -1 770
box -8 -3 16 105
use FILL  FILL_4759
timestamp 1745462530
transform 1 0 1384 0 -1 770
box -8 -3 16 105
use FILL  FILL_4760
timestamp 1745462530
transform 1 0 1376 0 -1 770
box -8 -3 16 105
use FILL  FILL_4761
timestamp 1745462530
transform 1 0 1328 0 -1 770
box -8 -3 16 105
use FILL  FILL_4762
timestamp 1745462530
transform 1 0 1320 0 -1 770
box -8 -3 16 105
use FILL  FILL_4763
timestamp 1745462530
transform 1 0 1296 0 -1 770
box -8 -3 16 105
use FILL  FILL_4764
timestamp 1745462530
transform 1 0 1288 0 -1 770
box -8 -3 16 105
use FILL  FILL_4765
timestamp 1745462530
transform 1 0 1240 0 -1 770
box -8 -3 16 105
use FILL  FILL_4766
timestamp 1745462530
transform 1 0 1232 0 -1 770
box -8 -3 16 105
use FILL  FILL_4767
timestamp 1745462530
transform 1 0 1224 0 -1 770
box -8 -3 16 105
use FILL  FILL_4768
timestamp 1745462530
transform 1 0 1200 0 -1 770
box -8 -3 16 105
use FILL  FILL_4769
timestamp 1745462530
transform 1 0 1096 0 -1 770
box -8 -3 16 105
use FILL  FILL_4770
timestamp 1745462530
transform 1 0 1088 0 -1 770
box -8 -3 16 105
use FILL  FILL_4771
timestamp 1745462530
transform 1 0 1080 0 -1 770
box -8 -3 16 105
use FILL  FILL_4772
timestamp 1745462530
transform 1 0 1032 0 -1 770
box -8 -3 16 105
use FILL  FILL_4773
timestamp 1745462530
transform 1 0 1024 0 -1 770
box -8 -3 16 105
use FILL  FILL_4774
timestamp 1745462530
transform 1 0 1016 0 -1 770
box -8 -3 16 105
use FILL  FILL_4775
timestamp 1745462530
transform 1 0 968 0 -1 770
box -8 -3 16 105
use FILL  FILL_4776
timestamp 1745462530
transform 1 0 960 0 -1 770
box -8 -3 16 105
use FILL  FILL_4777
timestamp 1745462530
transform 1 0 952 0 -1 770
box -8 -3 16 105
use FILL  FILL_4778
timestamp 1745462530
transform 1 0 920 0 -1 770
box -8 -3 16 105
use FILL  FILL_4779
timestamp 1745462530
transform 1 0 912 0 -1 770
box -8 -3 16 105
use FILL  FILL_4780
timestamp 1745462530
transform 1 0 880 0 -1 770
box -8 -3 16 105
use FILL  FILL_4781
timestamp 1745462530
transform 1 0 872 0 -1 770
box -8 -3 16 105
use FILL  FILL_4782
timestamp 1745462530
transform 1 0 840 0 -1 770
box -8 -3 16 105
use FILL  FILL_4783
timestamp 1745462530
transform 1 0 832 0 -1 770
box -8 -3 16 105
use FILL  FILL_4784
timestamp 1745462530
transform 1 0 792 0 -1 770
box -8 -3 16 105
use FILL  FILL_4785
timestamp 1745462530
transform 1 0 784 0 -1 770
box -8 -3 16 105
use FILL  FILL_4786
timestamp 1745462530
transform 1 0 776 0 -1 770
box -8 -3 16 105
use FILL  FILL_4787
timestamp 1745462530
transform 1 0 728 0 -1 770
box -8 -3 16 105
use FILL  FILL_4788
timestamp 1745462530
transform 1 0 720 0 -1 770
box -8 -3 16 105
use FILL  FILL_4789
timestamp 1745462530
transform 1 0 712 0 -1 770
box -8 -3 16 105
use FILL  FILL_4790
timestamp 1745462530
transform 1 0 664 0 -1 770
box -8 -3 16 105
use FILL  FILL_4791
timestamp 1745462530
transform 1 0 656 0 -1 770
box -8 -3 16 105
use FILL  FILL_4792
timestamp 1745462530
transform 1 0 648 0 -1 770
box -8 -3 16 105
use FILL  FILL_4793
timestamp 1745462530
transform 1 0 608 0 -1 770
box -8 -3 16 105
use FILL  FILL_4794
timestamp 1745462530
transform 1 0 600 0 -1 770
box -8 -3 16 105
use FILL  FILL_4795
timestamp 1745462530
transform 1 0 560 0 -1 770
box -8 -3 16 105
use FILL  FILL_4796
timestamp 1745462530
transform 1 0 552 0 -1 770
box -8 -3 16 105
use FILL  FILL_4797
timestamp 1745462530
transform 1 0 544 0 -1 770
box -8 -3 16 105
use FILL  FILL_4798
timestamp 1745462530
transform 1 0 496 0 -1 770
box -8 -3 16 105
use FILL  FILL_4799
timestamp 1745462530
transform 1 0 488 0 -1 770
box -8 -3 16 105
use FILL  FILL_4800
timestamp 1745462530
transform 1 0 480 0 -1 770
box -8 -3 16 105
use FILL  FILL_4801
timestamp 1745462530
transform 1 0 448 0 -1 770
box -8 -3 16 105
use FILL  FILL_4802
timestamp 1745462530
transform 1 0 440 0 -1 770
box -8 -3 16 105
use FILL  FILL_4803
timestamp 1745462530
transform 1 0 392 0 -1 770
box -8 -3 16 105
use FILL  FILL_4804
timestamp 1745462530
transform 1 0 384 0 -1 770
box -8 -3 16 105
use FILL  FILL_4805
timestamp 1745462530
transform 1 0 376 0 -1 770
box -8 -3 16 105
use FILL  FILL_4806
timestamp 1745462530
transform 1 0 344 0 -1 770
box -8 -3 16 105
use FILL  FILL_4807
timestamp 1745462530
transform 1 0 336 0 -1 770
box -8 -3 16 105
use FILL  FILL_4808
timestamp 1745462530
transform 1 0 288 0 -1 770
box -8 -3 16 105
use FILL  FILL_4809
timestamp 1745462530
transform 1 0 280 0 -1 770
box -8 -3 16 105
use FILL  FILL_4810
timestamp 1745462530
transform 1 0 272 0 -1 770
box -8 -3 16 105
use FILL  FILL_4811
timestamp 1745462530
transform 1 0 248 0 -1 770
box -8 -3 16 105
use FILL  FILL_4812
timestamp 1745462530
transform 1 0 240 0 -1 770
box -8 -3 16 105
use FILL  FILL_4813
timestamp 1745462530
transform 1 0 232 0 -1 770
box -8 -3 16 105
use FILL  FILL_4814
timestamp 1745462530
transform 1 0 128 0 -1 770
box -8 -3 16 105
use FILL  FILL_4815
timestamp 1745462530
transform 1 0 120 0 -1 770
box -8 -3 16 105
use FILL  FILL_4816
timestamp 1745462530
transform 1 0 112 0 -1 770
box -8 -3 16 105
use FILL  FILL_4817
timestamp 1745462530
transform 1 0 104 0 -1 770
box -8 -3 16 105
use FILL  FILL_4818
timestamp 1745462530
transform 1 0 96 0 -1 770
box -8 -3 16 105
use FILL  FILL_4819
timestamp 1745462530
transform 1 0 88 0 -1 770
box -8 -3 16 105
use FILL  FILL_4820
timestamp 1745462530
transform 1 0 80 0 -1 770
box -8 -3 16 105
use FILL  FILL_4821
timestamp 1745462530
transform 1 0 72 0 -1 770
box -8 -3 16 105
use FILL  FILL_4822
timestamp 1745462530
transform 1 0 4368 0 1 570
box -8 -3 16 105
use FILL  FILL_4823
timestamp 1745462530
transform 1 0 4360 0 1 570
box -8 -3 16 105
use FILL  FILL_4824
timestamp 1745462530
transform 1 0 4352 0 1 570
box -8 -3 16 105
use FILL  FILL_4825
timestamp 1745462530
transform 1 0 4304 0 1 570
box -8 -3 16 105
use FILL  FILL_4826
timestamp 1745462530
transform 1 0 4296 0 1 570
box -8 -3 16 105
use FILL  FILL_4827
timestamp 1745462530
transform 1 0 4288 0 1 570
box -8 -3 16 105
use FILL  FILL_4828
timestamp 1745462530
transform 1 0 4184 0 1 570
box -8 -3 16 105
use FILL  FILL_4829
timestamp 1745462530
transform 1 0 4176 0 1 570
box -8 -3 16 105
use FILL  FILL_4830
timestamp 1745462530
transform 1 0 4128 0 1 570
box -8 -3 16 105
use FILL  FILL_4831
timestamp 1745462530
transform 1 0 4120 0 1 570
box -8 -3 16 105
use FILL  FILL_4832
timestamp 1745462530
transform 1 0 4072 0 1 570
box -8 -3 16 105
use FILL  FILL_4833
timestamp 1745462530
transform 1 0 4048 0 1 570
box -8 -3 16 105
use FILL  FILL_4834
timestamp 1745462530
transform 1 0 4040 0 1 570
box -8 -3 16 105
use FILL  FILL_4835
timestamp 1745462530
transform 1 0 3936 0 1 570
box -8 -3 16 105
use FILL  FILL_4836
timestamp 1745462530
transform 1 0 3928 0 1 570
box -8 -3 16 105
use FILL  FILL_4837
timestamp 1745462530
transform 1 0 3824 0 1 570
box -8 -3 16 105
use FILL  FILL_4838
timestamp 1745462530
transform 1 0 3816 0 1 570
box -8 -3 16 105
use FILL  FILL_4839
timestamp 1745462530
transform 1 0 3808 0 1 570
box -8 -3 16 105
use FILL  FILL_4840
timestamp 1745462530
transform 1 0 3760 0 1 570
box -8 -3 16 105
use FILL  FILL_4841
timestamp 1745462530
transform 1 0 3752 0 1 570
box -8 -3 16 105
use FILL  FILL_4842
timestamp 1745462530
transform 1 0 3744 0 1 570
box -8 -3 16 105
use FILL  FILL_4843
timestamp 1745462530
transform 1 0 3696 0 1 570
box -8 -3 16 105
use FILL  FILL_4844
timestamp 1745462530
transform 1 0 3664 0 1 570
box -8 -3 16 105
use FILL  FILL_4845
timestamp 1745462530
transform 1 0 3656 0 1 570
box -8 -3 16 105
use FILL  FILL_4846
timestamp 1745462530
transform 1 0 3608 0 1 570
box -8 -3 16 105
use FILL  FILL_4847
timestamp 1745462530
transform 1 0 3600 0 1 570
box -8 -3 16 105
use FILL  FILL_4848
timestamp 1745462530
transform 1 0 3552 0 1 570
box -8 -3 16 105
use FILL  FILL_4849
timestamp 1745462530
transform 1 0 3544 0 1 570
box -8 -3 16 105
use FILL  FILL_4850
timestamp 1745462530
transform 1 0 3496 0 1 570
box -8 -3 16 105
use FILL  FILL_4851
timestamp 1745462530
transform 1 0 3488 0 1 570
box -8 -3 16 105
use FILL  FILL_4852
timestamp 1745462530
transform 1 0 3456 0 1 570
box -8 -3 16 105
use FILL  FILL_4853
timestamp 1745462530
transform 1 0 3408 0 1 570
box -8 -3 16 105
use FILL  FILL_4854
timestamp 1745462530
transform 1 0 3400 0 1 570
box -8 -3 16 105
use FILL  FILL_4855
timestamp 1745462530
transform 1 0 3352 0 1 570
box -8 -3 16 105
use FILL  FILL_4856
timestamp 1745462530
transform 1 0 3328 0 1 570
box -8 -3 16 105
use FILL  FILL_4857
timestamp 1745462530
transform 1 0 3296 0 1 570
box -8 -3 16 105
use FILL  FILL_4858
timestamp 1745462530
transform 1 0 3264 0 1 570
box -8 -3 16 105
use FILL  FILL_4859
timestamp 1745462530
transform 1 0 3256 0 1 570
box -8 -3 16 105
use FILL  FILL_4860
timestamp 1745462530
transform 1 0 3224 0 1 570
box -8 -3 16 105
use FILL  FILL_4861
timestamp 1745462530
transform 1 0 3192 0 1 570
box -8 -3 16 105
use FILL  FILL_4862
timestamp 1745462530
transform 1 0 3184 0 1 570
box -8 -3 16 105
use FILL  FILL_4863
timestamp 1745462530
transform 1 0 3080 0 1 570
box -8 -3 16 105
use FILL  FILL_4864
timestamp 1745462530
transform 1 0 3056 0 1 570
box -8 -3 16 105
use FILL  FILL_4865
timestamp 1745462530
transform 1 0 3008 0 1 570
box -8 -3 16 105
use FILL  FILL_4866
timestamp 1745462530
transform 1 0 3000 0 1 570
box -8 -3 16 105
use FILL  FILL_4867
timestamp 1745462530
transform 1 0 2992 0 1 570
box -8 -3 16 105
use FILL  FILL_4868
timestamp 1745462530
transform 1 0 2944 0 1 570
box -8 -3 16 105
use FILL  FILL_4869
timestamp 1745462530
transform 1 0 2912 0 1 570
box -8 -3 16 105
use FILL  FILL_4870
timestamp 1745462530
transform 1 0 2904 0 1 570
box -8 -3 16 105
use FILL  FILL_4871
timestamp 1745462530
transform 1 0 2856 0 1 570
box -8 -3 16 105
use FILL  FILL_4872
timestamp 1745462530
transform 1 0 2848 0 1 570
box -8 -3 16 105
use FILL  FILL_4873
timestamp 1745462530
transform 1 0 2840 0 1 570
box -8 -3 16 105
use FILL  FILL_4874
timestamp 1745462530
transform 1 0 2808 0 1 570
box -8 -3 16 105
use FILL  FILL_4875
timestamp 1745462530
transform 1 0 2800 0 1 570
box -8 -3 16 105
use FILL  FILL_4876
timestamp 1745462530
transform 1 0 2752 0 1 570
box -8 -3 16 105
use FILL  FILL_4877
timestamp 1745462530
transform 1 0 2744 0 1 570
box -8 -3 16 105
use FILL  FILL_4878
timestamp 1745462530
transform 1 0 2736 0 1 570
box -8 -3 16 105
use FILL  FILL_4879
timestamp 1745462530
transform 1 0 2688 0 1 570
box -8 -3 16 105
use FILL  FILL_4880
timestamp 1745462530
transform 1 0 2680 0 1 570
box -8 -3 16 105
use FILL  FILL_4881
timestamp 1745462530
transform 1 0 2648 0 1 570
box -8 -3 16 105
use FILL  FILL_4882
timestamp 1745462530
transform 1 0 2640 0 1 570
box -8 -3 16 105
use FILL  FILL_4883
timestamp 1745462530
transform 1 0 2608 0 1 570
box -8 -3 16 105
use FILL  FILL_4884
timestamp 1745462530
transform 1 0 2600 0 1 570
box -8 -3 16 105
use FILL  FILL_4885
timestamp 1745462530
transform 1 0 2568 0 1 570
box -8 -3 16 105
use FILL  FILL_4886
timestamp 1745462530
transform 1 0 2560 0 1 570
box -8 -3 16 105
use FILL  FILL_4887
timestamp 1745462530
transform 1 0 2552 0 1 570
box -8 -3 16 105
use FILL  FILL_4888
timestamp 1745462530
transform 1 0 2504 0 1 570
box -8 -3 16 105
use FILL  FILL_4889
timestamp 1745462530
transform 1 0 2496 0 1 570
box -8 -3 16 105
use FILL  FILL_4890
timestamp 1745462530
transform 1 0 2488 0 1 570
box -8 -3 16 105
use FILL  FILL_4891
timestamp 1745462530
transform 1 0 2456 0 1 570
box -8 -3 16 105
use FILL  FILL_4892
timestamp 1745462530
transform 1 0 2424 0 1 570
box -8 -3 16 105
use FILL  FILL_4893
timestamp 1745462530
transform 1 0 2416 0 1 570
box -8 -3 16 105
use FILL  FILL_4894
timestamp 1745462530
transform 1 0 2408 0 1 570
box -8 -3 16 105
use FILL  FILL_4895
timestamp 1745462530
transform 1 0 2360 0 1 570
box -8 -3 16 105
use FILL  FILL_4896
timestamp 1745462530
transform 1 0 2352 0 1 570
box -8 -3 16 105
use FILL  FILL_4897
timestamp 1745462530
transform 1 0 2304 0 1 570
box -8 -3 16 105
use FILL  FILL_4898
timestamp 1745462530
transform 1 0 2296 0 1 570
box -8 -3 16 105
use FILL  FILL_4899
timestamp 1745462530
transform 1 0 2288 0 1 570
box -8 -3 16 105
use FILL  FILL_4900
timestamp 1745462530
transform 1 0 2240 0 1 570
box -8 -3 16 105
use FILL  FILL_4901
timestamp 1745462530
transform 1 0 2232 0 1 570
box -8 -3 16 105
use FILL  FILL_4902
timestamp 1745462530
transform 1 0 2224 0 1 570
box -8 -3 16 105
use FILL  FILL_4903
timestamp 1745462530
transform 1 0 2176 0 1 570
box -8 -3 16 105
use FILL  FILL_4904
timestamp 1745462530
transform 1 0 2152 0 1 570
box -8 -3 16 105
use FILL  FILL_4905
timestamp 1745462530
transform 1 0 2048 0 1 570
box -8 -3 16 105
use FILL  FILL_4906
timestamp 1745462530
transform 1 0 2040 0 1 570
box -8 -3 16 105
use FILL  FILL_4907
timestamp 1745462530
transform 1 0 1992 0 1 570
box -8 -3 16 105
use FILL  FILL_4908
timestamp 1745462530
transform 1 0 1984 0 1 570
box -8 -3 16 105
use FILL  FILL_4909
timestamp 1745462530
transform 1 0 1976 0 1 570
box -8 -3 16 105
use FILL  FILL_4910
timestamp 1745462530
transform 1 0 1928 0 1 570
box -8 -3 16 105
use FILL  FILL_4911
timestamp 1745462530
transform 1 0 1920 0 1 570
box -8 -3 16 105
use FILL  FILL_4912
timestamp 1745462530
transform 1 0 1880 0 1 570
box -8 -3 16 105
use FILL  FILL_4913
timestamp 1745462530
transform 1 0 1848 0 1 570
box -8 -3 16 105
use FILL  FILL_4914
timestamp 1745462530
transform 1 0 1840 0 1 570
box -8 -3 16 105
use FILL  FILL_4915
timestamp 1745462530
transform 1 0 1832 0 1 570
box -8 -3 16 105
use FILL  FILL_4916
timestamp 1745462530
transform 1 0 1784 0 1 570
box -8 -3 16 105
use FILL  FILL_4917
timestamp 1745462530
transform 1 0 1776 0 1 570
box -8 -3 16 105
use FILL  FILL_4918
timestamp 1745462530
transform 1 0 1728 0 1 570
box -8 -3 16 105
use FILL  FILL_4919
timestamp 1745462530
transform 1 0 1720 0 1 570
box -8 -3 16 105
use FILL  FILL_4920
timestamp 1745462530
transform 1 0 1672 0 1 570
box -8 -3 16 105
use FILL  FILL_4921
timestamp 1745462530
transform 1 0 1664 0 1 570
box -8 -3 16 105
use FILL  FILL_4922
timestamp 1745462530
transform 1 0 1656 0 1 570
box -8 -3 16 105
use FILL  FILL_4923
timestamp 1745462530
transform 1 0 1608 0 1 570
box -8 -3 16 105
use FILL  FILL_4924
timestamp 1745462530
transform 1 0 1600 0 1 570
box -8 -3 16 105
use FILL  FILL_4925
timestamp 1745462530
transform 1 0 1568 0 1 570
box -8 -3 16 105
use FILL  FILL_4926
timestamp 1745462530
transform 1 0 1536 0 1 570
box -8 -3 16 105
use FILL  FILL_4927
timestamp 1745462530
transform 1 0 1504 0 1 570
box -8 -3 16 105
use FILL  FILL_4928
timestamp 1745462530
transform 1 0 1496 0 1 570
box -8 -3 16 105
use FILL  FILL_4929
timestamp 1745462530
transform 1 0 1464 0 1 570
box -8 -3 16 105
use FILL  FILL_4930
timestamp 1745462530
transform 1 0 1456 0 1 570
box -8 -3 16 105
use FILL  FILL_4931
timestamp 1745462530
transform 1 0 1408 0 1 570
box -8 -3 16 105
use FILL  FILL_4932
timestamp 1745462530
transform 1 0 1400 0 1 570
box -8 -3 16 105
use FILL  FILL_4933
timestamp 1745462530
transform 1 0 1352 0 1 570
box -8 -3 16 105
use FILL  FILL_4934
timestamp 1745462530
transform 1 0 1344 0 1 570
box -8 -3 16 105
use FILL  FILL_4935
timestamp 1745462530
transform 1 0 1296 0 1 570
box -8 -3 16 105
use FILL  FILL_4936
timestamp 1745462530
transform 1 0 1288 0 1 570
box -8 -3 16 105
use FILL  FILL_4937
timestamp 1745462530
transform 1 0 1280 0 1 570
box -8 -3 16 105
use FILL  FILL_4938
timestamp 1745462530
transform 1 0 1232 0 1 570
box -8 -3 16 105
use FILL  FILL_4939
timestamp 1745462530
transform 1 0 1224 0 1 570
box -8 -3 16 105
use FILL  FILL_4940
timestamp 1745462530
transform 1 0 1192 0 1 570
box -8 -3 16 105
use FILL  FILL_4941
timestamp 1745462530
transform 1 0 1160 0 1 570
box -8 -3 16 105
use FILL  FILL_4942
timestamp 1745462530
transform 1 0 1152 0 1 570
box -8 -3 16 105
use FILL  FILL_4943
timestamp 1745462530
transform 1 0 1104 0 1 570
box -8 -3 16 105
use FILL  FILL_4944
timestamp 1745462530
transform 1 0 1096 0 1 570
box -8 -3 16 105
use FILL  FILL_4945
timestamp 1745462530
transform 1 0 1048 0 1 570
box -8 -3 16 105
use FILL  FILL_4946
timestamp 1745462530
transform 1 0 944 0 1 570
box -8 -3 16 105
use FILL  FILL_4947
timestamp 1745462530
transform 1 0 840 0 1 570
box -8 -3 16 105
use FILL  FILL_4948
timestamp 1745462530
transform 1 0 808 0 1 570
box -8 -3 16 105
use FILL  FILL_4949
timestamp 1745462530
transform 1 0 760 0 1 570
box -8 -3 16 105
use FILL  FILL_4950
timestamp 1745462530
transform 1 0 752 0 1 570
box -8 -3 16 105
use FILL  FILL_4951
timestamp 1745462530
transform 1 0 632 0 1 570
box -8 -3 16 105
use FILL  FILL_4952
timestamp 1745462530
transform 1 0 624 0 1 570
box -8 -3 16 105
use FILL  FILL_4953
timestamp 1745462530
transform 1 0 560 0 1 570
box -8 -3 16 105
use FILL  FILL_4954
timestamp 1745462530
transform 1 0 552 0 1 570
box -8 -3 16 105
use FILL  FILL_4955
timestamp 1745462530
transform 1 0 544 0 1 570
box -8 -3 16 105
use FILL  FILL_4956
timestamp 1745462530
transform 1 0 456 0 1 570
box -8 -3 16 105
use FILL  FILL_4957
timestamp 1745462530
transform 1 0 448 0 1 570
box -8 -3 16 105
use FILL  FILL_4958
timestamp 1745462530
transform 1 0 408 0 1 570
box -8 -3 16 105
use FILL  FILL_4959
timestamp 1745462530
transform 1 0 360 0 1 570
box -8 -3 16 105
use FILL  FILL_4960
timestamp 1745462530
transform 1 0 352 0 1 570
box -8 -3 16 105
use FILL  FILL_4961
timestamp 1745462530
transform 1 0 288 0 1 570
box -8 -3 16 105
use FILL  FILL_4962
timestamp 1745462530
transform 1 0 280 0 1 570
box -8 -3 16 105
use FILL  FILL_4963
timestamp 1745462530
transform 1 0 232 0 1 570
box -8 -3 16 105
use FILL  FILL_4964
timestamp 1745462530
transform 1 0 184 0 1 570
box -8 -3 16 105
use FILL  FILL_4965
timestamp 1745462530
transform 1 0 176 0 1 570
box -8 -3 16 105
use FILL  FILL_4966
timestamp 1745462530
transform 1 0 72 0 1 570
box -8 -3 16 105
use FILL  FILL_4967
timestamp 1745462530
transform 1 0 4272 0 -1 570
box -8 -3 16 105
use FILL  FILL_4968
timestamp 1745462530
transform 1 0 4248 0 -1 570
box -8 -3 16 105
use FILL  FILL_4969
timestamp 1745462530
transform 1 0 4200 0 -1 570
box -8 -3 16 105
use FILL  FILL_4970
timestamp 1745462530
transform 1 0 4080 0 -1 570
box -8 -3 16 105
use FILL  FILL_4971
timestamp 1745462530
transform 1 0 3976 0 -1 570
box -8 -3 16 105
use FILL  FILL_4972
timestamp 1745462530
transform 1 0 3952 0 -1 570
box -8 -3 16 105
use FILL  FILL_4973
timestamp 1745462530
transform 1 0 3944 0 -1 570
box -8 -3 16 105
use FILL  FILL_4974
timestamp 1745462530
transform 1 0 3896 0 -1 570
box -8 -3 16 105
use FILL  FILL_4975
timestamp 1745462530
transform 1 0 3888 0 -1 570
box -8 -3 16 105
use FILL  FILL_4976
timestamp 1745462530
transform 1 0 3880 0 -1 570
box -8 -3 16 105
use FILL  FILL_4977
timestamp 1745462530
transform 1 0 3832 0 -1 570
box -8 -3 16 105
use FILL  FILL_4978
timestamp 1745462530
transform 1 0 3824 0 -1 570
box -8 -3 16 105
use FILL  FILL_4979
timestamp 1745462530
transform 1 0 3784 0 -1 570
box -8 -3 16 105
use FILL  FILL_4980
timestamp 1745462530
transform 1 0 3776 0 -1 570
box -8 -3 16 105
use FILL  FILL_4981
timestamp 1745462530
transform 1 0 3672 0 -1 570
box -8 -3 16 105
use FILL  FILL_4982
timestamp 1745462530
transform 1 0 3648 0 -1 570
box -8 -3 16 105
use FILL  FILL_4983
timestamp 1745462530
transform 1 0 3640 0 -1 570
box -8 -3 16 105
use FILL  FILL_4984
timestamp 1745462530
transform 1 0 3592 0 -1 570
box -8 -3 16 105
use FILL  FILL_4985
timestamp 1745462530
transform 1 0 3584 0 -1 570
box -8 -3 16 105
use FILL  FILL_4986
timestamp 1745462530
transform 1 0 3576 0 -1 570
box -8 -3 16 105
use FILL  FILL_4987
timestamp 1745462530
transform 1 0 3536 0 -1 570
box -8 -3 16 105
use FILL  FILL_4988
timestamp 1745462530
transform 1 0 3496 0 -1 570
box -8 -3 16 105
use FILL  FILL_4989
timestamp 1745462530
transform 1 0 3488 0 -1 570
box -8 -3 16 105
use FILL  FILL_4990
timestamp 1745462530
transform 1 0 3480 0 -1 570
box -8 -3 16 105
use FILL  FILL_4991
timestamp 1745462530
transform 1 0 3432 0 -1 570
box -8 -3 16 105
use FILL  FILL_4992
timestamp 1745462530
transform 1 0 3408 0 -1 570
box -8 -3 16 105
use FILL  FILL_4993
timestamp 1745462530
transform 1 0 3400 0 -1 570
box -8 -3 16 105
use FILL  FILL_4994
timestamp 1745462530
transform 1 0 3352 0 -1 570
box -8 -3 16 105
use FILL  FILL_4995
timestamp 1745462530
transform 1 0 3344 0 -1 570
box -8 -3 16 105
use FILL  FILL_4996
timestamp 1745462530
transform 1 0 3336 0 -1 570
box -8 -3 16 105
use FILL  FILL_4997
timestamp 1745462530
transform 1 0 3304 0 -1 570
box -8 -3 16 105
use FILL  FILL_4998
timestamp 1745462530
transform 1 0 3256 0 -1 570
box -8 -3 16 105
use FILL  FILL_4999
timestamp 1745462530
transform 1 0 3248 0 -1 570
box -8 -3 16 105
use FILL  FILL_5000
timestamp 1745462530
transform 1 0 3240 0 -1 570
box -8 -3 16 105
use FILL  FILL_5001
timestamp 1745462530
transform 1 0 3192 0 -1 570
box -8 -3 16 105
use FILL  FILL_5002
timestamp 1745462530
transform 1 0 3168 0 -1 570
box -8 -3 16 105
use FILL  FILL_5003
timestamp 1745462530
transform 1 0 3160 0 -1 570
box -8 -3 16 105
use FILL  FILL_5004
timestamp 1745462530
transform 1 0 3056 0 -1 570
box -8 -3 16 105
use FILL  FILL_5005
timestamp 1745462530
transform 1 0 3032 0 -1 570
box -8 -3 16 105
use FILL  FILL_5006
timestamp 1745462530
transform 1 0 2984 0 -1 570
box -8 -3 16 105
use FILL  FILL_5007
timestamp 1745462530
transform 1 0 2976 0 -1 570
box -8 -3 16 105
use FILL  FILL_5008
timestamp 1745462530
transform 1 0 2968 0 -1 570
box -8 -3 16 105
use FILL  FILL_5009
timestamp 1745462530
transform 1 0 2920 0 -1 570
box -8 -3 16 105
use FILL  FILL_5010
timestamp 1745462530
transform 1 0 2912 0 -1 570
box -8 -3 16 105
use FILL  FILL_5011
timestamp 1745462530
transform 1 0 2864 0 -1 570
box -8 -3 16 105
use FILL  FILL_5012
timestamp 1745462530
transform 1 0 2816 0 -1 570
box -8 -3 16 105
use FILL  FILL_5013
timestamp 1745462530
transform 1 0 2808 0 -1 570
box -8 -3 16 105
use FILL  FILL_5014
timestamp 1745462530
transform 1 0 2800 0 -1 570
box -8 -3 16 105
use FILL  FILL_5015
timestamp 1745462530
transform 1 0 2736 0 -1 570
box -8 -3 16 105
use FILL  FILL_5016
timestamp 1745462530
transform 1 0 2728 0 -1 570
box -8 -3 16 105
use FILL  FILL_5017
timestamp 1745462530
transform 1 0 2680 0 -1 570
box -8 -3 16 105
use FILL  FILL_5018
timestamp 1745462530
transform 1 0 2640 0 -1 570
box -8 -3 16 105
use FILL  FILL_5019
timestamp 1745462530
transform 1 0 2600 0 -1 570
box -8 -3 16 105
use FILL  FILL_5020
timestamp 1745462530
transform 1 0 2560 0 -1 570
box -8 -3 16 105
use FILL  FILL_5021
timestamp 1745462530
transform 1 0 2552 0 -1 570
box -8 -3 16 105
use FILL  FILL_5022
timestamp 1745462530
transform 1 0 2544 0 -1 570
box -8 -3 16 105
use FILL  FILL_5023
timestamp 1745462530
transform 1 0 2496 0 -1 570
box -8 -3 16 105
use FILL  FILL_5024
timestamp 1745462530
transform 1 0 2488 0 -1 570
box -8 -3 16 105
use FILL  FILL_5025
timestamp 1745462530
transform 1 0 2440 0 -1 570
box -8 -3 16 105
use FILL  FILL_5026
timestamp 1745462530
transform 1 0 2432 0 -1 570
box -8 -3 16 105
use FILL  FILL_5027
timestamp 1745462530
transform 1 0 2424 0 -1 570
box -8 -3 16 105
use FILL  FILL_5028
timestamp 1745462530
transform 1 0 2376 0 -1 570
box -8 -3 16 105
use FILL  FILL_5029
timestamp 1745462530
transform 1 0 2368 0 -1 570
box -8 -3 16 105
use FILL  FILL_5030
timestamp 1745462530
transform 1 0 2328 0 -1 570
box -8 -3 16 105
use FILL  FILL_5031
timestamp 1745462530
transform 1 0 2320 0 -1 570
box -8 -3 16 105
use FILL  FILL_5032
timestamp 1745462530
transform 1 0 2272 0 -1 570
box -8 -3 16 105
use FILL  FILL_5033
timestamp 1745462530
transform 1 0 2264 0 -1 570
box -8 -3 16 105
use FILL  FILL_5034
timestamp 1745462530
transform 1 0 2256 0 -1 570
box -8 -3 16 105
use FILL  FILL_5035
timestamp 1745462530
transform 1 0 2208 0 -1 570
box -8 -3 16 105
use FILL  FILL_5036
timestamp 1745462530
transform 1 0 2200 0 -1 570
box -8 -3 16 105
use FILL  FILL_5037
timestamp 1745462530
transform 1 0 2192 0 -1 570
box -8 -3 16 105
use FILL  FILL_5038
timestamp 1745462530
transform 1 0 2088 0 -1 570
box -8 -3 16 105
use FILL  FILL_5039
timestamp 1745462530
transform 1 0 2080 0 -1 570
box -8 -3 16 105
use FILL  FILL_5040
timestamp 1745462530
transform 1 0 2056 0 -1 570
box -8 -3 16 105
use FILL  FILL_5041
timestamp 1745462530
transform 1 0 2024 0 -1 570
box -8 -3 16 105
use FILL  FILL_5042
timestamp 1745462530
transform 1 0 2016 0 -1 570
box -8 -3 16 105
use FILL  FILL_5043
timestamp 1745462530
transform 1 0 2008 0 -1 570
box -8 -3 16 105
use FILL  FILL_5044
timestamp 1745462530
transform 1 0 1968 0 -1 570
box -8 -3 16 105
use FILL  FILL_5045
timestamp 1745462530
transform 1 0 1960 0 -1 570
box -8 -3 16 105
use FILL  FILL_5046
timestamp 1745462530
transform 1 0 1912 0 -1 570
box -8 -3 16 105
use FILL  FILL_5047
timestamp 1745462530
transform 1 0 1904 0 -1 570
box -8 -3 16 105
use FILL  FILL_5048
timestamp 1745462530
transform 1 0 1896 0 -1 570
box -8 -3 16 105
use FILL  FILL_5049
timestamp 1745462530
transform 1 0 1888 0 -1 570
box -8 -3 16 105
use FILL  FILL_5050
timestamp 1745462530
transform 1 0 1840 0 -1 570
box -8 -3 16 105
use FILL  FILL_5051
timestamp 1745462530
transform 1 0 1832 0 -1 570
box -8 -3 16 105
use FILL  FILL_5052
timestamp 1745462530
transform 1 0 1712 0 -1 570
box -8 -3 16 105
use FILL  FILL_5053
timestamp 1745462530
transform 1 0 1704 0 -1 570
box -8 -3 16 105
use FILL  FILL_5054
timestamp 1745462530
transform 1 0 1656 0 -1 570
box -8 -3 16 105
use FILL  FILL_5055
timestamp 1745462530
transform 1 0 1648 0 -1 570
box -8 -3 16 105
use FILL  FILL_5056
timestamp 1745462530
transform 1 0 1640 0 -1 570
box -8 -3 16 105
use FILL  FILL_5057
timestamp 1745462530
transform 1 0 1592 0 -1 570
box -8 -3 16 105
use FILL  FILL_5058
timestamp 1745462530
transform 1 0 1584 0 -1 570
box -8 -3 16 105
use FILL  FILL_5059
timestamp 1745462530
transform 1 0 1480 0 -1 570
box -8 -3 16 105
use FILL  FILL_5060
timestamp 1745462530
transform 1 0 1456 0 -1 570
box -8 -3 16 105
use FILL  FILL_5061
timestamp 1745462530
transform 1 0 1408 0 -1 570
box -8 -3 16 105
use FILL  FILL_5062
timestamp 1745462530
transform 1 0 1400 0 -1 570
box -8 -3 16 105
use FILL  FILL_5063
timestamp 1745462530
transform 1 0 1392 0 -1 570
box -8 -3 16 105
use FILL  FILL_5064
timestamp 1745462530
transform 1 0 1384 0 -1 570
box -8 -3 16 105
use FILL  FILL_5065
timestamp 1745462530
transform 1 0 1336 0 -1 570
box -8 -3 16 105
use FILL  FILL_5066
timestamp 1745462530
transform 1 0 1328 0 -1 570
box -8 -3 16 105
use FILL  FILL_5067
timestamp 1745462530
transform 1 0 1320 0 -1 570
box -8 -3 16 105
use FILL  FILL_5068
timestamp 1745462530
transform 1 0 1280 0 -1 570
box -8 -3 16 105
use FILL  FILL_5069
timestamp 1745462530
transform 1 0 1272 0 -1 570
box -8 -3 16 105
use FILL  FILL_5070
timestamp 1745462530
transform 1 0 1264 0 -1 570
box -8 -3 16 105
use FILL  FILL_5071
timestamp 1745462530
transform 1 0 1224 0 -1 570
box -8 -3 16 105
use FILL  FILL_5072
timestamp 1745462530
transform 1 0 1216 0 -1 570
box -8 -3 16 105
use FILL  FILL_5073
timestamp 1745462530
transform 1 0 1208 0 -1 570
box -8 -3 16 105
use FILL  FILL_5074
timestamp 1745462530
transform 1 0 1200 0 -1 570
box -8 -3 16 105
use FILL  FILL_5075
timestamp 1745462530
transform 1 0 1152 0 -1 570
box -8 -3 16 105
use FILL  FILL_5076
timestamp 1745462530
transform 1 0 1144 0 -1 570
box -8 -3 16 105
use FILL  FILL_5077
timestamp 1745462530
transform 1 0 1136 0 -1 570
box -8 -3 16 105
use FILL  FILL_5078
timestamp 1745462530
transform 1 0 1128 0 -1 570
box -8 -3 16 105
use FILL  FILL_5079
timestamp 1745462530
transform 1 0 1080 0 -1 570
box -8 -3 16 105
use FILL  FILL_5080
timestamp 1745462530
transform 1 0 1072 0 -1 570
box -8 -3 16 105
use FILL  FILL_5081
timestamp 1745462530
transform 1 0 1064 0 -1 570
box -8 -3 16 105
use FILL  FILL_5082
timestamp 1745462530
transform 1 0 1056 0 -1 570
box -8 -3 16 105
use FILL  FILL_5083
timestamp 1745462530
transform 1 0 1008 0 -1 570
box -8 -3 16 105
use FILL  FILL_5084
timestamp 1745462530
transform 1 0 1000 0 -1 570
box -8 -3 16 105
use FILL  FILL_5085
timestamp 1745462530
transform 1 0 992 0 -1 570
box -8 -3 16 105
use FILL  FILL_5086
timestamp 1745462530
transform 1 0 952 0 -1 570
box -8 -3 16 105
use FILL  FILL_5087
timestamp 1745462530
transform 1 0 944 0 -1 570
box -8 -3 16 105
use FILL  FILL_5088
timestamp 1745462530
transform 1 0 896 0 -1 570
box -8 -3 16 105
use FILL  FILL_5089
timestamp 1745462530
transform 1 0 888 0 -1 570
box -8 -3 16 105
use FILL  FILL_5090
timestamp 1745462530
transform 1 0 824 0 -1 570
box -8 -3 16 105
use FILL  FILL_5091
timestamp 1745462530
transform 1 0 816 0 -1 570
box -8 -3 16 105
use FILL  FILL_5092
timestamp 1745462530
transform 1 0 712 0 -1 570
box -8 -3 16 105
use FILL  FILL_5093
timestamp 1745462530
transform 1 0 664 0 -1 570
box -8 -3 16 105
use FILL  FILL_5094
timestamp 1745462530
transform 1 0 656 0 -1 570
box -8 -3 16 105
use FILL  FILL_5095
timestamp 1745462530
transform 1 0 552 0 -1 570
box -8 -3 16 105
use FILL  FILL_5096
timestamp 1745462530
transform 1 0 544 0 -1 570
box -8 -3 16 105
use FILL  FILL_5097
timestamp 1745462530
transform 1 0 504 0 -1 570
box -8 -3 16 105
use FILL  FILL_5098
timestamp 1745462530
transform 1 0 496 0 -1 570
box -8 -3 16 105
use FILL  FILL_5099
timestamp 1745462530
transform 1 0 448 0 -1 570
box -8 -3 16 105
use FILL  FILL_5100
timestamp 1745462530
transform 1 0 440 0 -1 570
box -8 -3 16 105
use FILL  FILL_5101
timestamp 1745462530
transform 1 0 400 0 -1 570
box -8 -3 16 105
use FILL  FILL_5102
timestamp 1745462530
transform 1 0 392 0 -1 570
box -8 -3 16 105
use FILL  FILL_5103
timestamp 1745462530
transform 1 0 344 0 -1 570
box -8 -3 16 105
use FILL  FILL_5104
timestamp 1745462530
transform 1 0 336 0 -1 570
box -8 -3 16 105
use FILL  FILL_5105
timestamp 1745462530
transform 1 0 288 0 -1 570
box -8 -3 16 105
use FILL  FILL_5106
timestamp 1745462530
transform 1 0 280 0 -1 570
box -8 -3 16 105
use FILL  FILL_5107
timestamp 1745462530
transform 1 0 272 0 -1 570
box -8 -3 16 105
use FILL  FILL_5108
timestamp 1745462530
transform 1 0 264 0 -1 570
box -8 -3 16 105
use FILL  FILL_5109
timestamp 1745462530
transform 1 0 216 0 -1 570
box -8 -3 16 105
use FILL  FILL_5110
timestamp 1745462530
transform 1 0 192 0 -1 570
box -8 -3 16 105
use FILL  FILL_5111
timestamp 1745462530
transform 1 0 184 0 -1 570
box -8 -3 16 105
use FILL  FILL_5112
timestamp 1745462530
transform 1 0 80 0 -1 570
box -8 -3 16 105
use FILL  FILL_5113
timestamp 1745462530
transform 1 0 72 0 -1 570
box -8 -3 16 105
use FILL  FILL_5114
timestamp 1745462530
transform 1 0 4368 0 1 370
box -8 -3 16 105
use FILL  FILL_5115
timestamp 1745462530
transform 1 0 4248 0 1 370
box -8 -3 16 105
use FILL  FILL_5116
timestamp 1745462530
transform 1 0 4200 0 1 370
box -8 -3 16 105
use FILL  FILL_5117
timestamp 1745462530
transform 1 0 4192 0 1 370
box -8 -3 16 105
use FILL  FILL_5118
timestamp 1745462530
transform 1 0 4184 0 1 370
box -8 -3 16 105
use FILL  FILL_5119
timestamp 1745462530
transform 1 0 4136 0 1 370
box -8 -3 16 105
use FILL  FILL_5120
timestamp 1745462530
transform 1 0 4112 0 1 370
box -8 -3 16 105
use FILL  FILL_5121
timestamp 1745462530
transform 1 0 4104 0 1 370
box -8 -3 16 105
use FILL  FILL_5122
timestamp 1745462530
transform 1 0 4056 0 1 370
box -8 -3 16 105
use FILL  FILL_5123
timestamp 1745462530
transform 1 0 4048 0 1 370
box -8 -3 16 105
use FILL  FILL_5124
timestamp 1745462530
transform 1 0 4040 0 1 370
box -8 -3 16 105
use FILL  FILL_5125
timestamp 1745462530
transform 1 0 3992 0 1 370
box -8 -3 16 105
use FILL  FILL_5126
timestamp 1745462530
transform 1 0 3984 0 1 370
box -8 -3 16 105
use FILL  FILL_5127
timestamp 1745462530
transform 1 0 3960 0 1 370
box -8 -3 16 105
use FILL  FILL_5128
timestamp 1745462530
transform 1 0 3952 0 1 370
box -8 -3 16 105
use FILL  FILL_5129
timestamp 1745462530
transform 1 0 3944 0 1 370
box -8 -3 16 105
use FILL  FILL_5130
timestamp 1745462530
transform 1 0 3896 0 1 370
box -8 -3 16 105
use FILL  FILL_5131
timestamp 1745462530
transform 1 0 3888 0 1 370
box -8 -3 16 105
use FILL  FILL_5132
timestamp 1745462530
transform 1 0 3880 0 1 370
box -8 -3 16 105
use FILL  FILL_5133
timestamp 1745462530
transform 1 0 3848 0 1 370
box -8 -3 16 105
use FILL  FILL_5134
timestamp 1745462530
transform 1 0 3840 0 1 370
box -8 -3 16 105
use FILL  FILL_5135
timestamp 1745462530
transform 1 0 3792 0 1 370
box -8 -3 16 105
use FILL  FILL_5136
timestamp 1745462530
transform 1 0 3784 0 1 370
box -8 -3 16 105
use FILL  FILL_5137
timestamp 1745462530
transform 1 0 3776 0 1 370
box -8 -3 16 105
use FILL  FILL_5138
timestamp 1745462530
transform 1 0 3768 0 1 370
box -8 -3 16 105
use FILL  FILL_5139
timestamp 1745462530
transform 1 0 3720 0 1 370
box -8 -3 16 105
use FILL  FILL_5140
timestamp 1745462530
transform 1 0 3712 0 1 370
box -8 -3 16 105
use FILL  FILL_5141
timestamp 1745462530
transform 1 0 3704 0 1 370
box -8 -3 16 105
use FILL  FILL_5142
timestamp 1745462530
transform 1 0 3656 0 1 370
box -8 -3 16 105
use FILL  FILL_5143
timestamp 1745462530
transform 1 0 3648 0 1 370
box -8 -3 16 105
use FILL  FILL_5144
timestamp 1745462530
transform 1 0 3640 0 1 370
box -8 -3 16 105
use FILL  FILL_5145
timestamp 1745462530
transform 1 0 3608 0 1 370
box -8 -3 16 105
use FILL  FILL_5146
timestamp 1745462530
transform 1 0 3568 0 1 370
box -8 -3 16 105
use FILL  FILL_5147
timestamp 1745462530
transform 1 0 3560 0 1 370
box -8 -3 16 105
use FILL  FILL_5148
timestamp 1745462530
transform 1 0 3552 0 1 370
box -8 -3 16 105
use FILL  FILL_5149
timestamp 1745462530
transform 1 0 3504 0 1 370
box -8 -3 16 105
use FILL  FILL_5150
timestamp 1745462530
transform 1 0 3496 0 1 370
box -8 -3 16 105
use FILL  FILL_5151
timestamp 1745462530
transform 1 0 3392 0 1 370
box -8 -3 16 105
use FILL  FILL_5152
timestamp 1745462530
transform 1 0 3384 0 1 370
box -8 -3 16 105
use FILL  FILL_5153
timestamp 1745462530
transform 1 0 3336 0 1 370
box -8 -3 16 105
use FILL  FILL_5154
timestamp 1745462530
transform 1 0 3328 0 1 370
box -8 -3 16 105
use FILL  FILL_5155
timestamp 1745462530
transform 1 0 3208 0 1 370
box -8 -3 16 105
use FILL  FILL_5156
timestamp 1745462530
transform 1 0 3200 0 1 370
box -8 -3 16 105
use FILL  FILL_5157
timestamp 1745462530
transform 1 0 3096 0 1 370
box -8 -3 16 105
use FILL  FILL_5158
timestamp 1745462530
transform 1 0 3088 0 1 370
box -8 -3 16 105
use FILL  FILL_5159
timestamp 1745462530
transform 1 0 2984 0 1 370
box -8 -3 16 105
use FILL  FILL_5160
timestamp 1745462530
transform 1 0 2960 0 1 370
box -8 -3 16 105
use FILL  FILL_5161
timestamp 1745462530
transform 1 0 2912 0 1 370
box -8 -3 16 105
use FILL  FILL_5162
timestamp 1745462530
transform 1 0 2904 0 1 370
box -8 -3 16 105
use FILL  FILL_5163
timestamp 1745462530
transform 1 0 2896 0 1 370
box -8 -3 16 105
use FILL  FILL_5164
timestamp 1745462530
transform 1 0 2872 0 1 370
box -8 -3 16 105
use FILL  FILL_5165
timestamp 1745462530
transform 1 0 2824 0 1 370
box -8 -3 16 105
use FILL  FILL_5166
timestamp 1745462530
transform 1 0 2816 0 1 370
box -8 -3 16 105
use FILL  FILL_5167
timestamp 1745462530
transform 1 0 2808 0 1 370
box -8 -3 16 105
use FILL  FILL_5168
timestamp 1745462530
transform 1 0 2704 0 1 370
box -8 -3 16 105
use FILL  FILL_5169
timestamp 1745462530
transform 1 0 2680 0 1 370
box -8 -3 16 105
use FILL  FILL_5170
timestamp 1745462530
transform 1 0 2576 0 1 370
box -8 -3 16 105
use FILL  FILL_5171
timestamp 1745462530
transform 1 0 2568 0 1 370
box -8 -3 16 105
use FILL  FILL_5172
timestamp 1745462530
transform 1 0 2544 0 1 370
box -8 -3 16 105
use FILL  FILL_5173
timestamp 1745462530
transform 1 0 2440 0 1 370
box -8 -3 16 105
use FILL  FILL_5174
timestamp 1745462530
transform 1 0 2336 0 1 370
box -8 -3 16 105
use FILL  FILL_5175
timestamp 1745462530
transform 1 0 2328 0 1 370
box -8 -3 16 105
use FILL  FILL_5176
timestamp 1745462530
transform 1 0 2280 0 1 370
box -8 -3 16 105
use FILL  FILL_5177
timestamp 1745462530
transform 1 0 2272 0 1 370
box -8 -3 16 105
use FILL  FILL_5178
timestamp 1745462530
transform 1 0 2264 0 1 370
box -8 -3 16 105
use FILL  FILL_5179
timestamp 1745462530
transform 1 0 2216 0 1 370
box -8 -3 16 105
use FILL  FILL_5180
timestamp 1745462530
transform 1 0 2208 0 1 370
box -8 -3 16 105
use FILL  FILL_5181
timestamp 1745462530
transform 1 0 2184 0 1 370
box -8 -3 16 105
use FILL  FILL_5182
timestamp 1745462530
transform 1 0 2080 0 1 370
box -8 -3 16 105
use FILL  FILL_5183
timestamp 1745462530
transform 1 0 2072 0 1 370
box -8 -3 16 105
use FILL  FILL_5184
timestamp 1745462530
transform 1 0 1968 0 1 370
box -8 -3 16 105
use FILL  FILL_5185
timestamp 1745462530
transform 1 0 1960 0 1 370
box -8 -3 16 105
use FILL  FILL_5186
timestamp 1745462530
transform 1 0 1952 0 1 370
box -8 -3 16 105
use FILL  FILL_5187
timestamp 1745462530
transform 1 0 1904 0 1 370
box -8 -3 16 105
use FILL  FILL_5188
timestamp 1745462530
transform 1 0 1896 0 1 370
box -8 -3 16 105
use FILL  FILL_5189
timestamp 1745462530
transform 1 0 1888 0 1 370
box -8 -3 16 105
use FILL  FILL_5190
timestamp 1745462530
transform 1 0 1864 0 1 370
box -8 -3 16 105
use FILL  FILL_5191
timestamp 1745462530
transform 1 0 1816 0 1 370
box -8 -3 16 105
use FILL  FILL_5192
timestamp 1745462530
transform 1 0 1808 0 1 370
box -8 -3 16 105
use FILL  FILL_5193
timestamp 1745462530
transform 1 0 1800 0 1 370
box -8 -3 16 105
use FILL  FILL_5194
timestamp 1745462530
transform 1 0 1696 0 1 370
box -8 -3 16 105
use FILL  FILL_5195
timestamp 1745462530
transform 1 0 1688 0 1 370
box -8 -3 16 105
use FILL  FILL_5196
timestamp 1745462530
transform 1 0 1640 0 1 370
box -8 -3 16 105
use FILL  FILL_5197
timestamp 1745462530
transform 1 0 1632 0 1 370
box -8 -3 16 105
use FILL  FILL_5198
timestamp 1745462530
transform 1 0 1624 0 1 370
box -8 -3 16 105
use FILL  FILL_5199
timestamp 1745462530
transform 1 0 1504 0 1 370
box -8 -3 16 105
use FILL  FILL_5200
timestamp 1745462530
transform 1 0 1496 0 1 370
box -8 -3 16 105
use FILL  FILL_5201
timestamp 1745462530
transform 1 0 1488 0 1 370
box -8 -3 16 105
use FILL  FILL_5202
timestamp 1745462530
transform 1 0 1448 0 1 370
box -8 -3 16 105
use FILL  FILL_5203
timestamp 1745462530
transform 1 0 1440 0 1 370
box -8 -3 16 105
use FILL  FILL_5204
timestamp 1745462530
transform 1 0 1336 0 1 370
box -8 -3 16 105
use FILL  FILL_5205
timestamp 1745462530
transform 1 0 1328 0 1 370
box -8 -3 16 105
use FILL  FILL_5206
timestamp 1745462530
transform 1 0 1224 0 1 370
box -8 -3 16 105
use FILL  FILL_5207
timestamp 1745462530
transform 1 0 1200 0 1 370
box -8 -3 16 105
use FILL  FILL_5208
timestamp 1745462530
transform 1 0 1192 0 1 370
box -8 -3 16 105
use FILL  FILL_5209
timestamp 1745462530
transform 1 0 1184 0 1 370
box -8 -3 16 105
use FILL  FILL_5210
timestamp 1745462530
transform 1 0 1136 0 1 370
box -8 -3 16 105
use FILL  FILL_5211
timestamp 1745462530
transform 1 0 1128 0 1 370
box -8 -3 16 105
use FILL  FILL_5212
timestamp 1745462530
transform 1 0 1120 0 1 370
box -8 -3 16 105
use FILL  FILL_5213
timestamp 1745462530
transform 1 0 1096 0 1 370
box -8 -3 16 105
use FILL  FILL_5214
timestamp 1745462530
transform 1 0 992 0 1 370
box -8 -3 16 105
use FILL  FILL_5215
timestamp 1745462530
transform 1 0 984 0 1 370
box -8 -3 16 105
use FILL  FILL_5216
timestamp 1745462530
transform 1 0 976 0 1 370
box -8 -3 16 105
use FILL  FILL_5217
timestamp 1745462530
transform 1 0 872 0 1 370
box -8 -3 16 105
use FILL  FILL_5218
timestamp 1745462530
transform 1 0 864 0 1 370
box -8 -3 16 105
use FILL  FILL_5219
timestamp 1745462530
transform 1 0 856 0 1 370
box -8 -3 16 105
use FILL  FILL_5220
timestamp 1745462530
transform 1 0 752 0 1 370
box -8 -3 16 105
use FILL  FILL_5221
timestamp 1745462530
transform 1 0 744 0 1 370
box -8 -3 16 105
use FILL  FILL_5222
timestamp 1745462530
transform 1 0 736 0 1 370
box -8 -3 16 105
use FILL  FILL_5223
timestamp 1745462530
transform 1 0 672 0 1 370
box -8 -3 16 105
use FILL  FILL_5224
timestamp 1745462530
transform 1 0 664 0 1 370
box -8 -3 16 105
use FILL  FILL_5225
timestamp 1745462530
transform 1 0 656 0 1 370
box -8 -3 16 105
use FILL  FILL_5226
timestamp 1745462530
transform 1 0 552 0 1 370
box -8 -3 16 105
use FILL  FILL_5227
timestamp 1745462530
transform 1 0 544 0 1 370
box -8 -3 16 105
use FILL  FILL_5228
timestamp 1745462530
transform 1 0 520 0 1 370
box -8 -3 16 105
use FILL  FILL_5229
timestamp 1745462530
transform 1 0 512 0 1 370
box -8 -3 16 105
use FILL  FILL_5230
timestamp 1745462530
transform 1 0 464 0 1 370
box -8 -3 16 105
use FILL  FILL_5231
timestamp 1745462530
transform 1 0 456 0 1 370
box -8 -3 16 105
use FILL  FILL_5232
timestamp 1745462530
transform 1 0 432 0 1 370
box -8 -3 16 105
use FILL  FILL_5233
timestamp 1745462530
transform 1 0 384 0 1 370
box -8 -3 16 105
use FILL  FILL_5234
timestamp 1745462530
transform 1 0 376 0 1 370
box -8 -3 16 105
use FILL  FILL_5235
timestamp 1745462530
transform 1 0 352 0 1 370
box -8 -3 16 105
use FILL  FILL_5236
timestamp 1745462530
transform 1 0 304 0 1 370
box -8 -3 16 105
use FILL  FILL_5237
timestamp 1745462530
transform 1 0 296 0 1 370
box -8 -3 16 105
use FILL  FILL_5238
timestamp 1745462530
transform 1 0 288 0 1 370
box -8 -3 16 105
use FILL  FILL_5239
timestamp 1745462530
transform 1 0 248 0 1 370
box -8 -3 16 105
use FILL  FILL_5240
timestamp 1745462530
transform 1 0 240 0 1 370
box -8 -3 16 105
use FILL  FILL_5241
timestamp 1745462530
transform 1 0 192 0 1 370
box -8 -3 16 105
use FILL  FILL_5242
timestamp 1745462530
transform 1 0 184 0 1 370
box -8 -3 16 105
use FILL  FILL_5243
timestamp 1745462530
transform 1 0 80 0 1 370
box -8 -3 16 105
use FILL  FILL_5244
timestamp 1745462530
transform 1 0 72 0 1 370
box -8 -3 16 105
use FILL  FILL_5245
timestamp 1745462530
transform 1 0 4352 0 -1 370
box -8 -3 16 105
use FILL  FILL_5246
timestamp 1745462530
transform 1 0 4344 0 -1 370
box -8 -3 16 105
use FILL  FILL_5247
timestamp 1745462530
transform 1 0 4336 0 -1 370
box -8 -3 16 105
use FILL  FILL_5248
timestamp 1745462530
transform 1 0 4288 0 -1 370
box -8 -3 16 105
use FILL  FILL_5249
timestamp 1745462530
transform 1 0 4280 0 -1 370
box -8 -3 16 105
use FILL  FILL_5250
timestamp 1745462530
transform 1 0 4256 0 -1 370
box -8 -3 16 105
use FILL  FILL_5251
timestamp 1745462530
transform 1 0 4248 0 -1 370
box -8 -3 16 105
use FILL  FILL_5252
timestamp 1745462530
transform 1 0 4144 0 -1 370
box -8 -3 16 105
use FILL  FILL_5253
timestamp 1745462530
transform 1 0 4136 0 -1 370
box -8 -3 16 105
use FILL  FILL_5254
timestamp 1745462530
transform 1 0 4032 0 -1 370
box -8 -3 16 105
use FILL  FILL_5255
timestamp 1745462530
transform 1 0 4024 0 -1 370
box -8 -3 16 105
use FILL  FILL_5256
timestamp 1745462530
transform 1 0 4016 0 -1 370
box -8 -3 16 105
use FILL  FILL_5257
timestamp 1745462530
transform 1 0 3968 0 -1 370
box -8 -3 16 105
use FILL  FILL_5258
timestamp 1745462530
transform 1 0 3960 0 -1 370
box -8 -3 16 105
use FILL  FILL_5259
timestamp 1745462530
transform 1 0 3952 0 -1 370
box -8 -3 16 105
use FILL  FILL_5260
timestamp 1745462530
transform 1 0 3944 0 -1 370
box -8 -3 16 105
use FILL  FILL_5261
timestamp 1745462530
transform 1 0 3896 0 -1 370
box -8 -3 16 105
use FILL  FILL_5262
timestamp 1745462530
transform 1 0 3888 0 -1 370
box -8 -3 16 105
use FILL  FILL_5263
timestamp 1745462530
transform 1 0 3880 0 -1 370
box -8 -3 16 105
use FILL  FILL_5264
timestamp 1745462530
transform 1 0 3848 0 -1 370
box -8 -3 16 105
use FILL  FILL_5265
timestamp 1745462530
transform 1 0 3840 0 -1 370
box -8 -3 16 105
use FILL  FILL_5266
timestamp 1745462530
transform 1 0 3800 0 -1 370
box -8 -3 16 105
use FILL  FILL_5267
timestamp 1745462530
transform 1 0 3792 0 -1 370
box -8 -3 16 105
use FILL  FILL_5268
timestamp 1745462530
transform 1 0 3744 0 -1 370
box -8 -3 16 105
use FILL  FILL_5269
timestamp 1745462530
transform 1 0 3736 0 -1 370
box -8 -3 16 105
use FILL  FILL_5270
timestamp 1745462530
transform 1 0 3728 0 -1 370
box -8 -3 16 105
use FILL  FILL_5271
timestamp 1745462530
transform 1 0 3720 0 -1 370
box -8 -3 16 105
use FILL  FILL_5272
timestamp 1745462530
transform 1 0 3680 0 -1 370
box -8 -3 16 105
use FILL  FILL_5273
timestamp 1745462530
transform 1 0 3672 0 -1 370
box -8 -3 16 105
use FILL  FILL_5274
timestamp 1745462530
transform 1 0 3624 0 -1 370
box -8 -3 16 105
use FILL  FILL_5275
timestamp 1745462530
transform 1 0 3616 0 -1 370
box -8 -3 16 105
use FILL  FILL_5276
timestamp 1745462530
transform 1 0 3552 0 -1 370
box -8 -3 16 105
use FILL  FILL_5277
timestamp 1745462530
transform 1 0 3544 0 -1 370
box -8 -3 16 105
use FILL  FILL_5278
timestamp 1745462530
transform 1 0 3536 0 -1 370
box -8 -3 16 105
use FILL  FILL_5279
timestamp 1745462530
transform 1 0 3416 0 -1 370
box -8 -3 16 105
use FILL  FILL_5280
timestamp 1745462530
transform 1 0 3408 0 -1 370
box -8 -3 16 105
use FILL  FILL_5281
timestamp 1745462530
transform 1 0 3360 0 -1 370
box -8 -3 16 105
use FILL  FILL_5282
timestamp 1745462530
transform 1 0 3352 0 -1 370
box -8 -3 16 105
use FILL  FILL_5283
timestamp 1745462530
transform 1 0 3304 0 -1 370
box -8 -3 16 105
use FILL  FILL_5284
timestamp 1745462530
transform 1 0 3296 0 -1 370
box -8 -3 16 105
use FILL  FILL_5285
timestamp 1745462530
transform 1 0 3248 0 -1 370
box -8 -3 16 105
use FILL  FILL_5286
timestamp 1745462530
transform 1 0 3240 0 -1 370
box -8 -3 16 105
use FILL  FILL_5287
timestamp 1745462530
transform 1 0 3120 0 -1 370
box -8 -3 16 105
use FILL  FILL_5288
timestamp 1745462530
transform 1 0 3016 0 -1 370
box -8 -3 16 105
use FILL  FILL_5289
timestamp 1745462530
transform 1 0 3008 0 -1 370
box -8 -3 16 105
use FILL  FILL_5290
timestamp 1745462530
transform 1 0 2944 0 -1 370
box -8 -3 16 105
use FILL  FILL_5291
timestamp 1745462530
transform 1 0 2936 0 -1 370
box -8 -3 16 105
use FILL  FILL_5292
timestamp 1745462530
transform 1 0 2832 0 -1 370
box -8 -3 16 105
use FILL  FILL_5293
timestamp 1745462530
transform 1 0 2824 0 -1 370
box -8 -3 16 105
use FILL  FILL_5294
timestamp 1745462530
transform 1 0 2704 0 -1 370
box -8 -3 16 105
use FILL  FILL_5295
timestamp 1745462530
transform 1 0 2696 0 -1 370
box -8 -3 16 105
use FILL  FILL_5296
timestamp 1745462530
transform 1 0 2648 0 -1 370
box -8 -3 16 105
use FILL  FILL_5297
timestamp 1745462530
transform 1 0 2640 0 -1 370
box -8 -3 16 105
use FILL  FILL_5298
timestamp 1745462530
transform 1 0 2632 0 -1 370
box -8 -3 16 105
use FILL  FILL_5299
timestamp 1745462530
transform 1 0 2552 0 -1 370
box -8 -3 16 105
use FILL  FILL_5300
timestamp 1745462530
transform 1 0 2544 0 -1 370
box -8 -3 16 105
use FILL  FILL_5301
timestamp 1745462530
transform 1 0 2496 0 -1 370
box -8 -3 16 105
use FILL  FILL_5302
timestamp 1745462530
transform 1 0 2488 0 -1 370
box -8 -3 16 105
use FILL  FILL_5303
timestamp 1745462530
transform 1 0 2480 0 -1 370
box -8 -3 16 105
use FILL  FILL_5304
timestamp 1745462530
transform 1 0 2432 0 -1 370
box -8 -3 16 105
use FILL  FILL_5305
timestamp 1745462530
transform 1 0 2424 0 -1 370
box -8 -3 16 105
use FILL  FILL_5306
timestamp 1745462530
transform 1 0 2400 0 -1 370
box -8 -3 16 105
use FILL  FILL_5307
timestamp 1745462530
transform 1 0 2392 0 -1 370
box -8 -3 16 105
use FILL  FILL_5308
timestamp 1745462530
transform 1 0 2344 0 -1 370
box -8 -3 16 105
use FILL  FILL_5309
timestamp 1745462530
transform 1 0 2336 0 -1 370
box -8 -3 16 105
use FILL  FILL_5310
timestamp 1745462530
transform 1 0 2328 0 -1 370
box -8 -3 16 105
use FILL  FILL_5311
timestamp 1745462530
transform 1 0 2280 0 -1 370
box -8 -3 16 105
use FILL  FILL_5312
timestamp 1745462530
transform 1 0 2272 0 -1 370
box -8 -3 16 105
use FILL  FILL_5313
timestamp 1745462530
transform 1 0 2264 0 -1 370
box -8 -3 16 105
use FILL  FILL_5314
timestamp 1745462530
transform 1 0 2216 0 -1 370
box -8 -3 16 105
use FILL  FILL_5315
timestamp 1745462530
transform 1 0 2208 0 -1 370
box -8 -3 16 105
use FILL  FILL_5316
timestamp 1745462530
transform 1 0 2184 0 -1 370
box -8 -3 16 105
use FILL  FILL_5317
timestamp 1745462530
transform 1 0 2080 0 -1 370
box -8 -3 16 105
use FILL  FILL_5318
timestamp 1745462530
transform 1 0 2072 0 -1 370
box -8 -3 16 105
use FILL  FILL_5319
timestamp 1745462530
transform 1 0 1968 0 -1 370
box -8 -3 16 105
use FILL  FILL_5320
timestamp 1745462530
transform 1 0 1960 0 -1 370
box -8 -3 16 105
use FILL  FILL_5321
timestamp 1745462530
transform 1 0 1936 0 -1 370
box -8 -3 16 105
use FILL  FILL_5322
timestamp 1745462530
transform 1 0 1928 0 -1 370
box -8 -3 16 105
use FILL  FILL_5323
timestamp 1745462530
transform 1 0 1880 0 -1 370
box -8 -3 16 105
use FILL  FILL_5324
timestamp 1745462530
transform 1 0 1872 0 -1 370
box -8 -3 16 105
use FILL  FILL_5325
timestamp 1745462530
transform 1 0 1768 0 -1 370
box -8 -3 16 105
use FILL  FILL_5326
timestamp 1745462530
transform 1 0 1760 0 -1 370
box -8 -3 16 105
use FILL  FILL_5327
timestamp 1745462530
transform 1 0 1752 0 -1 370
box -8 -3 16 105
use FILL  FILL_5328
timestamp 1745462530
transform 1 0 1704 0 -1 370
box -8 -3 16 105
use FILL  FILL_5329
timestamp 1745462530
transform 1 0 1696 0 -1 370
box -8 -3 16 105
use FILL  FILL_5330
timestamp 1745462530
transform 1 0 1672 0 -1 370
box -8 -3 16 105
use FILL  FILL_5331
timestamp 1745462530
transform 1 0 1664 0 -1 370
box -8 -3 16 105
use FILL  FILL_5332
timestamp 1745462530
transform 1 0 1656 0 -1 370
box -8 -3 16 105
use FILL  FILL_5333
timestamp 1745462530
transform 1 0 1608 0 -1 370
box -8 -3 16 105
use FILL  FILL_5334
timestamp 1745462530
transform 1 0 1600 0 -1 370
box -8 -3 16 105
use FILL  FILL_5335
timestamp 1745462530
transform 1 0 1592 0 -1 370
box -8 -3 16 105
use FILL  FILL_5336
timestamp 1745462530
transform 1 0 1584 0 -1 370
box -8 -3 16 105
use FILL  FILL_5337
timestamp 1745462530
transform 1 0 1544 0 -1 370
box -8 -3 16 105
use FILL  FILL_5338
timestamp 1745462530
transform 1 0 1536 0 -1 370
box -8 -3 16 105
use FILL  FILL_5339
timestamp 1745462530
transform 1 0 1528 0 -1 370
box -8 -3 16 105
use FILL  FILL_5340
timestamp 1745462530
transform 1 0 1520 0 -1 370
box -8 -3 16 105
use FILL  FILL_5341
timestamp 1745462530
transform 1 0 1472 0 -1 370
box -8 -3 16 105
use FILL  FILL_5342
timestamp 1745462530
transform 1 0 1464 0 -1 370
box -8 -3 16 105
use FILL  FILL_5343
timestamp 1745462530
transform 1 0 1456 0 -1 370
box -8 -3 16 105
use FILL  FILL_5344
timestamp 1745462530
transform 1 0 1448 0 -1 370
box -8 -3 16 105
use FILL  FILL_5345
timestamp 1745462530
transform 1 0 1400 0 -1 370
box -8 -3 16 105
use FILL  FILL_5346
timestamp 1745462530
transform 1 0 1392 0 -1 370
box -8 -3 16 105
use FILL  FILL_5347
timestamp 1745462530
transform 1 0 1384 0 -1 370
box -8 -3 16 105
use FILL  FILL_5348
timestamp 1745462530
transform 1 0 1360 0 -1 370
box -8 -3 16 105
use FILL  FILL_5349
timestamp 1745462530
transform 1 0 1352 0 -1 370
box -8 -3 16 105
use FILL  FILL_5350
timestamp 1745462530
transform 1 0 1304 0 -1 370
box -8 -3 16 105
use FILL  FILL_5351
timestamp 1745462530
transform 1 0 1296 0 -1 370
box -8 -3 16 105
use FILL  FILL_5352
timestamp 1745462530
transform 1 0 1288 0 -1 370
box -8 -3 16 105
use FILL  FILL_5353
timestamp 1745462530
transform 1 0 1280 0 -1 370
box -8 -3 16 105
use FILL  FILL_5354
timestamp 1745462530
transform 1 0 1176 0 -1 370
box -8 -3 16 105
use FILL  FILL_5355
timestamp 1745462530
transform 1 0 1168 0 -1 370
box -8 -3 16 105
use FILL  FILL_5356
timestamp 1745462530
transform 1 0 1160 0 -1 370
box -8 -3 16 105
use FILL  FILL_5357
timestamp 1745462530
transform 1 0 1152 0 -1 370
box -8 -3 16 105
use FILL  FILL_5358
timestamp 1745462530
transform 1 0 1104 0 -1 370
box -8 -3 16 105
use FILL  FILL_5359
timestamp 1745462530
transform 1 0 1096 0 -1 370
box -8 -3 16 105
use FILL  FILL_5360
timestamp 1745462530
transform 1 0 1072 0 -1 370
box -8 -3 16 105
use FILL  FILL_5361
timestamp 1745462530
transform 1 0 1064 0 -1 370
box -8 -3 16 105
use FILL  FILL_5362
timestamp 1745462530
transform 1 0 960 0 -1 370
box -8 -3 16 105
use FILL  FILL_5363
timestamp 1745462530
transform 1 0 952 0 -1 370
box -8 -3 16 105
use FILL  FILL_5364
timestamp 1745462530
transform 1 0 928 0 -1 370
box -8 -3 16 105
use FILL  FILL_5365
timestamp 1745462530
transform 1 0 880 0 -1 370
box -8 -3 16 105
use FILL  FILL_5366
timestamp 1745462530
transform 1 0 872 0 -1 370
box -8 -3 16 105
use FILL  FILL_5367
timestamp 1745462530
transform 1 0 848 0 -1 370
box -8 -3 16 105
use FILL  FILL_5368
timestamp 1745462530
transform 1 0 800 0 -1 370
box -8 -3 16 105
use FILL  FILL_5369
timestamp 1745462530
transform 1 0 792 0 -1 370
box -8 -3 16 105
use FILL  FILL_5370
timestamp 1745462530
transform 1 0 784 0 -1 370
box -8 -3 16 105
use FILL  FILL_5371
timestamp 1745462530
transform 1 0 744 0 -1 370
box -8 -3 16 105
use FILL  FILL_5372
timestamp 1745462530
transform 1 0 736 0 -1 370
box -8 -3 16 105
use FILL  FILL_5373
timestamp 1745462530
transform 1 0 688 0 -1 370
box -8 -3 16 105
use FILL  FILL_5374
timestamp 1745462530
transform 1 0 680 0 -1 370
box -8 -3 16 105
use FILL  FILL_5375
timestamp 1745462530
transform 1 0 656 0 -1 370
box -8 -3 16 105
use FILL  FILL_5376
timestamp 1745462530
transform 1 0 608 0 -1 370
box -8 -3 16 105
use FILL  FILL_5377
timestamp 1745462530
transform 1 0 600 0 -1 370
box -8 -3 16 105
use FILL  FILL_5378
timestamp 1745462530
transform 1 0 592 0 -1 370
box -8 -3 16 105
use FILL  FILL_5379
timestamp 1745462530
transform 1 0 488 0 -1 370
box -8 -3 16 105
use FILL  FILL_5380
timestamp 1745462530
transform 1 0 480 0 -1 370
box -8 -3 16 105
use FILL  FILL_5381
timestamp 1745462530
transform 1 0 472 0 -1 370
box -8 -3 16 105
use FILL  FILL_5382
timestamp 1745462530
transform 1 0 368 0 -1 370
box -8 -3 16 105
use FILL  FILL_5383
timestamp 1745462530
transform 1 0 360 0 -1 370
box -8 -3 16 105
use FILL  FILL_5384
timestamp 1745462530
transform 1 0 352 0 -1 370
box -8 -3 16 105
use FILL  FILL_5385
timestamp 1745462530
transform 1 0 248 0 -1 370
box -8 -3 16 105
use FILL  FILL_5386
timestamp 1745462530
transform 1 0 240 0 -1 370
box -8 -3 16 105
use FILL  FILL_5387
timestamp 1745462530
transform 1 0 232 0 -1 370
box -8 -3 16 105
use FILL  FILL_5388
timestamp 1745462530
transform 1 0 184 0 -1 370
box -8 -3 16 105
use FILL  FILL_5389
timestamp 1745462530
transform 1 0 176 0 -1 370
box -8 -3 16 105
use FILL  FILL_5390
timestamp 1745462530
transform 1 0 168 0 -1 370
box -8 -3 16 105
use FILL  FILL_5391
timestamp 1745462530
transform 1 0 144 0 -1 370
box -8 -3 16 105
use FILL  FILL_5392
timestamp 1745462530
transform 1 0 136 0 -1 370
box -8 -3 16 105
use FILL  FILL_5393
timestamp 1745462530
transform 1 0 128 0 -1 370
box -8 -3 16 105
use FILL  FILL_5394
timestamp 1745462530
transform 1 0 120 0 -1 370
box -8 -3 16 105
use FILL  FILL_5395
timestamp 1745462530
transform 1 0 112 0 -1 370
box -8 -3 16 105
use FILL  FILL_5396
timestamp 1745462530
transform 1 0 104 0 -1 370
box -8 -3 16 105
use FILL  FILL_5397
timestamp 1745462530
transform 1 0 96 0 -1 370
box -8 -3 16 105
use FILL  FILL_5398
timestamp 1745462530
transform 1 0 88 0 -1 370
box -8 -3 16 105
use FILL  FILL_5399
timestamp 1745462530
transform 1 0 80 0 -1 370
box -8 -3 16 105
use FILL  FILL_5400
timestamp 1745462530
transform 1 0 72 0 -1 370
box -8 -3 16 105
use FILL  FILL_5401
timestamp 1745462530
transform 1 0 4368 0 1 170
box -8 -3 16 105
use FILL  FILL_5402
timestamp 1745462530
transform 1 0 4264 0 1 170
box -8 -3 16 105
use FILL  FILL_5403
timestamp 1745462530
transform 1 0 4256 0 1 170
box -8 -3 16 105
use FILL  FILL_5404
timestamp 1745462530
transform 1 0 4248 0 1 170
box -8 -3 16 105
use FILL  FILL_5405
timestamp 1745462530
transform 1 0 4200 0 1 170
box -8 -3 16 105
use FILL  FILL_5406
timestamp 1745462530
transform 1 0 4192 0 1 170
box -8 -3 16 105
use FILL  FILL_5407
timestamp 1745462530
transform 1 0 4184 0 1 170
box -8 -3 16 105
use FILL  FILL_5408
timestamp 1745462530
transform 1 0 4176 0 1 170
box -8 -3 16 105
use FILL  FILL_5409
timestamp 1745462530
transform 1 0 4128 0 1 170
box -8 -3 16 105
use FILL  FILL_5410
timestamp 1745462530
transform 1 0 4120 0 1 170
box -8 -3 16 105
use FILL  FILL_5411
timestamp 1745462530
transform 1 0 4096 0 1 170
box -8 -3 16 105
use FILL  FILL_5412
timestamp 1745462530
transform 1 0 4072 0 1 170
box -8 -3 16 105
use FILL  FILL_5413
timestamp 1745462530
transform 1 0 4064 0 1 170
box -8 -3 16 105
use FILL  FILL_5414
timestamp 1745462530
transform 1 0 4040 0 1 170
box -8 -3 16 105
use FILL  FILL_5415
timestamp 1745462530
transform 1 0 4032 0 1 170
box -8 -3 16 105
use FILL  FILL_5416
timestamp 1745462530
transform 1 0 4024 0 1 170
box -8 -3 16 105
use FILL  FILL_5417
timestamp 1745462530
transform 1 0 4016 0 1 170
box -8 -3 16 105
use FILL  FILL_5418
timestamp 1745462530
transform 1 0 3968 0 1 170
box -8 -3 16 105
use FILL  FILL_5419
timestamp 1745462530
transform 1 0 3960 0 1 170
box -8 -3 16 105
use FILL  FILL_5420
timestamp 1745462530
transform 1 0 3952 0 1 170
box -8 -3 16 105
use FILL  FILL_5421
timestamp 1745462530
transform 1 0 3928 0 1 170
box -8 -3 16 105
use FILL  FILL_5422
timestamp 1745462530
transform 1 0 3920 0 1 170
box -8 -3 16 105
use FILL  FILL_5423
timestamp 1745462530
transform 1 0 3912 0 1 170
box -8 -3 16 105
use FILL  FILL_5424
timestamp 1745462530
transform 1 0 3864 0 1 170
box -8 -3 16 105
use FILL  FILL_5425
timestamp 1745462530
transform 1 0 3856 0 1 170
box -8 -3 16 105
use FILL  FILL_5426
timestamp 1745462530
transform 1 0 3848 0 1 170
box -8 -3 16 105
use FILL  FILL_5427
timestamp 1745462530
transform 1 0 3840 0 1 170
box -8 -3 16 105
use FILL  FILL_5428
timestamp 1745462530
transform 1 0 3792 0 1 170
box -8 -3 16 105
use FILL  FILL_5429
timestamp 1745462530
transform 1 0 3784 0 1 170
box -8 -3 16 105
use FILL  FILL_5430
timestamp 1745462530
transform 1 0 3776 0 1 170
box -8 -3 16 105
use FILL  FILL_5431
timestamp 1745462530
transform 1 0 3728 0 1 170
box -8 -3 16 105
use FILL  FILL_5432
timestamp 1745462530
transform 1 0 3720 0 1 170
box -8 -3 16 105
use FILL  FILL_5433
timestamp 1745462530
transform 1 0 3696 0 1 170
box -8 -3 16 105
use FILL  FILL_5434
timestamp 1745462530
transform 1 0 3688 0 1 170
box -8 -3 16 105
use FILL  FILL_5435
timestamp 1745462530
transform 1 0 3584 0 1 170
box -8 -3 16 105
use FILL  FILL_5436
timestamp 1745462530
transform 1 0 3576 0 1 170
box -8 -3 16 105
use FILL  FILL_5437
timestamp 1745462530
transform 1 0 3568 0 1 170
box -8 -3 16 105
use FILL  FILL_5438
timestamp 1745462530
transform 1 0 3520 0 1 170
box -8 -3 16 105
use FILL  FILL_5439
timestamp 1745462530
transform 1 0 3512 0 1 170
box -8 -3 16 105
use FILL  FILL_5440
timestamp 1745462530
transform 1 0 3504 0 1 170
box -8 -3 16 105
use FILL  FILL_5441
timestamp 1745462530
transform 1 0 3480 0 1 170
box -8 -3 16 105
use FILL  FILL_5442
timestamp 1745462530
transform 1 0 3472 0 1 170
box -8 -3 16 105
use FILL  FILL_5443
timestamp 1745462530
transform 1 0 3464 0 1 170
box -8 -3 16 105
use FILL  FILL_5444
timestamp 1745462530
transform 1 0 3416 0 1 170
box -8 -3 16 105
use FILL  FILL_5445
timestamp 1745462530
transform 1 0 3408 0 1 170
box -8 -3 16 105
use FILL  FILL_5446
timestamp 1745462530
transform 1 0 3400 0 1 170
box -8 -3 16 105
use FILL  FILL_5447
timestamp 1745462530
transform 1 0 3392 0 1 170
box -8 -3 16 105
use FILL  FILL_5448
timestamp 1745462530
transform 1 0 3352 0 1 170
box -8 -3 16 105
use FILL  FILL_5449
timestamp 1745462530
transform 1 0 3344 0 1 170
box -8 -3 16 105
use FILL  FILL_5450
timestamp 1745462530
transform 1 0 3336 0 1 170
box -8 -3 16 105
use FILL  FILL_5451
timestamp 1745462530
transform 1 0 3288 0 1 170
box -8 -3 16 105
use FILL  FILL_5452
timestamp 1745462530
transform 1 0 3280 0 1 170
box -8 -3 16 105
use FILL  FILL_5453
timestamp 1745462530
transform 1 0 3256 0 1 170
box -8 -3 16 105
use FILL  FILL_5454
timestamp 1745462530
transform 1 0 3248 0 1 170
box -8 -3 16 105
use FILL  FILL_5455
timestamp 1745462530
transform 1 0 3240 0 1 170
box -8 -3 16 105
use FILL  FILL_5456
timestamp 1745462530
transform 1 0 3192 0 1 170
box -8 -3 16 105
use FILL  FILL_5457
timestamp 1745462530
transform 1 0 3184 0 1 170
box -8 -3 16 105
use FILL  FILL_5458
timestamp 1745462530
transform 1 0 3176 0 1 170
box -8 -3 16 105
use FILL  FILL_5459
timestamp 1745462530
transform 1 0 3168 0 1 170
box -8 -3 16 105
use FILL  FILL_5460
timestamp 1745462530
transform 1 0 3144 0 1 170
box -8 -3 16 105
use FILL  FILL_5461
timestamp 1745462530
transform 1 0 3136 0 1 170
box -8 -3 16 105
use FILL  FILL_5462
timestamp 1745462530
transform 1 0 3088 0 1 170
box -8 -3 16 105
use FILL  FILL_5463
timestamp 1745462530
transform 1 0 3080 0 1 170
box -8 -3 16 105
use FILL  FILL_5464
timestamp 1745462530
transform 1 0 3072 0 1 170
box -8 -3 16 105
use FILL  FILL_5465
timestamp 1745462530
transform 1 0 3064 0 1 170
box -8 -3 16 105
use FILL  FILL_5466
timestamp 1745462530
transform 1 0 3016 0 1 170
box -8 -3 16 105
use FILL  FILL_5467
timestamp 1745462530
transform 1 0 3008 0 1 170
box -8 -3 16 105
use FILL  FILL_5468
timestamp 1745462530
transform 1 0 3000 0 1 170
box -8 -3 16 105
use FILL  FILL_5469
timestamp 1745462530
transform 1 0 2992 0 1 170
box -8 -3 16 105
use FILL  FILL_5470
timestamp 1745462530
transform 1 0 2952 0 1 170
box -8 -3 16 105
use FILL  FILL_5471
timestamp 1745462530
transform 1 0 2944 0 1 170
box -8 -3 16 105
use FILL  FILL_5472
timestamp 1745462530
transform 1 0 2936 0 1 170
box -8 -3 16 105
use FILL  FILL_5473
timestamp 1745462530
transform 1 0 2928 0 1 170
box -8 -3 16 105
use FILL  FILL_5474
timestamp 1745462530
transform 1 0 2880 0 1 170
box -8 -3 16 105
use FILL  FILL_5475
timestamp 1745462530
transform 1 0 2872 0 1 170
box -8 -3 16 105
use FILL  FILL_5476
timestamp 1745462530
transform 1 0 2848 0 1 170
box -8 -3 16 105
use FILL  FILL_5477
timestamp 1745462530
transform 1 0 2840 0 1 170
box -8 -3 16 105
use FILL  FILL_5478
timestamp 1745462530
transform 1 0 2792 0 1 170
box -8 -3 16 105
use FILL  FILL_5479
timestamp 1745462530
transform 1 0 2784 0 1 170
box -8 -3 16 105
use FILL  FILL_5480
timestamp 1745462530
transform 1 0 2776 0 1 170
box -8 -3 16 105
use FILL  FILL_5481
timestamp 1745462530
transform 1 0 2768 0 1 170
box -8 -3 16 105
use FILL  FILL_5482
timestamp 1745462530
transform 1 0 2720 0 1 170
box -8 -3 16 105
use FILL  FILL_5483
timestamp 1745462530
transform 1 0 2712 0 1 170
box -8 -3 16 105
use FILL  FILL_5484
timestamp 1745462530
transform 1 0 2704 0 1 170
box -8 -3 16 105
use FILL  FILL_5485
timestamp 1745462530
transform 1 0 2648 0 1 170
box -8 -3 16 105
use FILL  FILL_5486
timestamp 1745462530
transform 1 0 2640 0 1 170
box -8 -3 16 105
use FILL  FILL_5487
timestamp 1745462530
transform 1 0 2592 0 1 170
box -8 -3 16 105
use FILL  FILL_5488
timestamp 1745462530
transform 1 0 2584 0 1 170
box -8 -3 16 105
use FILL  FILL_5489
timestamp 1745462530
transform 1 0 2576 0 1 170
box -8 -3 16 105
use FILL  FILL_5490
timestamp 1745462530
transform 1 0 2552 0 1 170
box -8 -3 16 105
use FILL  FILL_5491
timestamp 1745462530
transform 1 0 2448 0 1 170
box -8 -3 16 105
use FILL  FILL_5492
timestamp 1745462530
transform 1 0 2440 0 1 170
box -8 -3 16 105
use FILL  FILL_5493
timestamp 1745462530
transform 1 0 2336 0 1 170
box -8 -3 16 105
use FILL  FILL_5494
timestamp 1745462530
transform 1 0 2328 0 1 170
box -8 -3 16 105
use FILL  FILL_5495
timestamp 1745462530
transform 1 0 2280 0 1 170
box -8 -3 16 105
use FILL  FILL_5496
timestamp 1745462530
transform 1 0 2272 0 1 170
box -8 -3 16 105
use FILL  FILL_5497
timestamp 1745462530
transform 1 0 2264 0 1 170
box -8 -3 16 105
use FILL  FILL_5498
timestamp 1745462530
transform 1 0 2256 0 1 170
box -8 -3 16 105
use FILL  FILL_5499
timestamp 1745462530
transform 1 0 2208 0 1 170
box -8 -3 16 105
use FILL  FILL_5500
timestamp 1745462530
transform 1 0 2184 0 1 170
box -8 -3 16 105
use FILL  FILL_5501
timestamp 1745462530
transform 1 0 2176 0 1 170
box -8 -3 16 105
use FILL  FILL_5502
timestamp 1745462530
transform 1 0 2072 0 1 170
box -8 -3 16 105
use FILL  FILL_5503
timestamp 1745462530
transform 1 0 2064 0 1 170
box -8 -3 16 105
use FILL  FILL_5504
timestamp 1745462530
transform 1 0 1960 0 1 170
box -8 -3 16 105
use FILL  FILL_5505
timestamp 1745462530
transform 1 0 1936 0 1 170
box -8 -3 16 105
use FILL  FILL_5506
timestamp 1745462530
transform 1 0 1928 0 1 170
box -8 -3 16 105
use FILL  FILL_5507
timestamp 1745462530
transform 1 0 1920 0 1 170
box -8 -3 16 105
use FILL  FILL_5508
timestamp 1745462530
transform 1 0 1872 0 1 170
box -8 -3 16 105
use FILL  FILL_5509
timestamp 1745462530
transform 1 0 1864 0 1 170
box -8 -3 16 105
use FILL  FILL_5510
timestamp 1745462530
transform 1 0 1856 0 1 170
box -8 -3 16 105
use FILL  FILL_5511
timestamp 1745462530
transform 1 0 1832 0 1 170
box -8 -3 16 105
use FILL  FILL_5512
timestamp 1745462530
transform 1 0 1824 0 1 170
box -8 -3 16 105
use FILL  FILL_5513
timestamp 1745462530
transform 1 0 1776 0 1 170
box -8 -3 16 105
use FILL  FILL_5514
timestamp 1745462530
transform 1 0 1768 0 1 170
box -8 -3 16 105
use FILL  FILL_5515
timestamp 1745462530
transform 1 0 1760 0 1 170
box -8 -3 16 105
use FILL  FILL_5516
timestamp 1745462530
transform 1 0 1736 0 1 170
box -8 -3 16 105
use FILL  FILL_5517
timestamp 1745462530
transform 1 0 1728 0 1 170
box -8 -3 16 105
use FILL  FILL_5518
timestamp 1745462530
transform 1 0 1720 0 1 170
box -8 -3 16 105
use FILL  FILL_5519
timestamp 1745462530
transform 1 0 1672 0 1 170
box -8 -3 16 105
use FILL  FILL_5520
timestamp 1745462530
transform 1 0 1664 0 1 170
box -8 -3 16 105
use FILL  FILL_5521
timestamp 1745462530
transform 1 0 1656 0 1 170
box -8 -3 16 105
use FILL  FILL_5522
timestamp 1745462530
transform 1 0 1552 0 1 170
box -8 -3 16 105
use FILL  FILL_5523
timestamp 1745462530
transform 1 0 1544 0 1 170
box -8 -3 16 105
use FILL  FILL_5524
timestamp 1745462530
transform 1 0 1504 0 1 170
box -8 -3 16 105
use FILL  FILL_5525
timestamp 1745462530
transform 1 0 1496 0 1 170
box -8 -3 16 105
use FILL  FILL_5526
timestamp 1745462530
transform 1 0 1488 0 1 170
box -8 -3 16 105
use FILL  FILL_5527
timestamp 1745462530
transform 1 0 1480 0 1 170
box -8 -3 16 105
use FILL  FILL_5528
timestamp 1745462530
transform 1 0 1432 0 1 170
box -8 -3 16 105
use FILL  FILL_5529
timestamp 1745462530
transform 1 0 1424 0 1 170
box -8 -3 16 105
use FILL  FILL_5530
timestamp 1745462530
transform 1 0 1400 0 1 170
box -8 -3 16 105
use FILL  FILL_5531
timestamp 1745462530
transform 1 0 1392 0 1 170
box -8 -3 16 105
use FILL  FILL_5532
timestamp 1745462530
transform 1 0 1344 0 1 170
box -8 -3 16 105
use FILL  FILL_5533
timestamp 1745462530
transform 1 0 1336 0 1 170
box -8 -3 16 105
use FILL  FILL_5534
timestamp 1745462530
transform 1 0 1232 0 1 170
box -8 -3 16 105
use FILL  FILL_5535
timestamp 1745462530
transform 1 0 1208 0 1 170
box -8 -3 16 105
use FILL  FILL_5536
timestamp 1745462530
transform 1 0 1200 0 1 170
box -8 -3 16 105
use FILL  FILL_5537
timestamp 1745462530
transform 1 0 1192 0 1 170
box -8 -3 16 105
use FILL  FILL_5538
timestamp 1745462530
transform 1 0 1144 0 1 170
box -8 -3 16 105
use FILL  FILL_5539
timestamp 1745462530
transform 1 0 1136 0 1 170
box -8 -3 16 105
use FILL  FILL_5540
timestamp 1745462530
transform 1 0 1088 0 1 170
box -8 -3 16 105
use FILL  FILL_5541
timestamp 1745462530
transform 1 0 1080 0 1 170
box -8 -3 16 105
use FILL  FILL_5542
timestamp 1745462530
transform 1 0 960 0 1 170
box -8 -3 16 105
use FILL  FILL_5543
timestamp 1745462530
transform 1 0 952 0 1 170
box -8 -3 16 105
use FILL  FILL_5544
timestamp 1745462530
transform 1 0 944 0 1 170
box -8 -3 16 105
use FILL  FILL_5545
timestamp 1745462530
transform 1 0 880 0 1 170
box -8 -3 16 105
use FILL  FILL_5546
timestamp 1745462530
transform 1 0 816 0 1 170
box -8 -3 16 105
use FILL  FILL_5547
timestamp 1745462530
transform 1 0 808 0 1 170
box -8 -3 16 105
use FILL  FILL_5548
timestamp 1745462530
transform 1 0 704 0 1 170
box -8 -3 16 105
use FILL  FILL_5549
timestamp 1745462530
transform 1 0 680 0 1 170
box -8 -3 16 105
use FILL  FILL_5550
timestamp 1745462530
transform 1 0 576 0 1 170
box -8 -3 16 105
use FILL  FILL_5551
timestamp 1745462530
transform 1 0 568 0 1 170
box -8 -3 16 105
use FILL  FILL_5552
timestamp 1745462530
transform 1 0 544 0 1 170
box -8 -3 16 105
use FILL  FILL_5553
timestamp 1745462530
transform 1 0 440 0 1 170
box -8 -3 16 105
use FILL  FILL_5554
timestamp 1745462530
transform 1 0 432 0 1 170
box -8 -3 16 105
use FILL  FILL_5555
timestamp 1745462530
transform 1 0 424 0 1 170
box -8 -3 16 105
use FILL  FILL_5556
timestamp 1745462530
transform 1 0 376 0 1 170
box -8 -3 16 105
use FILL  FILL_5557
timestamp 1745462530
transform 1 0 368 0 1 170
box -8 -3 16 105
use FILL  FILL_5558
timestamp 1745462530
transform 1 0 304 0 1 170
box -8 -3 16 105
use FILL  FILL_5559
timestamp 1745462530
transform 1 0 296 0 1 170
box -8 -3 16 105
use FILL  FILL_5560
timestamp 1745462530
transform 1 0 288 0 1 170
box -8 -3 16 105
use FILL  FILL_5561
timestamp 1745462530
transform 1 0 280 0 1 170
box -8 -3 16 105
use FILL  FILL_5562
timestamp 1745462530
transform 1 0 232 0 1 170
box -8 -3 16 105
use FILL  FILL_5563
timestamp 1745462530
transform 1 0 224 0 1 170
box -8 -3 16 105
use FILL  FILL_5564
timestamp 1745462530
transform 1 0 200 0 1 170
box -8 -3 16 105
use FILL  FILL_5565
timestamp 1745462530
transform 1 0 192 0 1 170
box -8 -3 16 105
use FILL  FILL_5566
timestamp 1745462530
transform 1 0 184 0 1 170
box -8 -3 16 105
use FILL  FILL_5567
timestamp 1745462530
transform 1 0 80 0 1 170
box -8 -3 16 105
use FILL  FILL_5568
timestamp 1745462530
transform 1 0 72 0 1 170
box -8 -3 16 105
use FILL  FILL_5569
timestamp 1745462530
transform 1 0 4368 0 -1 170
box -8 -3 16 105
use FILL  FILL_5570
timestamp 1745462530
transform 1 0 4360 0 -1 170
box -8 -3 16 105
use FILL  FILL_5571
timestamp 1745462530
transform 1 0 4256 0 -1 170
box -8 -3 16 105
use FILL  FILL_5572
timestamp 1745462530
transform 1 0 4232 0 -1 170
box -8 -3 16 105
use FILL  FILL_5573
timestamp 1745462530
transform 1 0 4224 0 -1 170
box -8 -3 16 105
use FILL  FILL_5574
timestamp 1745462530
transform 1 0 4120 0 -1 170
box -8 -3 16 105
use FILL  FILL_5575
timestamp 1745462530
transform 1 0 4016 0 -1 170
box -8 -3 16 105
use FILL  FILL_5576
timestamp 1745462530
transform 1 0 4008 0 -1 170
box -8 -3 16 105
use FILL  FILL_5577
timestamp 1745462530
transform 1 0 4000 0 -1 170
box -8 -3 16 105
use FILL  FILL_5578
timestamp 1745462530
transform 1 0 3896 0 -1 170
box -8 -3 16 105
use FILL  FILL_5579
timestamp 1745462530
transform 1 0 3888 0 -1 170
box -8 -3 16 105
use FILL  FILL_5580
timestamp 1745462530
transform 1 0 3784 0 -1 170
box -8 -3 16 105
use FILL  FILL_5581
timestamp 1745462530
transform 1 0 3776 0 -1 170
box -8 -3 16 105
use FILL  FILL_5582
timestamp 1745462530
transform 1 0 3768 0 -1 170
box -8 -3 16 105
use FILL  FILL_5583
timestamp 1745462530
transform 1 0 3664 0 -1 170
box -8 -3 16 105
use FILL  FILL_5584
timestamp 1745462530
transform 1 0 3656 0 -1 170
box -8 -3 16 105
use FILL  FILL_5585
timestamp 1745462530
transform 1 0 3552 0 -1 170
box -8 -3 16 105
use FILL  FILL_5586
timestamp 1745462530
transform 1 0 3544 0 -1 170
box -8 -3 16 105
use FILL  FILL_5587
timestamp 1745462530
transform 1 0 3440 0 -1 170
box -8 -3 16 105
use FILL  FILL_5588
timestamp 1745462530
transform 1 0 3432 0 -1 170
box -8 -3 16 105
use FILL  FILL_5589
timestamp 1745462530
transform 1 0 3328 0 -1 170
box -8 -3 16 105
use FILL  FILL_5590
timestamp 1745462530
transform 1 0 3320 0 -1 170
box -8 -3 16 105
use FILL  FILL_5591
timestamp 1745462530
transform 1 0 3216 0 -1 170
box -8 -3 16 105
use FILL  FILL_5592
timestamp 1745462530
transform 1 0 3208 0 -1 170
box -8 -3 16 105
use FILL  FILL_5593
timestamp 1745462530
transform 1 0 3104 0 -1 170
box -8 -3 16 105
use FILL  FILL_5594
timestamp 1745462530
transform 1 0 3096 0 -1 170
box -8 -3 16 105
use FILL  FILL_5595
timestamp 1745462530
transform 1 0 2992 0 -1 170
box -8 -3 16 105
use FILL  FILL_5596
timestamp 1745462530
transform 1 0 2888 0 -1 170
box -8 -3 16 105
use FILL  FILL_5597
timestamp 1745462530
transform 1 0 2880 0 -1 170
box -8 -3 16 105
use FILL  FILL_5598
timestamp 1745462530
transform 1 0 2776 0 -1 170
box -8 -3 16 105
use FILL  FILL_5599
timestamp 1745462530
transform 1 0 2672 0 -1 170
box -8 -3 16 105
use FILL  FILL_5600
timestamp 1745462530
transform 1 0 2664 0 -1 170
box -8 -3 16 105
use FILL  FILL_5601
timestamp 1745462530
transform 1 0 2640 0 -1 170
box -8 -3 16 105
use FILL  FILL_5602
timestamp 1745462530
transform 1 0 2536 0 -1 170
box -8 -3 16 105
use FILL  FILL_5603
timestamp 1745462530
transform 1 0 2528 0 -1 170
box -8 -3 16 105
use FILL  FILL_5604
timestamp 1745462530
transform 1 0 2480 0 -1 170
box -8 -3 16 105
use FILL  FILL_5605
timestamp 1745462530
transform 1 0 2472 0 -1 170
box -8 -3 16 105
use FILL  FILL_5606
timestamp 1745462530
transform 1 0 2448 0 -1 170
box -8 -3 16 105
use FILL  FILL_5607
timestamp 1745462530
transform 1 0 2440 0 -1 170
box -8 -3 16 105
use FILL  FILL_5608
timestamp 1745462530
transform 1 0 2336 0 -1 170
box -8 -3 16 105
use FILL  FILL_5609
timestamp 1745462530
transform 1 0 2312 0 -1 170
box -8 -3 16 105
use FILL  FILL_5610
timestamp 1745462530
transform 1 0 2208 0 -1 170
box -8 -3 16 105
use FILL  FILL_5611
timestamp 1745462530
transform 1 0 2184 0 -1 170
box -8 -3 16 105
use FILL  FILL_5612
timestamp 1745462530
transform 1 0 2176 0 -1 170
box -8 -3 16 105
use FILL  FILL_5613
timestamp 1745462530
transform 1 0 2072 0 -1 170
box -8 -3 16 105
use FILL  FILL_5614
timestamp 1745462530
transform 1 0 2064 0 -1 170
box -8 -3 16 105
use FILL  FILL_5615
timestamp 1745462530
transform 1 0 1960 0 -1 170
box -8 -3 16 105
use FILL  FILL_5616
timestamp 1745462530
transform 1 0 1936 0 -1 170
box -8 -3 16 105
use FILL  FILL_5617
timestamp 1745462530
transform 1 0 1928 0 -1 170
box -8 -3 16 105
use FILL  FILL_5618
timestamp 1745462530
transform 1 0 1880 0 -1 170
box -8 -3 16 105
use FILL  FILL_5619
timestamp 1745462530
transform 1 0 1872 0 -1 170
box -8 -3 16 105
use FILL  FILL_5620
timestamp 1745462530
transform 1 0 1768 0 -1 170
box -8 -3 16 105
use FILL  FILL_5621
timestamp 1745462530
transform 1 0 1760 0 -1 170
box -8 -3 16 105
use FILL  FILL_5622
timestamp 1745462530
transform 1 0 1656 0 -1 170
box -8 -3 16 105
use FILL  FILL_5623
timestamp 1745462530
transform 1 0 1552 0 -1 170
box -8 -3 16 105
use FILL  FILL_5624
timestamp 1745462530
transform 1 0 1528 0 -1 170
box -8 -3 16 105
use FILL  FILL_5625
timestamp 1745462530
transform 1 0 1520 0 -1 170
box -8 -3 16 105
use FILL  FILL_5626
timestamp 1745462530
transform 1 0 1472 0 -1 170
box -8 -3 16 105
use FILL  FILL_5627
timestamp 1745462530
transform 1 0 1464 0 -1 170
box -8 -3 16 105
use FILL  FILL_5628
timestamp 1745462530
transform 1 0 1360 0 -1 170
box -8 -3 16 105
use FILL  FILL_5629
timestamp 1745462530
transform 1 0 1352 0 -1 170
box -8 -3 16 105
use FILL  FILL_5630
timestamp 1745462530
transform 1 0 1344 0 -1 170
box -8 -3 16 105
use FILL  FILL_5631
timestamp 1745462530
transform 1 0 1296 0 -1 170
box -8 -3 16 105
use FILL  FILL_5632
timestamp 1745462530
transform 1 0 1288 0 -1 170
box -8 -3 16 105
use FILL  FILL_5633
timestamp 1745462530
transform 1 0 1264 0 -1 170
box -8 -3 16 105
use FILL  FILL_5634
timestamp 1745462530
transform 1 0 1160 0 -1 170
box -8 -3 16 105
use FILL  FILL_5635
timestamp 1745462530
transform 1 0 1152 0 -1 170
box -8 -3 16 105
use FILL  FILL_5636
timestamp 1745462530
transform 1 0 1128 0 -1 170
box -8 -3 16 105
use FILL  FILL_5637
timestamp 1745462530
transform 1 0 1120 0 -1 170
box -8 -3 16 105
use FILL  FILL_5638
timestamp 1745462530
transform 1 0 1016 0 -1 170
box -8 -3 16 105
use FILL  FILL_5639
timestamp 1745462530
transform 1 0 1008 0 -1 170
box -8 -3 16 105
use FILL  FILL_5640
timestamp 1745462530
transform 1 0 904 0 -1 170
box -8 -3 16 105
use FILL  FILL_5641
timestamp 1745462530
transform 1 0 896 0 -1 170
box -8 -3 16 105
use FILL  FILL_5642
timestamp 1745462530
transform 1 0 792 0 -1 170
box -8 -3 16 105
use FILL  FILL_5643
timestamp 1745462530
transform 1 0 784 0 -1 170
box -8 -3 16 105
use FILL  FILL_5644
timestamp 1745462530
transform 1 0 776 0 -1 170
box -8 -3 16 105
use FILL  FILL_5645
timestamp 1745462530
transform 1 0 672 0 -1 170
box -8 -3 16 105
use FILL  FILL_5646
timestamp 1745462530
transform 1 0 664 0 -1 170
box -8 -3 16 105
use FILL  FILL_5647
timestamp 1745462530
transform 1 0 600 0 -1 170
box -8 -3 16 105
use FILL  FILL_5648
timestamp 1745462530
transform 1 0 592 0 -1 170
box -8 -3 16 105
use FILL  FILL_5649
timestamp 1745462530
transform 1 0 584 0 -1 170
box -8 -3 16 105
use FILL  FILL_5650
timestamp 1745462530
transform 1 0 520 0 -1 170
box -8 -3 16 105
use FILL  FILL_5651
timestamp 1745462530
transform 1 0 512 0 -1 170
box -8 -3 16 105
use FILL  FILL_5652
timestamp 1745462530
transform 1 0 408 0 -1 170
box -8 -3 16 105
use FILL  FILL_5653
timestamp 1745462530
transform 1 0 400 0 -1 170
box -8 -3 16 105
use FILL  FILL_5654
timestamp 1745462530
transform 1 0 392 0 -1 170
box -8 -3 16 105
use FILL  FILL_5655
timestamp 1745462530
transform 1 0 288 0 -1 170
box -8 -3 16 105
use FILL  FILL_5656
timestamp 1745462530
transform 1 0 280 0 -1 170
box -8 -3 16 105
use FILL  FILL_5657
timestamp 1745462530
transform 1 0 256 0 -1 170
box -8 -3 16 105
use FILL  FILL_5658
timestamp 1745462530
transform 1 0 152 0 -1 170
box -8 -3 16 105
use FILL  FILL_5659
timestamp 1745462530
transform 1 0 144 0 -1 170
box -8 -3 16 105
use FILL  FILL_5660
timestamp 1745462530
transform 1 0 136 0 -1 170
box -8 -3 16 105
use FILL  FILL_5661
timestamp 1745462530
transform 1 0 128 0 -1 170
box -8 -3 16 105
use FILL  FILL_5662
timestamp 1745462530
transform 1 0 120 0 -1 170
box -8 -3 16 105
use FILL  FILL_5663
timestamp 1745462530
transform 1 0 112 0 -1 170
box -8 -3 16 105
use FILL  FILL_5664
timestamp 1745462530
transform 1 0 104 0 -1 170
box -8 -3 16 105
use FILL  FILL_5665
timestamp 1745462530
transform 1 0 96 0 -1 170
box -8 -3 16 105
use FILL  FILL_5666
timestamp 1745462530
transform 1 0 88 0 -1 170
box -8 -3 16 105
use FILL  FILL_5667
timestamp 1745462530
transform 1 0 80 0 -1 170
box -8 -3 16 105
use FILL  FILL_5668
timestamp 1745462530
transform 1 0 72 0 -1 170
box -8 -3 16 105
use HAX1  HAX1_0
timestamp 1745462530
transform 1 0 152 0 1 2970
box -5 -3 84 105
use HAX1  HAX1_1
timestamp 1745462530
transform 1 0 288 0 -1 3170
box -5 -3 84 105
use HAX1  HAX1_2
timestamp 1745462530
transform 1 0 392 0 -1 3170
box -5 -3 84 105
use HAX1  HAX1_3
timestamp 1745462530
transform 1 0 480 0 -1 3170
box -5 -3 84 105
use INVX2  INVX2_0
timestamp 1745462530
transform 1 0 288 0 -1 3570
box -9 -3 26 105
use INVX2  INVX2_1
timestamp 1745462530
transform 1 0 160 0 -1 3570
box -9 -3 26 105
use INVX2  INVX2_2
timestamp 1745462530
transform 1 0 416 0 -1 3570
box -9 -3 26 105
use INVX2  INVX2_3
timestamp 1745462530
transform 1 0 272 0 1 3370
box -9 -3 26 105
use INVX2  INVX2_4
timestamp 1745462530
transform 1 0 352 0 1 3570
box -9 -3 26 105
use INVX2  INVX2_5
timestamp 1745462530
transform 1 0 216 0 1 3570
box -9 -3 26 105
use INVX2  INVX2_6
timestamp 1745462530
transform 1 0 216 0 1 3370
box -9 -3 26 105
use INVX2  INVX2_7
timestamp 1745462530
transform 1 0 80 0 -1 3570
box -9 -3 26 105
use INVX2  INVX2_8
timestamp 1745462530
transform 1 0 1160 0 -1 3570
box -9 -3 26 105
use INVX2  INVX2_9
timestamp 1745462530
transform 1 0 2192 0 -1 3370
box -9 -3 26 105
use INVX2  INVX2_10
timestamp 1745462530
transform 1 0 2080 0 1 3370
box -9 -3 26 105
use INVX2  INVX2_11
timestamp 1745462530
transform 1 0 2048 0 1 3370
box -9 -3 26 105
use INVX2  INVX2_12
timestamp 1745462530
transform 1 0 3048 0 -1 3370
box -9 -3 26 105
use INVX2  INVX2_13
timestamp 1745462530
transform 1 0 3024 0 1 3170
box -9 -3 26 105
use INVX2  INVX2_14
timestamp 1745462530
transform 1 0 2968 0 1 3170
box -9 -3 26 105
use INVX2  INVX2_15
timestamp 1745462530
transform 1 0 1504 0 1 2970
box -9 -3 26 105
use INVX2  INVX2_16
timestamp 1745462530
transform 1 0 1576 0 -1 3370
box -9 -3 26 105
use INVX2  INVX2_17
timestamp 1745462530
transform 1 0 1632 0 -1 3570
box -9 -3 26 105
use INVX2  INVX2_18
timestamp 1745462530
transform 1 0 728 0 1 3170
box -9 -3 26 105
use INVX2  INVX2_19
timestamp 1745462530
transform 1 0 2192 0 1 2170
box -9 -3 26 105
use INVX2  INVX2_20
timestamp 1745462530
transform 1 0 2328 0 -1 2770
box -9 -3 26 105
use INVX2  INVX2_21
timestamp 1745462530
transform 1 0 2384 0 -1 2570
box -9 -3 26 105
use INVX2  INVX2_22
timestamp 1745462530
transform 1 0 2224 0 -1 2370
box -9 -3 26 105
use INVX2  INVX2_23
timestamp 1745462530
transform 1 0 2216 0 1 2170
box -9 -3 26 105
use INVX2  INVX2_24
timestamp 1745462530
transform 1 0 2560 0 1 2370
box -9 -3 26 105
use INVX2  INVX2_25
timestamp 1745462530
transform 1 0 2344 0 -1 2770
box -9 -3 26 105
use INVX2  INVX2_26
timestamp 1745462530
transform 1 0 2544 0 1 2370
box -9 -3 26 105
use INVX2  INVX2_27
timestamp 1745462530
transform 1 0 2208 0 1 2370
box -9 -3 26 105
use INVX2  INVX2_28
timestamp 1745462530
transform 1 0 2640 0 -1 2570
box -9 -3 26 105
use INVX2  INVX2_29
timestamp 1745462530
transform 1 0 1056 0 1 2370
box -9 -3 26 105
use INVX2  INVX2_30
timestamp 1745462530
transform 1 0 2384 0 1 2570
box -9 -3 26 105
use INVX2  INVX2_31
timestamp 1745462530
transform 1 0 2208 0 -1 2370
box -9 -3 26 105
use INVX2  INVX2_32
timestamp 1745462530
transform 1 0 2312 0 1 1770
box -9 -3 26 105
use INVX2  INVX2_33
timestamp 1745462530
transform 1 0 960 0 1 770
box -9 -3 26 105
use INVX2  INVX2_34
timestamp 1745462530
transform 1 0 1552 0 -1 770
box -9 -3 26 105
use INVX2  INVX2_35
timestamp 1745462530
transform 1 0 3248 0 -1 1370
box -9 -3 26 105
use INVX2  INVX2_36
timestamp 1745462530
transform 1 0 2608 0 -1 2370
box -9 -3 26 105
use INVX2  INVX2_37
timestamp 1745462530
transform 1 0 2232 0 1 2170
box -9 -3 26 105
use INVX2  INVX2_38
timestamp 1745462530
transform 1 0 3248 0 -1 770
box -9 -3 26 105
use INVX2  INVX2_39
timestamp 1745462530
transform 1 0 1008 0 1 2370
box -9 -3 26 105
use INVX2  INVX2_40
timestamp 1745462530
transform 1 0 2680 0 -1 770
box -9 -3 26 105
use INVX2  INVX2_41
timestamp 1745462530
transform 1 0 2120 0 1 2370
box -9 -3 26 105
use INVX2  INVX2_42
timestamp 1745462530
transform 1 0 2144 0 -1 1970
box -9 -3 26 105
use INVX2  INVX2_43
timestamp 1745462530
transform 1 0 2128 0 -1 1970
box -9 -3 26 105
use INVX2  INVX2_44
timestamp 1745462530
transform 1 0 1792 0 1 1970
box -9 -3 26 105
use INVX2  INVX2_45
timestamp 1745462530
transform 1 0 1424 0 -1 2570
box -9 -3 26 105
use INVX2  INVX2_46
timestamp 1745462530
transform 1 0 1480 0 -1 1970
box -9 -3 26 105
use INVX2  INVX2_47
timestamp 1745462530
transform 1 0 336 0 1 2770
box -9 -3 26 105
use INVX2  INVX2_48
timestamp 1745462530
transform 1 0 504 0 1 2770
box -9 -3 26 105
use INVX2  INVX2_49
timestamp 1745462530
transform 1 0 264 0 1 2770
box -9 -3 26 105
use INVX2  INVX2_50
timestamp 1745462530
transform 1 0 920 0 1 2770
box -9 -3 26 105
use INVX2  INVX2_51
timestamp 1745462530
transform 1 0 184 0 1 2370
box -9 -3 26 105
use INVX2  INVX2_52
timestamp 1745462530
transform 1 0 208 0 -1 970
box -9 -3 26 105
use INVX2  INVX2_53
timestamp 1745462530
transform 1 0 208 0 1 170
box -9 -3 26 105
use INVX2  INVX2_54
timestamp 1745462530
transform 1 0 256 0 1 370
box -9 -3 26 105
use INVX2  INVX2_55
timestamp 1745462530
transform 1 0 688 0 1 170
box -9 -3 26 105
use INVX2  INVX2_56
timestamp 1745462530
transform 1 0 1456 0 1 370
box -9 -3 26 105
use INVX2  INVX2_57
timestamp 1745462530
transform 1 0 1528 0 1 170
box -9 -3 26 105
use INVX2  INVX2_58
timestamp 1745462530
transform 1 0 1616 0 -1 770
box -9 -3 26 105
use INVX2  INVX2_59
timestamp 1745462530
transform 1 0 1552 0 -1 370
box -9 -3 26 105
use INVX2  INVX2_60
timestamp 1745462530
transform 1 0 2704 0 -1 770
box -9 -3 26 105
use INVX2  INVX2_61
timestamp 1745462530
transform 1 0 2672 0 1 170
box -9 -3 26 105
use INVX2  INVX2_62
timestamp 1745462530
transform 1 0 2688 0 1 370
box -9 -3 26 105
use INVX2  INVX2_63
timestamp 1745462530
transform 1 0 2656 0 1 170
box -9 -3 26 105
use INVX2  INVX2_64
timestamp 1745462530
transform 1 0 3808 0 -1 370
box -9 -3 26 105
use INVX2  INVX2_65
timestamp 1745462530
transform 1 0 4080 0 1 170
box -9 -3 26 105
use INVX2  INVX2_66
timestamp 1745462530
transform 1 0 3704 0 -1 370
box -9 -3 26 105
use INVX2  INVX2_67
timestamp 1745462530
transform 1 0 4264 0 -1 370
box -9 -3 26 105
use INVX2  INVX2_68
timestamp 1745462530
transform 1 0 3688 0 -1 1570
box -9 -3 26 105
use INVX2  INVX2_69
timestamp 1745462530
transform 1 0 4184 0 1 1770
box -9 -3 26 105
use INVX2  INVX2_70
timestamp 1745462530
transform 1 0 3840 0 -1 1770
box -9 -3 26 105
use INVX2  INVX2_71
timestamp 1745462530
transform 1 0 4168 0 1 1770
box -9 -3 26 105
use INVX2  INVX2_72
timestamp 1745462530
transform 1 0 4152 0 -1 2370
box -9 -3 26 105
use INVX2  INVX2_73
timestamp 1745462530
transform 1 0 3696 0 -1 2970
box -9 -3 26 105
use INVX2  INVX2_74
timestamp 1745462530
transform 1 0 1640 0 1 2770
box -9 -3 26 105
use INVX2  INVX2_75
timestamp 1745462530
transform 1 0 1640 0 1 2170
box -9 -3 26 105
use INVX2  INVX2_76
timestamp 1745462530
transform 1 0 1672 0 1 2570
box -9 -3 26 105
use INVX2  INVX2_77
timestamp 1745462530
transform 1 0 248 0 -1 2170
box -9 -3 26 105
use INVX2  INVX2_78
timestamp 1745462530
transform 1 0 224 0 1 1770
box -9 -3 26 105
use INVX2  INVX2_79
timestamp 1745462530
transform 1 0 592 0 -1 1770
box -9 -3 26 105
use INVX2  INVX2_80
timestamp 1745462530
transform 1 0 392 0 1 1570
box -9 -3 26 105
use INVX2  INVX2_81
timestamp 1745462530
transform 1 0 856 0 -1 370
box -9 -3 26 105
use INVX2  INVX2_82
timestamp 1745462530
transform 1 0 248 0 1 1170
box -9 -3 26 105
use INVX2  INVX2_83
timestamp 1745462530
transform 1 0 800 0 1 1370
box -9 -3 26 105
use INVX2  INVX2_84
timestamp 1745462530
transform 1 0 1512 0 1 170
box -9 -3 26 105
use INVX2  INVX2_85
timestamp 1745462530
transform 1 0 1944 0 -1 970
box -9 -3 26 105
use INVX2  INVX2_86
timestamp 1745462530
transform 1 0 1624 0 -1 1370
box -9 -3 26 105
use INVX2  INVX2_87
timestamp 1745462530
transform 1 0 1600 0 1 1370
box -9 -3 26 105
use INVX2  INVX2_88
timestamp 1745462530
transform 1 0 2560 0 -1 370
box -9 -3 26 105
use INVX2  INVX2_89
timestamp 1745462530
transform 1 0 2760 0 1 970
box -9 -3 26 105
use INVX2  INVX2_90
timestamp 1745462530
transform 1 0 2640 0 -1 1170
box -9 -3 26 105
use INVX2  INVX2_91
timestamp 1745462530
transform 1 0 2688 0 -1 1370
box -9 -3 26 105
use INVX2  INVX2_92
timestamp 1745462530
transform 1 0 3360 0 1 170
box -9 -3 26 105
use INVX2  INVX2_93
timestamp 1745462530
transform 1 0 4192 0 -1 970
box -9 -3 26 105
use INVX2  INVX2_94
timestamp 1745462530
transform 1 0 4104 0 1 970
box -9 -3 26 105
use INVX2  INVX2_95
timestamp 1745462530
transform 1 0 3816 0 1 1170
box -9 -3 26 105
use INVX2  INVX2_96
timestamp 1745462530
transform 1 0 4136 0 -1 1770
box -9 -3 26 105
use INVX2  INVX2_97
timestamp 1745462530
transform 1 0 3736 0 1 2170
box -9 -3 26 105
use INVX2  INVX2_98
timestamp 1745462530
transform 1 0 2976 0 -1 1970
box -9 -3 26 105
use INVX2  INVX2_99
timestamp 1745462530
transform 1 0 2696 0 -1 2170
box -9 -3 26 105
use INVX2  INVX2_100
timestamp 1745462530
transform 1 0 3736 0 -1 2770
box -9 -3 26 105
use INVX2  INVX2_101
timestamp 1745462530
transform 1 0 3888 0 1 2970
box -9 -3 26 105
use INVX2  INVX2_102
timestamp 1745462530
transform 1 0 4008 0 1 2770
box -9 -3 26 105
use INVX2  INVX2_103
timestamp 1745462530
transform 1 0 4200 0 -1 2970
box -9 -3 26 105
use INVX2  INVX2_104
timestamp 1745462530
transform 1 0 3944 0 1 2370
box -9 -3 26 105
use INVX2  INVX2_105
timestamp 1745462530
transform 1 0 2832 0 1 2570
box -9 -3 26 105
use INVX2  INVX2_106
timestamp 1745462530
transform 1 0 2824 0 -1 2770
box -9 -3 26 105
use INVX2  INVX2_107
timestamp 1745462530
transform 1 0 1064 0 1 3170
box -9 -3 26 105
use INVX2  INVX2_108
timestamp 1745462530
transform 1 0 1064 0 -1 3570
box -9 -3 26 105
use INVX2  INVX2_109
timestamp 1745462530
transform 1 0 1352 0 -1 3170
box -9 -3 26 105
use INVX2  INVX2_110
timestamp 1745462530
transform 1 0 816 0 1 3370
box -9 -3 26 105
use INVX2  INVX2_111
timestamp 1745462530
transform 1 0 1128 0 1 3570
box -9 -3 26 105
use INVX2  INVX2_112
timestamp 1745462530
transform 1 0 1024 0 1 3570
box -9 -3 26 105
use INVX2  INVX2_113
timestamp 1745462530
transform 1 0 856 0 1 3570
box -9 -3 26 105
use INVX2  INVX2_114
timestamp 1745462530
transform 1 0 792 0 -1 3570
box -9 -3 26 105
use INVX2  INVX2_115
timestamp 1745462530
transform 1 0 952 0 -1 3370
box -9 -3 26 105
use INVX2  INVX2_116
timestamp 1745462530
transform 1 0 1504 0 1 3170
box -9 -3 26 105
use INVX2  INVX2_117
timestamp 1745462530
transform 1 0 1584 0 1 3370
box -9 -3 26 105
use INVX2  INVX2_118
timestamp 1745462530
transform 1 0 1280 0 1 3170
box -9 -3 26 105
use INVX2  INVX2_119
timestamp 1745462530
transform 1 0 1592 0 -1 3370
box -9 -3 26 105
use INVX2  INVX2_120
timestamp 1745462530
transform 1 0 1712 0 -1 3170
box -9 -3 26 105
use INVX2  INVX2_121
timestamp 1745462530
transform 1 0 1568 0 1 2970
box -9 -3 26 105
use INVX2  INVX2_122
timestamp 1745462530
transform 1 0 1768 0 1 3370
box -9 -3 26 105
use INVX2  INVX2_123
timestamp 1745462530
transform 1 0 1768 0 -1 3770
box -9 -3 26 105
use INVX2  INVX2_124
timestamp 1745462530
transform 1 0 1256 0 1 2970
box -9 -3 26 105
use INVX2  INVX2_125
timestamp 1745462530
transform 1 0 1288 0 -1 3770
box -9 -3 26 105
use INVX2  INVX2_126
timestamp 1745462530
transform 1 0 1904 0 -1 3770
box -9 -3 26 105
use INVX2  INVX2_127
timestamp 1745462530
transform 1 0 616 0 1 3170
box -9 -3 26 105
use INVX2  INVX2_128
timestamp 1745462530
transform 1 0 208 0 1 3170
box -9 -3 26 105
use INVX2  INVX2_129
timestamp 1745462530
transform 1 0 216 0 -1 3170
box -9 -3 26 105
use INVX2  INVX2_130
timestamp 1745462530
transform 1 0 304 0 1 3170
box -9 -3 26 105
use INVX2  INVX2_131
timestamp 1745462530
transform 1 0 408 0 1 3170
box -9 -3 26 105
use INVX2  INVX2_132
timestamp 1745462530
transform 1 0 600 0 1 3170
box -9 -3 26 105
use INVX2  INVX2_133
timestamp 1745462530
transform 1 0 856 0 1 3170
box -9 -3 26 105
use INVX2  INVX2_134
timestamp 1745462530
transform 1 0 1616 0 1 3370
box -9 -3 26 105
use INVX2  INVX2_135
timestamp 1745462530
transform 1 0 1016 0 1 2770
box -9 -3 26 105
use INVX2  INVX2_136
timestamp 1745462530
transform 1 0 1152 0 1 2770
box -9 -3 26 105
use INVX2  INVX2_137
timestamp 1745462530
transform 1 0 1184 0 1 2170
box -9 -3 26 105
use INVX2  INVX2_138
timestamp 1745462530
transform 1 0 1200 0 -1 2770
box -9 -3 26 105
use INVX2  INVX2_139
timestamp 1745462530
transform 1 0 1128 0 -1 2170
box -9 -3 26 105
use INVX2  INVX2_140
timestamp 1745462530
transform 1 0 1152 0 -1 2570
box -9 -3 26 105
use INVX2  INVX2_141
timestamp 1745462530
transform 1 0 1120 0 -1 1970
box -9 -3 26 105
use INVX2  INVX2_142
timestamp 1745462530
transform 1 0 864 0 -1 2970
box -9 -3 26 105
use INVX2  INVX2_143
timestamp 1745462530
transform 1 0 808 0 1 2570
box -9 -3 26 105
use INVX2  INVX2_144
timestamp 1745462530
transform 1 0 176 0 -1 2770
box -9 -3 26 105
use INVX2  INVX2_145
timestamp 1745462530
transform 1 0 176 0 -1 2370
box -9 -3 26 105
use INVX2  INVX2_146
timestamp 1745462530
transform 1 0 184 0 -1 2170
box -9 -3 26 105
use INVX2  INVX2_147
timestamp 1745462530
transform 1 0 264 0 -1 1770
box -9 -3 26 105
use INVX2  INVX2_148
timestamp 1745462530
transform 1 0 744 0 1 1570
box -9 -3 26 105
use INVX2  INVX2_149
timestamp 1745462530
transform 1 0 176 0 1 1370
box -9 -3 26 105
use INVX2  INVX2_150
timestamp 1745462530
transform 1 0 232 0 1 970
box -9 -3 26 105
use INVX2  INVX2_151
timestamp 1745462530
transform 1 0 200 0 -1 570
box -9 -3 26 105
use INVX2  INVX2_152
timestamp 1745462530
transform 1 0 296 0 1 570
box -9 -3 26 105
use INVX2  INVX2_153
timestamp 1745462530
transform 1 0 736 0 1 570
box -9 -3 26 105
use INVX2  INVX2_154
timestamp 1745462530
transform 1 0 960 0 -1 570
box -9 -3 26 105
use INVX2  INVX2_155
timestamp 1745462530
transform 1 0 184 0 -1 1370
box -9 -3 26 105
use INVX2  INVX2_156
timestamp 1745462530
transform 1 0 984 0 -1 1370
box -9 -3 26 105
use INVX2  INVX2_157
timestamp 1745462530
transform 1 0 1080 0 -1 370
box -9 -3 26 105
use INVX2  INVX2_158
timestamp 1745462530
transform 1 0 1104 0 1 370
box -9 -3 26 105
use INVX2  INVX2_159
timestamp 1745462530
transform 1 0 1208 0 1 370
box -9 -3 26 105
use INVX2  INVX2_160
timestamp 1745462530
transform 1 0 1304 0 -1 770
box -9 -3 26 105
use INVX2  INVX2_161
timestamp 1745462530
transform 1 0 1368 0 -1 370
box -9 -3 26 105
use INVX2  INVX2_162
timestamp 1745462530
transform 1 0 1368 0 1 970
box -9 -3 26 105
use INVX2  INVX2_163
timestamp 1745462530
transform 1 0 1408 0 -1 1370
box -9 -3 26 105
use INVX2  INVX2_164
timestamp 1745462530
transform 1 0 1472 0 1 1370
box -9 -3 26 105
use INVX2  INVX2_165
timestamp 1745462530
transform 1 0 2192 0 -1 370
box -9 -3 26 105
use INVX2  INVX2_166
timestamp 1745462530
transform 1 0 2240 0 -1 770
box -9 -3 26 105
use INVX2  INVX2_167
timestamp 1745462530
transform 1 0 2192 0 1 170
box -9 -3 26 105
use INVX2  INVX2_168
timestamp 1745462530
transform 1 0 2336 0 -1 570
box -9 -3 26 105
use INVX2  INVX2_169
timestamp 1745462530
transform 1 0 2576 0 -1 370
box -9 -3 26 105
use INVX2  INVX2_170
timestamp 1745462530
transform 1 0 2520 0 -1 970
box -9 -3 26 105
use INVX2  INVX2_171
timestamp 1745462530
transform 1 0 2408 0 -1 1170
box -9 -3 26 105
use INVX2  INVX2_172
timestamp 1745462530
transform 1 0 2448 0 1 1370
box -9 -3 26 105
use INVX2  INVX2_173
timestamp 1745462530
transform 1 0 3312 0 1 370
box -9 -3 26 105
use INVX2  INVX2_174
timestamp 1745462530
transform 1 0 3416 0 -1 570
box -9 -3 26 105
use INVX2  INVX2_175
timestamp 1745462530
transform 1 0 3960 0 -1 570
box -9 -3 26 105
use INVX2  INVX2_176
timestamp 1745462530
transform 1 0 3568 0 -1 770
box -9 -3 26 105
use INVX2  INVX2_177
timestamp 1745462530
transform 1 0 4056 0 1 570
box -9 -3 26 105
use INVX2  INVX2_178
timestamp 1745462530
transform 1 0 3912 0 1 770
box -9 -3 26 105
use INVX2  INVX2_179
timestamp 1745462530
transform 1 0 3496 0 1 970
box -9 -3 26 105
use INVX2  INVX2_180
timestamp 1745462530
transform 1 0 3416 0 1 1170
box -9 -3 26 105
use INVX2  INVX2_181
timestamp 1745462530
transform 1 0 3936 0 -1 1570
box -9 -3 26 105
use INVX2  INVX2_182
timestamp 1745462530
transform 1 0 3448 0 -1 1970
box -9 -3 26 105
use INVX2  INVX2_183
timestamp 1745462530
transform 1 0 4088 0 -1 1970
box -9 -3 26 105
use INVX2  INVX2_184
timestamp 1745462530
transform 1 0 3640 0 1 1970
box -9 -3 26 105
use INVX2  INVX2_185
timestamp 1745462530
transform 1 0 4112 0 1 1970
box -9 -3 26 105
use INVX2  INVX2_186
timestamp 1745462530
transform 1 0 3320 0 1 2170
box -9 -3 26 105
use INVX2  INVX2_187
timestamp 1745462530
transform 1 0 2784 0 -1 2170
box -9 -3 26 105
use INVX2  INVX2_188
timestamp 1745462530
transform 1 0 2584 0 1 2170
box -9 -3 26 105
use INVX2  INVX2_189
timestamp 1745462530
transform 1 0 3480 0 -1 2770
box -9 -3 26 105
use INVX2  INVX2_190
timestamp 1745462530
transform 1 0 3256 0 -1 2970
box -9 -3 26 105
use INVX2  INVX2_191
timestamp 1745462530
transform 1 0 3368 0 1 2770
box -9 -3 26 105
use INVX2  INVX2_192
timestamp 1745462530
transform 1 0 3320 0 -1 2970
box -9 -3 26 105
use INVX2  INVX2_193
timestamp 1745462530
transform 1 0 3432 0 1 2370
box -9 -3 26 105
use INVX2  INVX2_194
timestamp 1745462530
transform 1 0 3336 0 1 2370
box -9 -3 26 105
use INVX2  INVX2_195
timestamp 1745462530
transform 1 0 3280 0 1 2770
box -9 -3 26 105
use INVX2  INVX2_196
timestamp 1745462530
transform 1 0 2816 0 -1 2570
box -9 -3 26 105
use INVX2  INVX2_197
timestamp 1745462530
transform 1 0 2960 0 1 2970
box -9 -3 26 105
use INVX2  INVX2_198
timestamp 1745462530
transform 1 0 2656 0 1 2770
box -9 -3 26 105
use INVX2  INVX2_199
timestamp 1745462530
transform 1 0 904 0 1 2770
box -9 -3 26 105
use INVX2  INVX2_200
timestamp 1745462530
transform 1 0 1840 0 1 2770
box -9 -3 26 105
use INVX2  INVX2_201
timestamp 1745462530
transform 1 0 1928 0 1 2170
box -9 -3 26 105
use INVX2  INVX2_202
timestamp 1745462530
transform 1 0 1864 0 1 2570
box -9 -3 26 105
use INVX2  INVX2_203
timestamp 1745462530
transform 1 0 1880 0 1 1970
box -9 -3 26 105
use INVX2  INVX2_204
timestamp 1745462530
transform 1 0 1832 0 -1 2570
box -9 -3 26 105
use INVX2  INVX2_205
timestamp 1745462530
transform 1 0 1848 0 -1 1970
box -9 -3 26 105
use INVX2  INVX2_206
timestamp 1745462530
transform 1 0 792 0 -1 2970
box -9 -3 26 105
use INVX2  INVX2_207
timestamp 1745462530
transform 1 0 712 0 -1 2970
box -9 -3 26 105
use INVX2  INVX2_208
timestamp 1745462530
transform 1 0 472 0 1 2770
box -9 -3 26 105
use INVX2  INVX2_209
timestamp 1745462530
transform 1 0 360 0 1 2170
box -9 -3 26 105
use INVX2  INVX2_210
timestamp 1745462530
transform 1 0 384 0 1 1970
box -9 -3 26 105
use INVX2  INVX2_211
timestamp 1745462530
transform 1 0 376 0 1 1770
box -9 -3 26 105
use INVX2  INVX2_212
timestamp 1745462530
transform 1 0 720 0 -1 1770
box -9 -3 26 105
use INVX2  INVX2_213
timestamp 1745462530
transform 1 0 296 0 1 1370
box -9 -3 26 105
use INVX2  INVX2_214
timestamp 1745462530
transform 1 0 232 0 1 770
box -9 -3 26 105
use INVX2  INVX2_215
timestamp 1745462530
transform 1 0 152 0 -1 370
box -9 -3 26 105
use INVX2  INVX2_216
timestamp 1745462530
transform 1 0 272 0 1 370
box -9 -3 26 105
use INVX2  INVX2_217
timestamp 1745462530
transform 1 0 752 0 -1 370
box -9 -3 26 105
use INVX2  INVX2_218
timestamp 1745462530
transform 1 0 936 0 -1 370
box -9 -3 26 105
use INVX2  INVX2_219
timestamp 1745462530
transform 1 0 144 0 -1 1170
box -9 -3 26 105
use INVX2  INVX2_220
timestamp 1745462530
transform 1 0 896 0 1 1370
box -9 -3 26 105
use INVX2  INVX2_221
timestamp 1745462530
transform 1 0 1568 0 -1 370
box -9 -3 26 105
use INVX2  INVX2_222
timestamp 1745462530
transform 1 0 2064 0 -1 570
box -9 -3 26 105
use INVX2  INVX2_223
timestamp 1745462530
transform 1 0 1944 0 1 170
box -9 -3 26 105
use INVX2  INVX2_224
timestamp 1745462530
transform 1 0 1936 0 -1 770
box -9 -3 26 105
use INVX2  INVX2_225
timestamp 1745462530
transform 1 0 1944 0 -1 370
box -9 -3 26 105
use INVX2  INVX2_226
timestamp 1745462530
transform 1 0 1960 0 -1 970
box -9 -3 26 105
use INVX2  INVX2_227
timestamp 1745462530
transform 1 0 2120 0 -1 1170
box -9 -3 26 105
use INVX2  INVX2_228
timestamp 1745462530
transform 1 0 2048 0 -1 1370
box -9 -3 26 105
use INVX2  INVX2_229
timestamp 1745462530
transform 1 0 2408 0 -1 370
box -9 -3 26 105
use INVX2  INVX2_230
timestamp 1745462530
transform 1 0 2432 0 -1 770
box -9 -3 26 105
use INVX2  INVX2_231
timestamp 1745462530
transform 1 0 2560 0 1 170
box -9 -3 26 105
use INVX2  INVX2_232
timestamp 1745462530
transform 1 0 2352 0 -1 570
box -9 -3 26 105
use INVX2  INVX2_233
timestamp 1745462530
transform 1 0 2552 0 1 370
box -9 -3 26 105
use INVX2  INVX2_234
timestamp 1745462530
transform 1 0 2296 0 1 770
box -9 -3 26 105
use INVX2  INVX2_235
timestamp 1745462530
transform 1 0 2560 0 -1 1170
box -9 -3 26 105
use INVX2  INVX2_236
timestamp 1745462530
transform 1 0 2560 0 -1 1370
box -9 -3 26 105
use INVX2  INVX2_237
timestamp 1745462530
transform 1 0 3520 0 -1 370
box -9 -3 26 105
use INVX2  INVX2_238
timestamp 1745462530
transform 1 0 3656 0 -1 570
box -9 -3 26 105
use INVX2  INVX2_239
timestamp 1745462530
transform 1 0 4256 0 1 370
box -9 -3 26 105
use INVX2  INVX2_240
timestamp 1745462530
transform 1 0 3800 0 -1 770
box -9 -3 26 105
use INVX2  INVX2_241
timestamp 1745462530
transform 1 0 4256 0 -1 570
box -9 -3 26 105
use INVX2  INVX2_242
timestamp 1745462530
transform 1 0 4104 0 1 770
box -9 -3 26 105
use INVX2  INVX2_243
timestamp 1745462530
transform 1 0 3752 0 1 970
box -9 -3 26 105
use INVX2  INVX2_244
timestamp 1745462530
transform 1 0 3736 0 1 1170
box -9 -3 26 105
use INVX2  INVX2_245
timestamp 1745462530
transform 1 0 4168 0 -1 1370
box -9 -3 26 105
use INVX2  INVX2_246
timestamp 1745462530
transform 1 0 3840 0 1 1370
box -9 -3 26 105
use INVX2  INVX2_247
timestamp 1745462530
transform 1 0 4248 0 1 1370
box -9 -3 26 105
use INVX2  INVX2_248
timestamp 1745462530
transform 1 0 3840 0 1 1570
box -9 -3 26 105
use INVX2  INVX2_249
timestamp 1745462530
transform 1 0 3920 0 -1 1570
box -9 -3 26 105
use INVX2  INVX2_250
timestamp 1745462530
transform 1 0 3912 0 -1 1770
box -9 -3 26 105
use INVX2  INVX2_251
timestamp 1745462530
transform 1 0 3024 0 1 1770
box -9 -3 26 105
use INVX2  INVX2_252
timestamp 1745462530
transform 1 0 2648 0 1 1770
box -9 -3 26 105
use INVX2  INVX2_253
timestamp 1745462530
transform 1 0 3824 0 -1 2770
box -9 -3 26 105
use INVX2  INVX2_254
timestamp 1745462530
transform 1 0 3736 0 1 2970
box -9 -3 26 105
use INVX2  INVX2_255
timestamp 1745462530
transform 1 0 3824 0 1 2770
box -9 -3 26 105
use INVX2  INVX2_256
timestamp 1745462530
transform 1 0 3760 0 -1 2970
box -9 -3 26 105
use INVX2  INVX2_257
timestamp 1745462530
transform 1 0 3800 0 -1 2570
box -9 -3 26 105
use INVX2  INVX2_258
timestamp 1745462530
transform 1 0 3904 0 -1 2370
box -9 -3 26 105
use INVX2  INVX2_259
timestamp 1745462530
transform 1 0 3816 0 1 2970
box -9 -3 26 105
use INVX2  INVX2_260
timestamp 1745462530
transform 1 0 3024 0 1 2370
box -9 -3 26 105
use INVX2  INVX2_261
timestamp 1745462530
transform 1 0 2944 0 1 2970
box -9 -3 26 105
use INVX2  INVX2_262
timestamp 1745462530
transform 1 0 2464 0 1 2770
box -9 -3 26 105
use INVX2  INVX2_263
timestamp 1745462530
transform 1 0 912 0 1 2570
box -9 -3 26 105
use INVX2  INVX2_264
timestamp 1745462530
transform 1 0 1712 0 1 2770
box -9 -3 26 105
use INVX2  INVX2_265
timestamp 1745462530
transform 1 0 1656 0 1 2170
box -9 -3 26 105
use INVX2  INVX2_266
timestamp 1745462530
transform 1 0 1648 0 -1 2770
box -9 -3 26 105
use INVX2  INVX2_267
timestamp 1745462530
transform 1 0 1640 0 1 1970
box -9 -3 26 105
use INVX2  INVX2_268
timestamp 1745462530
transform 1 0 1568 0 -1 2570
box -9 -3 26 105
use INVX2  INVX2_269
timestamp 1745462530
transform 1 0 1520 0 1 1770
box -9 -3 26 105
use INVX2  INVX2_270
timestamp 1745462530
transform 1 0 400 0 -1 2770
box -9 -3 26 105
use INVX2  INVX2_271
timestamp 1745462530
transform 1 0 544 0 1 2570
box -9 -3 26 105
use INVX2  INVX2_272
timestamp 1745462530
transform 1 0 312 0 1 2570
box -9 -3 26 105
use INVX2  INVX2_273
timestamp 1745462530
transform 1 0 384 0 -1 2370
box -9 -3 26 105
use INVX2  INVX2_274
timestamp 1745462530
transform 1 0 496 0 -1 2170
box -9 -3 26 105
use INVX2  INVX2_275
timestamp 1745462530
transform 1 0 456 0 -1 1770
box -9 -3 26 105
use INVX2  INVX2_276
timestamp 1745462530
transform 1 0 632 0 1 1570
box -9 -3 26 105
use INVX2  INVX2_277
timestamp 1745462530
transform 1 0 416 0 1 1370
box -9 -3 26 105
use INVX2  INVX2_278
timestamp 1745462530
transform 1 0 416 0 1 770
box -9 -3 26 105
use INVX2  INVX2_279
timestamp 1745462530
transform 1 0 264 0 -1 170
box -9 -3 26 105
use INVX2  INVX2_280
timestamp 1745462530
transform 1 0 360 0 1 370
box -9 -3 26 105
use INVX2  INVX2_281
timestamp 1745462530
transform 1 0 568 0 -1 170
box -9 -3 26 105
use INVX2  INVX2_282
timestamp 1745462530
transform 1 0 864 0 1 170
box -9 -3 26 105
use INVX2  INVX2_283
timestamp 1745462530
transform 1 0 360 0 1 1170
box -9 -3 26 105
use INVX2  INVX2_284
timestamp 1745462530
transform 1 0 760 0 -1 1570
box -9 -3 26 105
use INVX2  INVX2_285
timestamp 1745462530
transform 1 0 1744 0 1 170
box -9 -3 26 105
use INVX2  INVX2_286
timestamp 1745462530
transform 1 0 1872 0 1 370
box -9 -3 26 105
use INVX2  INVX2_287
timestamp 1745462530
transform 1 0 1840 0 1 170
box -9 -3 26 105
use INVX2  INVX2_288
timestamp 1745462530
transform 1 0 1784 0 -1 770
box -9 -3 26 105
use INVX2  INVX2_289
timestamp 1745462530
transform 1 0 1944 0 -1 170
box -9 -3 26 105
use INVX2  INVX2_290
timestamp 1745462530
transform 1 0 1992 0 1 970
box -9 -3 26 105
use INVX2  INVX2_291
timestamp 1745462530
transform 1 0 1944 0 1 1170
box -9 -3 26 105
use INVX2  INVX2_292
timestamp 1745462530
transform 1 0 1888 0 1 1370
box -9 -3 26 105
use INVX2  INVX2_293
timestamp 1745462530
transform 1 0 2192 0 -1 170
box -9 -3 26 105
use INVX2  INVX2_294
timestamp 1745462530
transform 1 0 2160 0 1 570
box -9 -3 26 105
use INVX2  INVX2_295
timestamp 1745462530
transform 1 0 2320 0 -1 170
box -9 -3 26 105
use INVX2  INVX2_296
timestamp 1745462530
transform 1 0 2192 0 1 370
box -9 -3 26 105
use INVX2  INVX2_297
timestamp 1745462530
transform 1 0 2456 0 -1 170
box -9 -3 26 105
use INVX2  INVX2_298
timestamp 1745462530
transform 1 0 2400 0 -1 970
box -9 -3 26 105
use INVX2  INVX2_299
timestamp 1745462530
transform 1 0 2248 0 -1 1170
box -9 -3 26 105
use INVX2  INVX2_300
timestamp 1745462530
transform 1 0 2320 0 -1 1370
box -9 -3 26 105
use INVX2  INVX2_301
timestamp 1745462530
transform 1 0 3488 0 1 170
box -9 -3 26 105
use INVX2  INVX2_302
timestamp 1745462530
transform 1 0 3824 0 -1 370
box -9 -3 26 105
use INVX2  INVX2_303
timestamp 1745462530
transform 1 0 4240 0 -1 170
box -9 -3 26 105
use INVX2  INVX2_304
timestamp 1745462530
transform 1 0 3968 0 1 370
box -9 -3 26 105
use INVX2  INVX2_305
timestamp 1745462530
transform 1 0 4360 0 -1 370
box -9 -3 26 105
use INVX2  INVX2_306
timestamp 1745462530
transform 1 0 4176 0 -1 970
box -9 -3 26 105
use INVX2  INVX2_307
timestamp 1745462530
transform 1 0 4256 0 1 970
box -9 -3 26 105
use INVX2  INVX2_308
timestamp 1745462530
transform 1 0 3960 0 1 1170
box -9 -3 26 105
use INVX2  INVX2_309
timestamp 1745462530
transform 1 0 4248 0 -1 1370
box -9 -3 26 105
use INVX2  INVX2_310
timestamp 1745462530
transform 1 0 3632 0 1 1370
box -9 -3 26 105
use INVX2  INVX2_311
timestamp 1745462530
transform 1 0 4264 0 -1 1570
box -9 -3 26 105
use INVX2  INVX2_312
timestamp 1745462530
transform 1 0 3616 0 1 1570
box -9 -3 26 105
use INVX2  INVX2_313
timestamp 1745462530
transform 1 0 4352 0 1 1570
box -9 -3 26 105
use INVX2  INVX2_314
timestamp 1745462530
transform 1 0 3328 0 1 1770
box -9 -3 26 105
use INVX2  INVX2_315
timestamp 1745462530
transform 1 0 2920 0 1 1770
box -9 -3 26 105
use INVX2  INVX2_316
timestamp 1745462530
transform 1 0 2712 0 -1 1970
box -9 -3 26 105
use INVX2  INVX2_317
timestamp 1745462530
transform 1 0 4168 0 1 2570
box -9 -3 26 105
use INVX2  INVX2_318
timestamp 1745462530
transform 1 0 3928 0 -1 2970
box -9 -3 26 105
use INVX2  INVX2_319
timestamp 1745462530
transform 1 0 4112 0 1 2770
box -9 -3 26 105
use INVX2  INVX2_320
timestamp 1745462530
transform 1 0 4256 0 -1 2970
box -9 -3 26 105
use INVX2  INVX2_321
timestamp 1745462530
transform 1 0 4184 0 1 2370
box -9 -3 26 105
use INVX2  INVX2_322
timestamp 1745462530
transform 1 0 4136 0 1 2170
box -9 -3 26 105
use INVX2  INVX2_323
timestamp 1745462530
transform 1 0 4088 0 -1 2970
box -9 -3 26 105
use INVX2  INVX2_324
timestamp 1745462530
transform 1 0 2888 0 1 2370
box -9 -3 26 105
use INVX2  INVX2_325
timestamp 1745462530
transform 1 0 2616 0 -1 2970
box -9 -3 26 105
use INVX2  INVX2_326
timestamp 1745462530
transform 1 0 2568 0 1 2770
box -9 -3 26 105
use INVX2  INVX2_327
timestamp 1745462530
transform 1 0 1000 0 1 2770
box -9 -3 26 105
use INVX2  INVX2_328
timestamp 1745462530
transform 1 0 1376 0 1 2770
box -9 -3 26 105
use INVX2  INVX2_329
timestamp 1745462530
transform 1 0 1336 0 1 2170
box -9 -3 26 105
use INVX2  INVX2_330
timestamp 1745462530
transform 1 0 1304 0 -1 2770
box -9 -3 26 105
use INVX2  INVX2_331
timestamp 1745462530
transform 1 0 1280 0 1 1970
box -9 -3 26 105
use INVX2  INVX2_332
timestamp 1745462530
transform 1 0 1272 0 -1 2570
box -9 -3 26 105
use INVX2  INVX2_333
timestamp 1745462530
transform 1 0 1200 0 1 1770
box -9 -3 26 105
use INVX2  INVX2_334
timestamp 1745462530
transform 1 0 360 0 1 2770
box -9 -3 26 105
use INVX2  INVX2_335
timestamp 1745462530
transform 1 0 624 0 1 2770
box -9 -3 26 105
use INVX2  INVX2_336
timestamp 1745462530
transform 1 0 288 0 -1 2970
box -9 -3 26 105
use INVX2  INVX2_337
timestamp 1745462530
transform 1 0 432 0 1 2370
box -9 -3 26 105
use INVX2  INVX2_338
timestamp 1745462530
transform 1 0 448 0 1 1970
box -9 -3 26 105
use INVX2  INVX2_339
timestamp 1745462530
transform 1 0 448 0 -1 1970
box -9 -3 26 105
use INVX2  INVX2_340
timestamp 1745462530
transform 1 0 768 0 1 1770
box -9 -3 26 105
use INVX2  INVX2_341
timestamp 1745462530
transform 1 0 528 0 1 1370
box -9 -3 26 105
use INVX2  INVX2_342
timestamp 1745462530
transform 1 0 424 0 1 970
box -9 -3 26 105
use INVX2  INVX2_343
timestamp 1745462530
transform 1 0 352 0 1 170
box -9 -3 26 105
use INVX2  INVX2_344
timestamp 1745462530
transform 1 0 440 0 1 370
box -9 -3 26 105
use INVX2  INVX2_345
timestamp 1745462530
transform 1 0 608 0 -1 170
box -9 -3 26 105
use INVX2  INVX2_346
timestamp 1745462530
transform 1 0 928 0 1 170
box -9 -3 26 105
use INVX2  INVX2_347
timestamp 1745462530
transform 1 0 408 0 -1 1170
box -9 -3 26 105
use INVX2  INVX2_348
timestamp 1745462530
transform 1 0 656 0 1 1370
box -9 -3 26 105
use INVX2  INVX2_349
timestamp 1745462530
transform 1 0 1136 0 -1 170
box -9 -3 26 105
use INVX2  INVX2_350
timestamp 1745462530
transform 1 0 1464 0 -1 570
box -9 -3 26 105
use INVX2  INVX2_351
timestamp 1745462530
transform 1 0 1408 0 1 170
box -9 -3 26 105
use INVX2  INVX2_352
timestamp 1745462530
transform 1 0 1464 0 -1 770
box -9 -3 26 105
use INVX2  INVX2_353
timestamp 1745462530
transform 1 0 1536 0 -1 170
box -9 -3 26 105
use INVX2  INVX2_354
timestamp 1745462530
transform 1 0 1552 0 -1 970
box -9 -3 26 105
use INVX2  INVX2_355
timestamp 1745462530
transform 1 0 1536 0 1 1170
box -9 -3 26 105
use INVX2  INVX2_356
timestamp 1745462530
transform 1 0 1664 0 -1 1370
box -9 -3 26 105
use INVX2  INVX2_357
timestamp 1745462530
transform 1 0 2880 0 1 370
box -9 -3 26 105
use INVX2  INVX2_358
timestamp 1745462530
transform 1 0 3112 0 -1 770
box -9 -3 26 105
use INVX2  INVX2_359
timestamp 1745462530
transform 1 0 2808 0 -1 370
box -9 -3 26 105
use INVX2  INVX2_360
timestamp 1745462530
transform 1 0 3040 0 -1 570
box -9 -3 26 105
use INVX2  INVX2_361
timestamp 1745462530
transform 1 0 2992 0 -1 370
box -9 -3 26 105
use INVX2  INVX2_362
timestamp 1745462530
transform 1 0 2880 0 1 770
box -9 -3 26 105
use INVX2  INVX2_363
timestamp 1745462530
transform 1 0 2864 0 -1 1170
box -9 -3 26 105
use INVX2  INVX2_364
timestamp 1745462530
transform 1 0 2888 0 1 1370
box -9 -3 26 105
use INVX2  INVX2_365
timestamp 1745462530
transform 1 0 3224 0 -1 370
box -9 -3 26 105
use INVX2  INVX2_366
timestamp 1745462530
transform 1 0 3176 0 -1 570
box -9 -3 26 105
use INVX2  INVX2_367
timestamp 1745462530
transform 1 0 4088 0 -1 570
box -9 -3 26 105
use INVX2  INVX2_368
timestamp 1745462530
transform 1 0 3336 0 1 570
box -9 -3 26 105
use INVX2  INVX2_369
timestamp 1745462530
transform 1 0 4096 0 -1 770
box -9 -3 26 105
use INVX2  INVX2_370
timestamp 1745462530
transform 1 0 4008 0 1 770
box -9 -3 26 105
use INVX2  INVX2_371
timestamp 1745462530
transform 1 0 3288 0 1 970
box -9 -3 26 105
use INVX2  INVX2_372
timestamp 1745462530
transform 1 0 3328 0 1 1170
box -9 -3 26 105
use INVX2  INVX2_373
timestamp 1745462530
transform 1 0 4048 0 1 1370
box -9 -3 26 105
use INVX2  INVX2_374
timestamp 1745462530
transform 1 0 3464 0 1 1370
box -9 -3 26 105
use INVX2  INVX2_375
timestamp 1745462530
transform 1 0 4032 0 -1 1570
box -9 -3 26 105
use INVX2  INVX2_376
timestamp 1745462530
transform 1 0 3408 0 1 1570
box -9 -3 26 105
use INVX2  INVX2_377
timestamp 1745462530
transform 1 0 4128 0 1 1570
box -9 -3 26 105
use INVX2  INVX2_378
timestamp 1745462530
transform 1 0 3248 0 -1 1770
box -9 -3 26 105
use INVX2  INVX2_379
timestamp 1745462530
transform 1 0 2816 0 -1 1770
box -9 -3 26 105
use INVX2  INVX2_380
timestamp 1745462530
transform 1 0 2816 0 1 1770
box -9 -3 26 105
use INVX2  INVX2_381
timestamp 1745462530
transform 1 0 3184 0 1 2570
box -9 -3 26 105
use INVX2  INVX2_382
timestamp 1745462530
transform 1 0 2976 0 -1 2970
box -9 -3 26 105
use INVX2  INVX2_383
timestamp 1745462530
transform 1 0 3168 0 1 2770
box -9 -3 26 105
use INVX2  INVX2_384
timestamp 1745462530
transform 1 0 3176 0 1 2970
box -9 -3 26 105
use INVX2  INVX2_385
timestamp 1745462530
transform 1 0 3248 0 1 2370
box -9 -3 26 105
use INVX2  INVX2_386
timestamp 1745462530
transform 1 0 3168 0 1 2370
box -9 -3 26 105
use INVX2  INVX2_387
timestamp 1745462530
transform 1 0 3152 0 -1 2970
box -9 -3 26 105
use INVX2  INVX2_388
timestamp 1745462530
transform 1 0 2696 0 1 2370
box -9 -3 26 105
use INVX2  INVX2_389
timestamp 1745462530
transform 1 0 2600 0 -1 2970
box -9 -3 26 105
use INVX2  INVX2_390
timestamp 1745462530
transform 1 0 2768 0 -1 2770
box -9 -3 26 105
use INVX2  INVX2_391
timestamp 1745462530
transform 1 0 1560 0 1 2770
box -9 -3 26 105
use INVX2  INVX2_392
timestamp 1745462530
transform 1 0 1512 0 1 2170
box -9 -3 26 105
use INVX2  INVX2_393
timestamp 1745462530
transform 1 0 1520 0 1 2570
box -9 -3 26 105
use INVX2  INVX2_394
timestamp 1745462530
transform 1 0 1488 0 1 1970
box -9 -3 26 105
use INVX2  INVX2_395
timestamp 1745462530
transform 1 0 1392 0 1 2570
box -9 -3 26 105
use INVX2  INVX2_396
timestamp 1745462530
transform 1 0 1408 0 1 1770
box -9 -3 26 105
use INVX2  INVX2_397
timestamp 1745462530
transform 1 0 192 0 -1 2770
box -9 -3 26 105
use INVX2  INVX2_398
timestamp 1745462530
transform 1 0 608 0 -1 2770
box -9 -3 26 105
use INVX2  INVX2_399
timestamp 1745462530
transform 1 0 184 0 1 2770
box -9 -3 26 105
use INVX2  INVX2_400
timestamp 1745462530
transform 1 0 952 0 -1 2770
box -9 -3 26 105
use INVX2  INVX2_401
timestamp 1745462530
transform 1 0 248 0 1 2370
box -9 -3 26 105
use INVX2  INVX2_402
timestamp 1745462530
transform 1 0 176 0 1 1970
box -9 -3 26 105
use INVX2  INVX2_403
timestamp 1745462530
transform 1 0 184 0 -1 1970
box -9 -3 26 105
use INVX2  INVX2_404
timestamp 1745462530
transform 1 0 576 0 -1 1770
box -9 -3 26 105
use INVX2  INVX2_405
timestamp 1745462530
transform 1 0 184 0 -1 1570
box -9 -3 26 105
use INVX2  INVX2_406
timestamp 1745462530
transform 1 0 408 0 1 970
box -9 -3 26 105
use INVX2  INVX2_407
timestamp 1745462530
transform 1 0 552 0 1 170
box -9 -3 26 105
use INVX2  INVX2_408
timestamp 1745462530
transform 1 0 528 0 1 370
box -9 -3 26 105
use INVX2  INVX2_409
timestamp 1745462530
transform 1 0 664 0 -1 370
box -9 -3 26 105
use INVX2  INVX2_410
timestamp 1745462530
transform 1 0 768 0 -1 370
box -9 -3 26 105
use INVX2  INVX2_411
timestamp 1745462530
transform 1 0 456 0 1 1170
box -9 -3 26 105
use INVX2  INVX2_412
timestamp 1745462530
transform 1 0 896 0 -1 1370
box -9 -3 26 105
use INVX2  INVX2_413
timestamp 1745462530
transform 1 0 1064 0 1 170
box -9 -3 26 105
use INVX2  INVX2_414
timestamp 1745462530
transform 1 0 976 0 -1 570
box -9 -3 26 105
use INVX2  INVX2_415
timestamp 1745462530
transform 1 0 1216 0 1 170
box -9 -3 26 105
use INVX2  INVX2_416
timestamp 1745462530
transform 1 0 1208 0 -1 770
box -9 -3 26 105
use INVX2  INVX2_417
timestamp 1745462530
transform 1 0 1272 0 -1 170
box -9 -3 26 105
use INVX2  INVX2_418
timestamp 1745462530
transform 1 0 1368 0 -1 970
box -9 -3 26 105
use INVX2  INVX2_419
timestamp 1745462530
transform 1 0 1344 0 1 1170
box -9 -3 26 105
use INVX2  INVX2_420
timestamp 1745462530
transform 1 0 1984 0 1 1370
box -9 -3 26 105
use INVX2  INVX2_421
timestamp 1745462530
transform 1 0 2688 0 1 170
box -9 -3 26 105
use INVX2  INVX2_422
timestamp 1745462530
transform 1 0 2784 0 -1 770
box -9 -3 26 105
use INVX2  INVX2_423
timestamp 1745462530
transform 1 0 2648 0 -1 170
box -9 -3 26 105
use INVX2  INVX2_424
timestamp 1745462530
transform 1 0 2744 0 -1 570
box -9 -3 26 105
use INVX2  INVX2_425
timestamp 1745462530
transform 1 0 2976 0 1 170
box -9 -3 26 105
use INVX2  INVX2_426
timestamp 1745462530
transform 1 0 2752 0 -1 970
box -9 -3 26 105
use INVX2  INVX2_427
timestamp 1745462530
transform 1 0 2712 0 -1 1170
box -9 -3 26 105
use INVX2  INVX2_428
timestamp 1745462530
transform 1 0 2688 0 1 1370
box -9 -3 26 105
use INVX2  INVX2_429
timestamp 1745462530
transform 1 0 3264 0 1 170
box -9 -3 26 105
use INVX2  INVX2_430
timestamp 1745462530
transform 1 0 3600 0 -1 370
box -9 -3 26 105
use INVX2  INVX2_431
timestamp 1745462530
transform 1 0 3704 0 1 170
box -9 -3 26 105
use INVX2  INVX2_432
timestamp 1745462530
transform 1 0 3688 0 -1 370
box -9 -3 26 105
use INVX2  INVX2_433
timestamp 1745462530
transform 1 0 4240 0 -1 770
box -9 -3 26 105
use INVX2  INVX2_434
timestamp 1745462530
transform 1 0 4192 0 1 770
box -9 -3 26 105
use INVX2  INVX2_435
timestamp 1745462530
transform 1 0 4120 0 1 970
box -9 -3 26 105
use INVX2  INVX2_436
timestamp 1745462530
transform 1 0 3584 0 1 1170
box -9 -3 26 105
use INVX2  INVX2_437
timestamp 1745462530
transform 1 0 4256 0 1 1770
box -9 -3 26 105
use INVX2  INVX2_438
timestamp 1745462530
transform 1 0 3632 0 1 1770
box -9 -3 26 105
use INVX2  INVX2_439
timestamp 1745462530
transform 1 0 4264 0 -1 1970
box -9 -3 26 105
use INVX2  INVX2_440
timestamp 1745462530
transform 1 0 3736 0 1 1970
box -9 -3 26 105
use INVX2  INVX2_441
timestamp 1745462530
transform 1 0 4320 0 1 1970
box -9 -3 26 105
use INVX2  INVX2_442
timestamp 1745462530
transform 1 0 3528 0 1 2170
box -9 -3 26 105
use INVX2  INVX2_443
timestamp 1745462530
transform 1 0 2896 0 -1 2170
box -9 -3 26 105
use INVX2  INVX2_444
timestamp 1745462530
transform 1 0 2680 0 -1 2170
box -9 -3 26 105
use INVX2  INVX2_445
timestamp 1745462530
transform 1 0 3632 0 -1 2770
box -9 -3 26 105
use INVX2  INVX2_446
timestamp 1745462530
transform 1 0 3672 0 1 2970
box -9 -3 26 105
use INVX2  INVX2_447
timestamp 1745462530
transform 1 0 3600 0 1 2770
box -9 -3 26 105
use INVX2  INVX2_448
timestamp 1745462530
transform 1 0 3560 0 -1 2970
box -9 -3 26 105
use INVX2  INVX2_449
timestamp 1745462530
transform 1 0 3608 0 1 2370
box -9 -3 26 105
use INVX2  INVX2_450
timestamp 1745462530
transform 1 0 3592 0 1 2370
box -9 -3 26 105
use INVX2  INVX2_451
timestamp 1745462530
transform 1 0 3496 0 -1 2970
box -9 -3 26 105
use INVX2  INVX2_452
timestamp 1745462530
transform 1 0 2920 0 -1 2570
box -9 -3 26 105
use INVX2  INVX2_453
timestamp 1745462530
transform 1 0 3152 0 -1 3170
box -9 -3 26 105
use INVX2  INVX2_454
timestamp 1745462530
transform 1 0 3176 0 -1 3170
box -9 -3 26 105
use INVX2  INVX2_455
timestamp 1745462530
transform 1 0 2784 0 -1 3170
box -9 -3 26 105
use INVX2  INVX2_456
timestamp 1745462530
transform 1 0 2872 0 1 2970
box -9 -3 26 105
use INVX2  INVX2_457
timestamp 1745462530
transform 1 0 2976 0 1 2970
box -9 -3 26 105
use INVX2  INVX2_458
timestamp 1745462530
transform 1 0 2952 0 -1 3170
box -9 -3 26 105
use INVX2  INVX2_459
timestamp 1745462530
transform 1 0 3184 0 1 3170
box -9 -3 26 105
use INVX2  INVX2_460
timestamp 1745462530
transform 1 0 3112 0 -1 3170
box -9 -3 26 105
use INVX2  INVX2_461
timestamp 1745462530
transform 1 0 2800 0 -1 3170
box -9 -3 26 105
use INVX2  INVX2_462
timestamp 1745462530
transform 1 0 2552 0 1 2770
box -9 -3 26 105
use INVX2  INVX2_463
timestamp 1745462530
transform 1 0 1864 0 1 3770
box -9 -3 26 105
use INVX2  INVX2_464
timestamp 1745462530
transform 1 0 1736 0 -1 3770
box -9 -3 26 105
use INVX2  INVX2_465
timestamp 1745462530
transform 1 0 2488 0 1 3770
box -9 -3 26 105
use INVX2  INVX2_466
timestamp 1745462530
transform 1 0 2472 0 1 3770
box -9 -3 26 105
use INVX2  INVX2_467
timestamp 1745462530
transform 1 0 1888 0 1 2970
box -9 -3 26 105
use INVX2  INVX2_468
timestamp 1745462530
transform 1 0 1968 0 -1 2770
box -9 -3 26 105
use INVX2  INVX2_469
timestamp 1745462530
transform 1 0 2016 0 1 2170
box -9 -3 26 105
use INVX2  INVX2_470
timestamp 1745462530
transform 1 0 2000 0 -1 2570
box -9 -3 26 105
use INVX2  INVX2_471
timestamp 1745462530
transform 1 0 2000 0 -1 2170
box -9 -3 26 105
use INVX2  INVX2_472
timestamp 1745462530
transform 1 0 1816 0 1 2370
box -9 -3 26 105
use INVX2  INVX2_473
timestamp 1745462530
transform 1 0 1840 0 1 1770
box -9 -3 26 105
use INVX2  INVX2_474
timestamp 1745462530
transform 1 0 344 0 -1 2570
box -9 -3 26 105
use INVX2  INVX2_475
timestamp 1745462530
transform 1 0 544 0 -1 2570
box -9 -3 26 105
use INVX2  INVX2_476
timestamp 1745462530
transform 1 0 176 0 -1 2570
box -9 -3 26 105
use INVX2  INVX2_477
timestamp 1745462530
transform 1 0 896 0 1 2370
box -9 -3 26 105
use INVX2  INVX2_478
timestamp 1745462530
transform 1 0 304 0 -1 2370
box -9 -3 26 105
use INVX2  INVX2_479
timestamp 1745462530
transform 1 0 312 0 -1 2170
box -9 -3 26 105
use INVX2  INVX2_480
timestamp 1745462530
transform 1 0 312 0 -1 1970
box -9 -3 26 105
use INVX2  INVX2_481
timestamp 1745462530
transform 1 0 664 0 1 1770
box -9 -3 26 105
use INVX2  INVX2_482
timestamp 1745462530
transform 1 0 304 0 1 1570
box -9 -3 26 105
use INVX2  INVX2_483
timestamp 1745462530
transform 1 0 288 0 -1 970
box -9 -3 26 105
use INVX2  INVX2_484
timestamp 1745462530
transform 1 0 256 0 -1 770
box -9 -3 26 105
use INVX2  INVX2_485
timestamp 1745462530
transform 1 0 608 0 1 570
box -9 -3 26 105
use INVX2  INVX2_486
timestamp 1745462530
transform 1 0 680 0 1 370
box -9 -3 26 105
use INVX2  INVX2_487
timestamp 1745462530
transform 1 0 872 0 -1 570
box -9 -3 26 105
use INVX2  INVX2_488
timestamp 1745462530
transform 1 0 512 0 -1 1370
box -9 -3 26 105
use INVX2  INVX2_489
timestamp 1745462530
transform 1 0 640 0 -1 1370
box -9 -3 26 105
use INVX2  INVX2_490
timestamp 1745462530
transform 1 0 1472 0 1 370
box -9 -3 26 105
use INVX2  INVX2_491
timestamp 1745462530
transform 1 0 1720 0 -1 570
box -9 -3 26 105
use INVX2  INVX2_492
timestamp 1745462530
transform 1 0 1608 0 1 370
box -9 -3 26 105
use INVX2  INVX2_493
timestamp 1745462530
transform 1 0 1688 0 -1 770
box -9 -3 26 105
use INVX2  INVX2_494
timestamp 1745462530
transform 1 0 1680 0 -1 370
box -9 -3 26 105
use INVX2  INVX2_495
timestamp 1745462530
transform 1 0 1760 0 1 970
box -9 -3 26 105
use INVX2  INVX2_496
timestamp 1745462530
transform 1 0 1792 0 1 1170
box -9 -3 26 105
use INVX2  INVX2_497
timestamp 1745462530
transform 1 0 1768 0 1 1370
box -9 -3 26 105
use INVX2  INVX2_498
timestamp 1745462530
transform 1 0 2960 0 1 170
box -9 -3 26 105
use INVX2  INVX2_499
timestamp 1745462530
transform 1 0 3064 0 1 570
box -9 -3 26 105
use INVX2  INVX2_500
timestamp 1745462530
transform 1 0 2856 0 1 170
box -9 -3 26 105
use INVX2  INVX2_501
timestamp 1745462530
transform 1 0 2968 0 1 370
box -9 -3 26 105
use INVX2  INVX2_502
timestamp 1745462530
transform 1 0 3152 0 1 170
box -9 -3 26 105
use INVX2  INVX2_503
timestamp 1745462530
transform 1 0 2952 0 1 970
box -9 -3 26 105
use INVX2  INVX2_504
timestamp 1745462530
transform 1 0 2888 0 1 1170
box -9 -3 26 105
use INVX2  INVX2_505
timestamp 1745462530
transform 1 0 2856 0 -1 1370
box -9 -3 26 105
use INVX2  INVX2_506
timestamp 1745462530
transform 1 0 3376 0 1 170
box -9 -3 26 105
use INVX2  INVX2_507
timestamp 1745462530
transform 1 0 3936 0 1 170
box -9 -3 26 105
use INVX2  INVX2_508
timestamp 1745462530
transform 1 0 4104 0 1 170
box -9 -3 26 105
use INVX2  INVX2_509
timestamp 1745462530
transform 1 0 4048 0 1 170
box -9 -3 26 105
use INVX2  INVX2_510
timestamp 1745462530
transform 1 0 4120 0 1 370
box -9 -3 26 105
use INVX2  INVX2_511
timestamp 1745462530
transform 1 0 4360 0 1 970
box -9 -3 26 105
use INVX2  INVX2_512
timestamp 1745462530
transform 1 0 4104 0 -1 1170
box -9 -3 26 105
use INVX2  INVX2_513
timestamp 1745462530
transform 1 0 3840 0 1 1170
box -9 -3 26 105
use INVX2  INVX2_514
timestamp 1745462530
transform 1 0 4248 0 -1 1770
box -9 -3 26 105
use INVX2  INVX2_515
timestamp 1745462530
transform 1 0 3920 0 1 1770
box -9 -3 26 105
use INVX2  INVX2_516
timestamp 1745462530
transform 1 0 4256 0 1 2170
box -9 -3 26 105
use INVX2  INVX2_517
timestamp 1745462530
transform 1 0 3896 0 1 1970
box -9 -3 26 105
use INVX2  INVX2_518
timestamp 1745462530
transform 1 0 4192 0 1 1970
box -9 -3 26 105
use INVX2  INVX2_519
timestamp 1745462530
transform 1 0 3888 0 1 2170
box -9 -3 26 105
use INVX2  INVX2_520
timestamp 1745462530
transform 1 0 3168 0 1 2170
box -9 -3 26 105
use INVX2  INVX2_521
timestamp 1745462530
transform 1 0 2976 0 1 2170
box -9 -3 26 105
use INVX2  INVX2_522
timestamp 1745462530
transform 1 0 4160 0 -1 2770
box -9 -3 26 105
use INVX2  INVX2_523
timestamp 1745462530
transform 1 0 3952 0 1 2970
box -9 -3 26 105
use INVX2  INVX2_524
timestamp 1745462530
transform 1 0 4088 0 -1 2770
box -9 -3 26 105
use INVX2  INVX2_525
timestamp 1745462530
transform 1 0 4200 0 1 2970
box -9 -3 26 105
use INVX2  INVX2_526
timestamp 1745462530
transform 1 0 4240 0 -1 2570
box -9 -3 26 105
use INVX2  INVX2_527
timestamp 1745462530
transform 1 0 4256 0 -1 2370
box -9 -3 26 105
use INVX2  INVX2_528
timestamp 1745462530
transform 1 0 4128 0 1 2970
box -9 -3 26 105
use INVX2  INVX2_529
timestamp 1745462530
transform 1 0 2928 0 1 2570
box -9 -3 26 105
use INVX2  INVX2_530
timestamp 1745462530
transform 1 0 1128 0 -1 3770
box -9 -3 26 105
use INVX2  INVX2_531
timestamp 1745462530
transform 1 0 2472 0 -1 3170
box -9 -3 26 105
use INVX2  INVX2_532
timestamp 1745462530
transform 1 0 2872 0 -1 3970
box -9 -3 26 105
use INVX2  INVX2_533
timestamp 1745462530
transform 1 0 3120 0 -1 3970
box -9 -3 26 105
use INVX2  INVX2_534
timestamp 1745462530
transform 1 0 3608 0 1 3770
box -9 -3 26 105
use INVX2  INVX2_535
timestamp 1745462530
transform 1 0 3632 0 -1 3970
box -9 -3 26 105
use INVX2  INVX2_536
timestamp 1745462530
transform 1 0 3624 0 -1 3770
box -9 -3 26 105
use INVX2  INVX2_537
timestamp 1745462530
transform 1 0 3264 0 -1 4170
box -9 -3 26 105
use INVX2  INVX2_538
timestamp 1745462530
transform 1 0 2408 0 1 3970
box -9 -3 26 105
use INVX2  INVX2_539
timestamp 1745462530
transform 1 0 2248 0 -1 3970
box -9 -3 26 105
use INVX2  INVX2_540
timestamp 1745462530
transform 1 0 2392 0 1 2970
box -9 -3 26 105
use INVX2  INVX2_541
timestamp 1745462530
transform 1 0 2720 0 -1 4170
box -9 -3 26 105
use INVX2  INVX2_542
timestamp 1745462530
transform 1 0 3048 0 -1 4170
box -9 -3 26 105
use INVX2  INVX2_543
timestamp 1745462530
transform 1 0 3464 0 -1 4170
box -9 -3 26 105
use INVX2  INVX2_544
timestamp 1745462530
transform 1 0 3360 0 -1 4170
box -9 -3 26 105
use INVX2  INVX2_545
timestamp 1745462530
transform 1 0 3472 0 1 3970
box -9 -3 26 105
use INVX2  INVX2_546
timestamp 1745462530
transform 1 0 3208 0 -1 4170
box -9 -3 26 105
use INVX2  INVX2_547
timestamp 1745462530
transform 1 0 2440 0 -1 4170
box -9 -3 26 105
use INVX2  INVX2_548
timestamp 1745462530
transform 1 0 2208 0 -1 4170
box -9 -3 26 105
use INVX2  INVX2_549
timestamp 1745462530
transform 1 0 2568 0 -1 3170
box -9 -3 26 105
use INVX2  INVX2_550
timestamp 1745462530
transform 1 0 2632 0 1 3970
box -9 -3 26 105
use INVX2  INVX2_551
timestamp 1745462530
transform 1 0 2952 0 -1 3970
box -9 -3 26 105
use INVX2  INVX2_552
timestamp 1745462530
transform 1 0 4280 0 -1 3770
box -9 -3 26 105
use INVX2  INVX2_553
timestamp 1745462530
transform 1 0 4192 0 1 3770
box -9 -3 26 105
use INVX2  INVX2_554
timestamp 1745462530
transform 1 0 4208 0 1 3570
box -9 -3 26 105
use INVX2  INVX2_555
timestamp 1745462530
transform 1 0 3936 0 -1 3570
box -9 -3 26 105
use INVX2  INVX2_556
timestamp 1745462530
transform 1 0 1960 0 -1 3770
box -9 -3 26 105
use INVX2  INVX2_557
timestamp 1745462530
transform 1 0 1992 0 -1 3970
box -9 -3 26 105
use INVX2  INVX2_558
timestamp 1745462530
transform 1 0 2584 0 -1 3170
box -9 -3 26 105
use INVX2  INVX2_559
timestamp 1745462530
transform 1 0 1744 0 -1 3970
box -9 -3 26 105
use INVX2  INVX2_560
timestamp 1745462530
transform 1 0 1736 0 1 3970
box -9 -3 26 105
use INVX2  INVX2_561
timestamp 1745462530
transform 1 0 4176 0 -1 3170
box -9 -3 26 105
use INVX2  INVX2_562
timestamp 1745462530
transform 1 0 4192 0 1 3170
box -9 -3 26 105
use INVX2  INVX2_563
timestamp 1745462530
transform 1 0 4064 0 -1 3370
box -9 -3 26 105
use INVX2  INVX2_564
timestamp 1745462530
transform 1 0 3800 0 -1 3770
box -9 -3 26 105
use INVX2  INVX2_565
timestamp 1745462530
transform 1 0 1592 0 -1 3770
box -9 -3 26 105
use INVX2  INVX2_566
timestamp 1745462530
transform 1 0 1624 0 1 3770
box -9 -3 26 105
use INVX2  INVX2_567
timestamp 1745462530
transform 1 0 2544 0 1 2970
box -9 -3 26 105
use INVX2  INVX2_568
timestamp 1745462530
transform 1 0 2736 0 -1 3170
box -9 -3 26 105
use INVX2  INVX2_569
timestamp 1745462530
transform 1 0 2712 0 -1 3970
box -9 -3 26 105
use INVX2  INVX2_570
timestamp 1745462530
transform 1 0 2888 0 -1 3770
box -9 -3 26 105
use INVX2  INVX2_571
timestamp 1745462530
transform 1 0 4024 0 -1 3570
box -9 -3 26 105
use INVX2  INVX2_572
timestamp 1745462530
transform 1 0 4024 0 1 3570
box -9 -3 26 105
use INVX2  INVX2_573
timestamp 1745462530
transform 1 0 4168 0 1 3370
box -9 -3 26 105
use INVX2  INVX2_574
timestamp 1745462530
transform 1 0 3944 0 1 3370
box -9 -3 26 105
use INVX2  INVX2_575
timestamp 1745462530
transform 1 0 2048 0 1 3570
box -9 -3 26 105
use INVX2  INVX2_576
timestamp 1745462530
transform 1 0 1960 0 -1 3970
box -9 -3 26 105
use INVX2  INVX2_577
timestamp 1745462530
transform 1 0 2768 0 -1 3170
box -9 -3 26 105
use INVX2  INVX2_578
timestamp 1745462530
transform 1 0 1896 0 -1 3970
box -9 -3 26 105
use INVX2  INVX2_579
timestamp 1745462530
transform 1 0 1816 0 -1 3970
box -9 -3 26 105
use INVX2  INVX2_580
timestamp 1745462530
transform 1 0 4200 0 -1 3370
box -9 -3 26 105
use INVX2  INVX2_581
timestamp 1745462530
transform 1 0 4192 0 1 3370
box -9 -3 26 105
use INVX2  INVX2_582
timestamp 1745462530
transform 1 0 4008 0 1 3170
box -9 -3 26 105
use INVX2  INVX2_583
timestamp 1745462530
transform 1 0 3928 0 1 3170
box -9 -3 26 105
use INVX2  INVX2_584
timestamp 1745462530
transform 1 0 1696 0 1 3770
box -9 -3 26 105
use INVX2  INVX2_585
timestamp 1745462530
transform 1 0 1680 0 -1 3970
box -9 -3 26 105
use INVX2  INVX2_586
timestamp 1745462530
transform 1 0 2720 0 -1 3170
box -9 -3 26 105
use INVX2  INVX2_587
timestamp 1745462530
transform 1 0 2704 0 -1 4170
box -9 -3 26 105
use INVX2  INVX2_588
timestamp 1745462530
transform 1 0 2960 0 1 3970
box -9 -3 26 105
use INVX2  INVX2_589
timestamp 1745462530
transform 1 0 3736 0 1 3970
box -9 -3 26 105
use INVX2  INVX2_590
timestamp 1745462530
transform 1 0 3888 0 -1 4170
box -9 -3 26 105
use INVX2  INVX2_591
timestamp 1745462530
transform 1 0 3664 0 -1 3970
box -9 -3 26 105
use INVX2  INVX2_592
timestamp 1745462530
transform 1 0 3688 0 -1 4170
box -9 -3 26 105
use INVX2  INVX2_593
timestamp 1745462530
transform 1 0 2520 0 -1 4170
box -9 -3 26 105
use INVX2  INVX2_594
timestamp 1745462530
transform 1 0 2320 0 -1 4170
box -9 -3 26 105
use INVX2  INVX2_595
timestamp 1745462530
transform 1 0 2656 0 -1 3170
box -9 -3 26 105
use INVX2  INVX2_596
timestamp 1745462530
transform 1 0 3152 0 1 3770
box -9 -3 26 105
use INVX2  INVX2_597
timestamp 1745462530
transform 1 0 3400 0 -1 3970
box -9 -3 26 105
use INVX2  INVX2_598
timestamp 1745462530
transform 1 0 3328 0 -1 3970
box -9 -3 26 105
use INVX2  INVX2_599
timestamp 1745462530
transform 1 0 3384 0 1 3770
box -9 -3 26 105
use INVX2  INVX2_600
timestamp 1745462530
transform 1 0 3192 0 -1 3970
box -9 -3 26 105
use INVX2  INVX2_601
timestamp 1745462530
transform 1 0 2416 0 -1 3970
box -9 -3 26 105
use INVX2  INVX2_602
timestamp 1745462530
transform 1 0 2104 0 -1 3970
box -9 -3 26 105
use INVX2  INVX2_603
timestamp 1745462530
transform 1 0 2816 0 -1 3770
box -9 -3 26 105
use INVX2  INVX2_604
timestamp 1745462530
transform 1 0 2744 0 1 2770
box -9 -3 26 105
use INVX2  INVX2_605
timestamp 1745462530
transform 1 0 3016 0 -1 3970
box -9 -3 26 105
use INVX2  INVX2_606
timestamp 1745462530
transform 1 0 1560 0 1 3770
box -9 -3 26 105
use INVX2  INVX2_607
timestamp 1745462530
transform 1 0 2808 0 -1 3970
box -9 -3 26 105
use INVX2  INVX2_608
timestamp 1745462530
transform 1 0 1520 0 -1 3770
box -9 -3 26 105
use INVX2  INVX2_609
timestamp 1745462530
transform 1 0 3872 0 -1 3770
box -9 -3 26 105
use INVX2  INVX2_610
timestamp 1745462530
transform 1 0 4088 0 -1 3370
box -9 -3 26 105
use INVX2  INVX2_611
timestamp 1745462530
transform 1 0 4256 0 1 3170
box -9 -3 26 105
use INVX2  INVX2_612
timestamp 1745462530
transform 1 0 4240 0 -1 3170
box -9 -3 26 105
use INVX2  INVX2_613
timestamp 1745462530
transform 1 0 1632 0 1 3970
box -9 -3 26 105
use INVX2  INVX2_614
timestamp 1745462530
transform 1 0 1752 0 1 3970
box -9 -3 26 105
use INVX2  INVX2_615
timestamp 1745462530
transform 1 0 1480 0 -1 3970
box -9 -3 26 105
use INVX2  INVX2_616
timestamp 1745462530
transform 1 0 1600 0 -1 3970
box -9 -3 26 105
use INVX2  INVX2_617
timestamp 1745462530
transform 1 0 4008 0 -1 3370
box -9 -3 26 105
use INVX2  INVX2_618
timestamp 1745462530
transform 1 0 4072 0 1 3170
box -9 -3 26 105
use INVX2  INVX2_619
timestamp 1745462530
transform 1 0 4256 0 1 3370
box -9 -3 26 105
use INVX2  INVX2_620
timestamp 1745462530
transform 1 0 4264 0 -1 3370
box -9 -3 26 105
use INVX2  INVX2_621
timestamp 1745462530
transform 1 0 1768 0 1 3970
box -9 -3 26 105
use INVX2  INVX2_622
timestamp 1745462530
transform 1 0 1840 0 -1 3970
box -9 -3 26 105
use INVX2  INVX2_623
timestamp 1745462530
transform 1 0 1936 0 1 3970
box -9 -3 26 105
use INVX2  INVX2_624
timestamp 1745462530
transform 1 0 2024 0 -1 3770
box -9 -3 26 105
use INVX2  INVX2_625
timestamp 1745462530
transform 1 0 4000 0 1 3370
box -9 -3 26 105
use INVX2  INVX2_626
timestamp 1745462530
transform 1 0 4128 0 -1 3570
box -9 -3 26 105
use INVX2  INVX2_627
timestamp 1745462530
transform 1 0 4088 0 1 3570
box -9 -3 26 105
use INVX2  INVX2_628
timestamp 1745462530
transform 1 0 4112 0 -1 3570
box -9 -3 26 105
use INVX2  INVX2_629
timestamp 1745462530
transform 1 0 2880 0 1 3770
box -9 -3 26 105
use INVX2  INVX2_630
timestamp 1745462530
transform 1 0 2552 0 -1 3970
box -9 -3 26 105
use INVX2  INVX2_631
timestamp 1745462530
transform 1 0 2048 0 -1 3970
box -9 -3 26 105
use INVX2  INVX2_632
timestamp 1745462530
transform 1 0 2000 0 1 3770
box -9 -3 26 105
use INVX2  INVX2_633
timestamp 1745462530
transform 1 0 3904 0 1 3570
box -9 -3 26 105
use INVX2  INVX2_634
timestamp 1745462530
transform 1 0 4264 0 1 3570
box -9 -3 26 105
use INVX2  INVX2_635
timestamp 1745462530
transform 1 0 4248 0 1 3770
box -9 -3 26 105
use INVX2  INVX2_636
timestamp 1745462530
transform 1 0 4360 0 -1 3770
box -9 -3 26 105
use INVX2  INVX2_637
timestamp 1745462530
transform 1 0 2896 0 -1 3970
box -9 -3 26 105
use INVX2  INVX2_638
timestamp 1745462530
transform 1 0 2560 0 1 3970
box -9 -3 26 105
use INVX2  INVX2_639
timestamp 1745462530
transform 1 0 2264 0 -1 4170
box -9 -3 26 105
use INVX2  INVX2_640
timestamp 1745462530
transform 1 0 2464 0 -1 4170
box -9 -3 26 105
use INVX2  INVX2_641
timestamp 1745462530
transform 1 0 3744 0 -1 4170
box -9 -3 26 105
use INVX2  INVX2_642
timestamp 1745462530
transform 1 0 3728 0 -1 3970
box -9 -3 26 105
use INVX2  INVX2_643
timestamp 1745462530
transform 1 0 3896 0 1 4170
box -9 -3 26 105
use INVX2  INVX2_644
timestamp 1745462530
transform 1 0 3800 0 1 3970
box -9 -3 26 105
use INVX2  INVX2_645
timestamp 1745462530
transform 1 0 2992 0 -1 4170
box -9 -3 26 105
use INVX2  INVX2_646
timestamp 1745462530
transform 1 0 2680 0 -1 4170
box -9 -3 26 105
use INVX2  INVX2_647
timestamp 1745462530
transform 1 0 2152 0 -1 4170
box -9 -3 26 105
use INVX2  INVX2_648
timestamp 1745462530
transform 1 0 2376 0 -1 4170
box -9 -3 26 105
use INVX2  INVX2_649
timestamp 1745462530
transform 1 0 3304 0 -1 4170
box -9 -3 26 105
use INVX2  INVX2_650
timestamp 1745462530
transform 1 0 3584 0 1 3970
box -9 -3 26 105
use INVX2  INVX2_651
timestamp 1745462530
transform 1 0 3472 0 1 4170
box -9 -3 26 105
use INVX2  INVX2_652
timestamp 1745462530
transform 1 0 3560 0 -1 4170
box -9 -3 26 105
use INVX2  INVX2_653
timestamp 1745462530
transform 1 0 3072 0 1 4170
box -9 -3 26 105
use INVX2  INVX2_654
timestamp 1745462530
transform 1 0 2776 0 -1 4170
box -9 -3 26 105
use INVX2  INVX2_655
timestamp 1745462530
transform 1 0 2200 0 1 3970
box -9 -3 26 105
use INVX2  INVX2_656
timestamp 1745462530
transform 1 0 2352 0 1 3970
box -9 -3 26 105
use INVX2  INVX2_657
timestamp 1745462530
transform 1 0 3288 0 -1 4170
box -9 -3 26 105
use INVX2  INVX2_658
timestamp 1745462530
transform 1 0 3688 0 1 3770
box -9 -3 26 105
use INVX2  INVX2_659
timestamp 1745462530
transform 1 0 3624 0 -1 4170
box -9 -3 26 105
use INVX2  INVX2_660
timestamp 1745462530
transform 1 0 3672 0 1 3770
box -9 -3 26 105
use INVX2  INVX2_661
timestamp 1745462530
transform 1 0 3080 0 1 3970
box -9 -3 26 105
use INVX2  INVX2_662
timestamp 1745462530
transform 1 0 2712 0 1 3970
box -9 -3 26 105
use INVX2  INVX2_663
timestamp 1745462530
transform 1 0 2088 0 1 3970
box -9 -3 26 105
use INVX2  INVX2_664
timestamp 1745462530
transform 1 0 2360 0 -1 3970
box -9 -3 26 105
use INVX2  INVX2_665
timestamp 1745462530
transform 1 0 3224 0 -1 3970
box -9 -3 26 105
use INVX2  INVX2_666
timestamp 1745462530
transform 1 0 3416 0 1 3770
box -9 -3 26 105
use INVX2  INVX2_667
timestamp 1745462530
transform 1 0 3456 0 1 3970
box -9 -3 26 105
use INVX2  INVX2_668
timestamp 1745462530
transform 1 0 3440 0 -1 3970
box -9 -3 26 105
use INVX2  INVX2_669
timestamp 1745462530
transform 1 0 2168 0 1 3770
box -9 -3 26 105
use INVX2  INVX2_670
timestamp 1745462530
transform 1 0 456 0 1 3970
box -9 -3 26 105
use INVX2  INVX2_671
timestamp 1745462530
transform 1 0 952 0 -1 3770
box -9 -3 26 105
use INVX2  INVX2_672
timestamp 1745462530
transform 1 0 336 0 -1 4170
box -9 -3 26 105
use INVX2  INVX2_673
timestamp 1745462530
transform 1 0 448 0 -1 4170
box -9 -3 26 105
use INVX2  INVX2_674
timestamp 1745462530
transform 1 0 480 0 1 3770
box -9 -3 26 105
use INVX2  INVX2_675
timestamp 1745462530
transform 1 0 1520 0 -1 3570
box -9 -3 26 105
use INVX2  INVX2_676
timestamp 1745462530
transform 1 0 1360 0 -1 3770
box -9 -3 26 105
use INVX2  INVX2_677
timestamp 1745462530
transform 1 0 1232 0 1 3770
box -9 -3 26 105
use INVX2  INVX2_678
timestamp 1745462530
transform 1 0 1496 0 -1 3570
box -9 -3 26 105
use INVX2  INVX2_679
timestamp 1745462530
transform 1 0 1496 0 -1 3770
box -9 -3 26 105
use INVX2  INVX2_680
timestamp 1745462530
transform 1 0 1320 0 1 3570
box -9 -3 26 105
use INVX2  INVX2_681
timestamp 1745462530
transform 1 0 1472 0 1 3370
box -9 -3 26 105
use INVX2  INVX2_682
timestamp 1745462530
transform 1 0 536 0 1 3970
box -9 -3 26 105
use INVX2  INVX2_683
timestamp 1745462530
transform 1 0 592 0 1 3970
box -9 -3 26 105
use INVX2  INVX2_684
timestamp 1745462530
transform 1 0 1032 0 -1 4170
box -9 -3 26 105
use INVX2  INVX2_685
timestamp 1745462530
transform 1 0 1056 0 1 3970
box -9 -3 26 105
use INVX2  INVX2_686
timestamp 1745462530
transform 1 0 584 0 -1 4170
box -9 -3 26 105
use INVX2  INVX2_687
timestamp 1745462530
transform 1 0 560 0 1 4170
box -9 -3 26 105
use INVX2  INVX2_688
timestamp 1745462530
transform 1 0 632 0 1 3970
box -9 -3 26 105
use INVX2  INVX2_689
timestamp 1745462530
transform 1 0 760 0 1 3770
box -9 -3 26 105
use INVX2  INVX2_690
timestamp 1745462530
transform 1 0 112 0 1 3970
box -9 -3 26 105
use INVX2  INVX2_691
timestamp 1745462530
transform 1 0 168 0 1 4170
box -9 -3 26 105
use INVX2  INVX2_692
timestamp 1745462530
transform 1 0 176 0 -1 4170
box -9 -3 26 105
use INVX2  INVX2_693
timestamp 1745462530
transform 1 0 80 0 1 3770
box -9 -3 26 105
use INVX2  INVX2_694
timestamp 1745462530
transform 1 0 144 0 1 4170
box -9 -3 26 105
use INVX2  INVX2_695
timestamp 1745462530
transform 1 0 120 0 -1 3970
box -9 -3 26 105
use INVX2  INVX2_696
timestamp 1745462530
transform 1 0 304 0 -1 3970
box -9 -3 26 105
use INVX2  INVX2_697
timestamp 1745462530
transform 1 0 320 0 -1 4170
box -9 -3 26 105
use INVX2  INVX2_698
timestamp 1745462530
transform 1 0 608 0 1 4170
box -9 -3 26 105
use INVX2  INVX2_699
timestamp 1745462530
transform 1 0 880 0 -1 4170
box -9 -3 26 105
use INVX2  INVX2_700
timestamp 1745462530
transform 1 0 832 0 -1 4170
box -9 -3 26 105
use INVX2  INVX2_701
timestamp 1745462530
transform 1 0 688 0 1 4170
box -9 -3 26 105
use INVX2  INVX2_702
timestamp 1745462530
transform 1 0 2432 0 -1 2170
box -9 -3 26 105
use INVX2  INVX2_703
timestamp 1745462530
transform 1 0 1064 0 -1 3970
box -9 -3 26 105
use INVX2  INVX2_704
timestamp 1745462530
transform 1 0 808 0 -1 4170
box -9 -3 26 105
use INVX2  INVX2_705
timestamp 1745462530
transform 1 0 1344 0 1 3970
box -9 -3 26 105
use INVX2  INVX2_706
timestamp 1745462530
transform 1 0 664 0 -1 3770
box -9 -3 26 105
use INVX2  INVX2_707
timestamp 1745462530
transform 1 0 2360 0 -1 2770
box -9 -3 26 105
use INVX2  INVX2_708
timestamp 1745462530
transform 1 0 3136 0 -1 3170
box -9 -3 26 105
use INVX2  INVX2_709
timestamp 1745462530
transform 1 0 1120 0 -1 3370
box -9 -3 26 105
use INVX2  INVX2_710
timestamp 1745462530
transform 1 0 1560 0 1 3170
box -9 -3 26 105
use INVX2  INVX2_711
timestamp 1745462530
transform 1 0 696 0 -1 3770
box -9 -3 26 105
use INVX2  INVX2_712
timestamp 1745462530
transform 1 0 680 0 -1 3770
box -9 -3 26 105
use INVX2  INVX2_713
timestamp 1745462530
transform 1 0 2080 0 1 3570
box -9 -3 26 105
use INVX2  INVX2_714
timestamp 1745462530
transform 1 0 2176 0 -1 3570
box -9 -3 26 105
use INVX2  INVX2_715
timestamp 1745462530
transform 1 0 1632 0 1 3370
box -9 -3 26 105
use INVX2  INVX2_716
timestamp 1745462530
transform 1 0 1368 0 1 3970
box -9 -3 26 105
use INVX2  INVX2_717
timestamp 1745462530
transform 1 0 1528 0 -1 4170
box -9 -3 26 105
use INVX2  INVX2_718
timestamp 1745462530
transform 1 0 1376 0 -1 4170
box -9 -3 26 105
use INVX2  INVX2_719
timestamp 1745462530
transform 1 0 2248 0 1 1970
box -9 -3 26 105
use INVX2  INVX2_720
timestamp 1745462530
transform 1 0 1080 0 1 2970
box -9 -3 26 105
use INVX2  INVX2_721
timestamp 1745462530
transform 1 0 1816 0 -1 3770
box -9 -3 26 105
use INVX2  INVX2_722
timestamp 1745462530
transform 1 0 968 0 1 3170
box -9 -3 26 105
use INVX2  INVX2_723
timestamp 1745462530
transform 1 0 2040 0 1 1170
box -9 -3 26 105
use INVX2  INVX2_724
timestamp 1745462530
transform 1 0 2856 0 -1 2770
box -9 -3 26 105
use M2_M1  M2_M1_0
timestamp 1745462530
transform 1 0 828 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_1
timestamp 1745462530
transform 1 0 604 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_2
timestamp 1745462530
transform 1 0 580 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3
timestamp 1745462530
transform 1 0 596 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_4
timestamp 1745462530
transform 1 0 564 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_5
timestamp 1745462530
transform 1 0 540 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_6
timestamp 1745462530
transform 1 0 556 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_7
timestamp 1745462530
transform 1 0 452 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_8
timestamp 1745462530
transform 1 0 428 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_9
timestamp 1745462530
transform 1 0 444 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_10
timestamp 1745462530
transform 1 0 348 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_11
timestamp 1745462530
transform 1 0 324 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_12
timestamp 1745462530
transform 1 0 340 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_13
timestamp 1745462530
transform 1 0 316 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_14
timestamp 1745462530
transform 1 0 508 0 1 3115
box -2 -2 2 2
use M2_M1  M2_M1_15
timestamp 1745462530
transform 1 0 404 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_16
timestamp 1745462530
transform 1 0 420 0 1 3115
box -2 -2 2 2
use M2_M1  M2_M1_17
timestamp 1745462530
transform 1 0 300 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_18
timestamp 1745462530
transform 1 0 316 0 1 3115
box -2 -2 2 2
use M2_M1  M2_M1_19
timestamp 1745462530
transform 1 0 164 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_20
timestamp 1745462530
transform 1 0 188 0 1 3025
box -2 -2 2 2
use M2_M1  M2_M1_21
timestamp 1745462530
transform 1 0 84 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_22
timestamp 1745462530
transform 1 0 1660 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_23
timestamp 1745462530
transform 1 0 1540 0 1 3315
box -2 -2 2 2
use M2_M1  M2_M1_24
timestamp 1745462530
transform 1 0 1508 0 1 3315
box -2 -2 2 2
use M2_M1  M2_M1_25
timestamp 1745462530
transform 1 0 1508 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_26
timestamp 1745462530
transform 1 0 1492 0 1 3315
box -2 -2 2 2
use M2_M1  M2_M1_27
timestamp 1745462530
transform 1 0 1492 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_28
timestamp 1745462530
transform 1 0 1444 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_29
timestamp 1745462530
transform 1 0 1364 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_30
timestamp 1745462530
transform 1 0 1276 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_31
timestamp 1745462530
transform 1 0 1580 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_32
timestamp 1745462530
transform 1 0 1532 0 1 3305
box -2 -2 2 2
use M2_M1  M2_M1_33
timestamp 1745462530
transform 1 0 1500 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_34
timestamp 1745462530
transform 1 0 1492 0 1 3305
box -2 -2 2 2
use M2_M1  M2_M1_35
timestamp 1745462530
transform 1 0 1484 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_36
timestamp 1745462530
transform 1 0 1460 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_37
timestamp 1745462530
transform 1 0 1436 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_38
timestamp 1745462530
transform 1 0 1996 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_39
timestamp 1745462530
transform 1 0 1948 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_40
timestamp 1745462530
transform 1 0 1924 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_41
timestamp 1745462530
transform 1 0 1716 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_42
timestamp 1745462530
transform 1 0 1700 0 1 3105
box -2 -2 2 2
use M2_M1  M2_M1_43
timestamp 1745462530
transform 1 0 1548 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_44
timestamp 1745462530
transform 1 0 1508 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_45
timestamp 1745462530
transform 1 0 1436 0 1 3315
box -2 -2 2 2
use M2_M1  M2_M1_46
timestamp 1745462530
transform 1 0 1684 0 1 3625
box -2 -2 2 2
use M2_M1  M2_M1_47
timestamp 1745462530
transform 1 0 1644 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_48
timestamp 1745462530
transform 1 0 1644 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_49
timestamp 1745462530
transform 1 0 1572 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_50
timestamp 1745462530
transform 1 0 1556 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_51
timestamp 1745462530
transform 1 0 1548 0 1 3625
box -2 -2 2 2
use M2_M1  M2_M1_52
timestamp 1745462530
transform 1 0 1492 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_53
timestamp 1745462530
transform 1 0 1372 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_54
timestamp 1745462530
transform 1 0 1372 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_55
timestamp 1745462530
transform 1 0 1692 0 1 3635
box -2 -2 2 2
use M2_M1  M2_M1_56
timestamp 1745462530
transform 1 0 1628 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_57
timestamp 1745462530
transform 1 0 1540 0 1 3645
box -2 -2 2 2
use M2_M1  M2_M1_58
timestamp 1745462530
transform 1 0 1404 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_59
timestamp 1745462530
transform 1 0 1388 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_60
timestamp 1745462530
transform 1 0 1244 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_61
timestamp 1745462530
transform 1 0 1244 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_62
timestamp 1745462530
transform 1 0 1996 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_63
timestamp 1745462530
transform 1 0 1972 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_64
timestamp 1745462530
transform 1 0 1940 0 1 3715
box -2 -2 2 2
use M2_M1  M2_M1_65
timestamp 1745462530
transform 1 0 1900 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_66
timestamp 1745462530
transform 1 0 1892 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_67
timestamp 1745462530
transform 1 0 1852 0 1 3715
box -2 -2 2 2
use M2_M1  M2_M1_68
timestamp 1745462530
transform 1 0 1804 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_69
timestamp 1745462530
transform 1 0 1700 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_70
timestamp 1745462530
transform 1 0 1676 0 1 3705
box -2 -2 2 2
use M2_M1  M2_M1_71
timestamp 1745462530
transform 1 0 1612 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_72
timestamp 1745462530
transform 1 0 1156 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_73
timestamp 1745462530
transform 1 0 940 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_74
timestamp 1745462530
transform 1 0 1084 0 1 3545
box -2 -2 2 2
use M2_M1  M2_M1_75
timestamp 1745462530
transform 1 0 836 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_76
timestamp 1745462530
transform 1 0 3124 0 1 3315
box -2 -2 2 2
use M2_M1  M2_M1_77
timestamp 1745462530
transform 1 0 3044 0 1 3225
box -2 -2 2 2
use M2_M1  M2_M1_78
timestamp 1745462530
transform 1 0 3036 0 1 3305
box -2 -2 2 2
use M2_M1  M2_M1_79
timestamp 1745462530
transform 1 0 2972 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_80
timestamp 1745462530
transform 1 0 2324 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_81
timestamp 1745462530
transform 1 0 868 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_82
timestamp 1745462530
transform 1 0 596 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_83
timestamp 1745462530
transform 1 0 3172 0 1 3235
box -2 -2 2 2
use M2_M1  M2_M1_84
timestamp 1745462530
transform 1 0 3132 0 1 3305
box -2 -2 2 2
use M2_M1  M2_M1_85
timestamp 1745462530
transform 1 0 3028 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_86
timestamp 1745462530
transform 1 0 2932 0 1 3225
box -2 -2 2 2
use M2_M1  M2_M1_87
timestamp 1745462530
transform 1 0 2316 0 1 3225
box -2 -2 2 2
use M2_M1  M2_M1_88
timestamp 1745462530
transform 1 0 996 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_89
timestamp 1745462530
transform 1 0 700 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_90
timestamp 1745462530
transform 1 0 3100 0 1 3235
box -2 -2 2 2
use M2_M1  M2_M1_91
timestamp 1745462530
transform 1 0 3068 0 1 3235
box -2 -2 2 2
use M2_M1  M2_M1_92
timestamp 1745462530
transform 1 0 3052 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_93
timestamp 1745462530
transform 1 0 2948 0 1 3235
box -2 -2 2 2
use M2_M1  M2_M1_94
timestamp 1745462530
transform 1 0 2916 0 1 3235
box -2 -2 2 2
use M2_M1  M2_M1_95
timestamp 1745462530
transform 1 0 2332 0 1 3235
box -2 -2 2 2
use M2_M1  M2_M1_96
timestamp 1745462530
transform 1 0 2292 0 1 3235
box -2 -2 2 2
use M2_M1  M2_M1_97
timestamp 1745462530
transform 1 0 924 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_98
timestamp 1745462530
transform 1 0 588 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_99
timestamp 1745462530
transform 1 0 2132 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_100
timestamp 1745462530
transform 1 0 2108 0 1 3345
box -2 -2 2 2
use M2_M1  M2_M1_101
timestamp 1745462530
transform 1 0 2076 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_102
timestamp 1745462530
transform 1 0 2052 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_103
timestamp 1745462530
transform 1 0 876 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_104
timestamp 1745462530
transform 1 0 676 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_105
timestamp 1745462530
transform 1 0 2284 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_106
timestamp 1745462530
transform 1 0 2236 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_107
timestamp 1745462530
transform 1 0 2124 0 1 3515
box -2 -2 2 2
use M2_M1  M2_M1_108
timestamp 1745462530
transform 1 0 2084 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_109
timestamp 1745462530
transform 1 0 2068 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_110
timestamp 1745462530
transform 1 0 2012 0 1 3345
box -2 -2 2 2
use M2_M1  M2_M1_111
timestamp 1745462530
transform 1 0 932 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_112
timestamp 1745462530
transform 1 0 716 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_113
timestamp 1745462530
transform 1 0 2276 0 1 3315
box -2 -2 2 2
use M2_M1  M2_M1_114
timestamp 1745462530
transform 1 0 2228 0 1 3315
box -2 -2 2 2
use M2_M1  M2_M1_115
timestamp 1745462530
transform 1 0 2180 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_116
timestamp 1745462530
transform 1 0 2084 0 1 3545
box -2 -2 2 2
use M2_M1  M2_M1_117
timestamp 1745462530
transform 1 0 2060 0 1 3315
box -2 -2 2 2
use M2_M1  M2_M1_118
timestamp 1745462530
transform 1 0 1148 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_119
timestamp 1745462530
transform 1 0 540 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_120
timestamp 1745462530
transform 1 0 1700 0 1 3315
box -2 -2 2 2
use M2_M1  M2_M1_121
timestamp 1745462530
transform 1 0 1684 0 1 3305
box -2 -2 2 2
use M2_M1  M2_M1_122
timestamp 1745462530
transform 1 0 1652 0 1 3425
box -2 -2 2 2
use M2_M1  M2_M1_123
timestamp 1745462530
transform 1 0 1644 0 1 3305
box -2 -2 2 2
use M2_M1  M2_M1_124
timestamp 1745462530
transform 1 0 1572 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_125
timestamp 1745462530
transform 1 0 1252 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_126
timestamp 1745462530
transform 1 0 1156 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_127
timestamp 1745462530
transform 1 0 1764 0 1 3235
box -2 -2 2 2
use M2_M1  M2_M1_128
timestamp 1745462530
transform 1 0 1708 0 1 3305
box -2 -2 2 2
use M2_M1  M2_M1_129
timestamp 1745462530
transform 1 0 1668 0 1 3435
box -2 -2 2 2
use M2_M1  M2_M1_130
timestamp 1745462530
transform 1 0 1636 0 1 3235
box -2 -2 2 2
use M2_M1  M2_M1_131
timestamp 1745462530
transform 1 0 1372 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_132
timestamp 1745462530
transform 1 0 1300 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_133
timestamp 1745462530
transform 1 0 1284 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_134
timestamp 1745462530
transform 1 0 1700 0 1 3235
box -2 -2 2 2
use M2_M1  M2_M1_135
timestamp 1745462530
transform 1 0 1668 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_136
timestamp 1745462530
transform 1 0 1652 0 1 3225
box -2 -2 2 2
use M2_M1  M2_M1_137
timestamp 1745462530
transform 1 0 1636 0 1 3315
box -2 -2 2 2
use M2_M1  M2_M1_138
timestamp 1745462530
transform 1 0 1596 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_139
timestamp 1745462530
transform 1 0 1260 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_140
timestamp 1745462530
transform 1 0 1052 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_141
timestamp 1745462530
transform 1 0 1788 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_142
timestamp 1745462530
transform 1 0 1772 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_143
timestamp 1745462530
transform 1 0 1732 0 1 3625
box -2 -2 2 2
use M2_M1  M2_M1_144
timestamp 1745462530
transform 1 0 1732 0 1 3425
box -2 -2 2 2
use M2_M1  M2_M1_145
timestamp 1745462530
transform 1 0 1652 0 1 3545
box -2 -2 2 2
use M2_M1  M2_M1_146
timestamp 1745462530
transform 1 0 1388 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_147
timestamp 1745462530
transform 1 0 1356 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_148
timestamp 1745462530
transform 1 0 1028 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_149
timestamp 1745462530
transform 1 0 1612 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_150
timestamp 1745462530
transform 1 0 1268 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_151
timestamp 1745462530
transform 1 0 1244 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_152
timestamp 1745462530
transform 1 0 1124 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_153
timestamp 1745462530
transform 1 0 1876 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_154
timestamp 1745462530
transform 1 0 1828 0 1 3435
box -2 -2 2 2
use M2_M1  M2_M1_155
timestamp 1745462530
transform 1 0 1788 0 1 3425
box -2 -2 2 2
use M2_M1  M2_M1_156
timestamp 1745462530
transform 1 0 1740 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_157
timestamp 1745462530
transform 1 0 1636 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_158
timestamp 1745462530
transform 1 0 1276 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_159
timestamp 1745462530
transform 1 0 876 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_160
timestamp 1745462530
transform 1 0 772 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_161
timestamp 1745462530
transform 1 0 732 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_162
timestamp 1745462530
transform 1 0 492 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_163
timestamp 1745462530
transform 1 0 692 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_164
timestamp 1745462530
transform 1 0 660 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_165
timestamp 1745462530
transform 1 0 588 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_166
timestamp 1745462530
transform 1 0 564 0 1 3145
box -2 -2 2 2
use M2_M1  M2_M1_167
timestamp 1745462530
transform 1 0 484 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_168
timestamp 1745462530
transform 1 0 620 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_169
timestamp 1745462530
transform 1 0 524 0 1 2995
box -2 -2 2 2
use M2_M1  M2_M1_170
timestamp 1745462530
transform 1 0 476 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_171
timestamp 1745462530
transform 1 0 476 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_172
timestamp 1745462530
transform 1 0 396 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_173
timestamp 1745462530
transform 1 0 516 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_174
timestamp 1745462530
transform 1 0 420 0 1 2995
box -2 -2 2 2
use M2_M1  M2_M1_175
timestamp 1745462530
transform 1 0 380 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_176
timestamp 1745462530
transform 1 0 364 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_177
timestamp 1745462530
transform 1 0 284 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_178
timestamp 1745462530
transform 1 0 412 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_179
timestamp 1745462530
transform 1 0 308 0 1 2995
box -2 -2 2 2
use M2_M1  M2_M1_180
timestamp 1745462530
transform 1 0 268 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_181
timestamp 1745462530
transform 1 0 180 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_182
timestamp 1745462530
transform 1 0 156 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_183
timestamp 1745462530
transform 1 0 268 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_184
timestamp 1745462530
transform 1 0 228 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_185
timestamp 1745462530
transform 1 0 172 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_186
timestamp 1745462530
transform 1 0 148 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_187
timestamp 1745462530
transform 1 0 2508 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_188
timestamp 1745462530
transform 1 0 2476 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_189
timestamp 1745462530
transform 1 0 2452 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_190
timestamp 1745462530
transform 1 0 2436 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_191
timestamp 1745462530
transform 1 0 2364 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_192
timestamp 1745462530
transform 1 0 2356 0 1 2305
box -2 -2 2 2
use M2_M1  M2_M1_193
timestamp 1745462530
transform 1 0 2348 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_194
timestamp 1745462530
transform 1 0 2348 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_195
timestamp 1745462530
transform 1 0 2324 0 1 2505
box -2 -2 2 2
use M2_M1  M2_M1_196
timestamp 1745462530
transform 1 0 2300 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_197
timestamp 1745462530
transform 1 0 2444 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_198
timestamp 1745462530
transform 1 0 2380 0 1 2435
box -2 -2 2 2
use M2_M1  M2_M1_199
timestamp 1745462530
transform 1 0 2356 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_200
timestamp 1745462530
transform 1 0 2340 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_201
timestamp 1745462530
transform 1 0 2332 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_202
timestamp 1745462530
transform 1 0 2316 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_203
timestamp 1745462530
transform 1 0 2308 0 1 2505
box -2 -2 2 2
use M2_M1  M2_M1_204
timestamp 1745462530
transform 1 0 2292 0 1 2505
box -2 -2 2 2
use M2_M1  M2_M1_205
timestamp 1745462530
transform 1 0 2284 0 1 2235
box -2 -2 2 2
use M2_M1  M2_M1_206
timestamp 1745462530
transform 1 0 2276 0 1 2505
box -2 -2 2 2
use M2_M1  M2_M1_207
timestamp 1745462530
transform 1 0 2372 0 1 2305
box -2 -2 2 2
use M2_M1  M2_M1_208
timestamp 1745462530
transform 1 0 2364 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_209
timestamp 1745462530
transform 1 0 2348 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_210
timestamp 1745462530
transform 1 0 2332 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_211
timestamp 1745462530
transform 1 0 2316 0 1 2305
box -2 -2 2 2
use M2_M1  M2_M1_212
timestamp 1745462530
transform 1 0 2300 0 1 2745
box -2 -2 2 2
use M2_M1  M2_M1_213
timestamp 1745462530
transform 1 0 2300 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_214
timestamp 1745462530
transform 1 0 2292 0 1 2435
box -2 -2 2 2
use M2_M1  M2_M1_215
timestamp 1745462530
transform 1 0 2292 0 1 2235
box -2 -2 2 2
use M2_M1  M2_M1_216
timestamp 1745462530
transform 1 0 2276 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_217
timestamp 1745462530
transform 1 0 2252 0 1 2555
box -2 -2 2 2
use M2_M1  M2_M1_218
timestamp 1745462530
transform 1 0 2244 0 1 2545
box -2 -2 2 2
use M2_M1  M2_M1_219
timestamp 1745462530
transform 1 0 2244 0 1 2305
box -2 -2 2 2
use M2_M1  M2_M1_220
timestamp 1745462530
transform 1 0 2228 0 1 2745
box -2 -2 2 2
use M2_M1  M2_M1_221
timestamp 1745462530
transform 1 0 2220 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_222
timestamp 1745462530
transform 1 0 2212 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_223
timestamp 1745462530
transform 1 0 2140 0 1 2235
box -2 -2 2 2
use M2_M1  M2_M1_224
timestamp 1745462530
transform 1 0 2092 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_225
timestamp 1745462530
transform 1 0 2276 0 1 2105
box -2 -2 2 2
use M2_M1  M2_M1_226
timestamp 1745462530
transform 1 0 2252 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_227
timestamp 1745462530
transform 1 0 2236 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_228
timestamp 1745462530
transform 1 0 2188 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_229
timestamp 1745462530
transform 1 0 2180 0 1 2545
box -2 -2 2 2
use M2_M1  M2_M1_230
timestamp 1745462530
transform 1 0 2140 0 1 2105
box -2 -2 2 2
use M2_M1  M2_M1_231
timestamp 1745462530
transform 1 0 2108 0 1 2105
box -2 -2 2 2
use M2_M1  M2_M1_232
timestamp 1745462530
transform 1 0 2100 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_233
timestamp 1745462530
transform 1 0 2076 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_234
timestamp 1745462530
transform 1 0 2300 0 1 2105
box -2 -2 2 2
use M2_M1  M2_M1_235
timestamp 1745462530
transform 1 0 2276 0 1 2305
box -2 -2 2 2
use M2_M1  M2_M1_236
timestamp 1745462530
transform 1 0 2228 0 1 2105
box -2 -2 2 2
use M2_M1  M2_M1_237
timestamp 1745462530
transform 1 0 2196 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_238
timestamp 1745462530
transform 1 0 2188 0 1 2745
box -2 -2 2 2
use M2_M1  M2_M1_239
timestamp 1745462530
transform 1 0 2188 0 1 2105
box -2 -2 2 2
use M2_M1  M2_M1_240
timestamp 1745462530
transform 1 0 2180 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_241
timestamp 1745462530
transform 1 0 2108 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_242
timestamp 1745462530
transform 1 0 1004 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_243
timestamp 1745462530
transform 1 0 972 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_244
timestamp 1745462530
transform 1 0 932 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_245
timestamp 1745462530
transform 1 0 1020 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_246
timestamp 1745462530
transform 1 0 996 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_247
timestamp 1745462530
transform 1 0 1180 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_248
timestamp 1745462530
transform 1 0 1132 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_249
timestamp 1745462530
transform 1 0 1116 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_250
timestamp 1745462530
transform 1 0 284 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_251
timestamp 1745462530
transform 1 0 244 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_252
timestamp 1745462530
transform 1 0 244 0 1 4025
box -2 -2 2 2
use M2_M1  M2_M1_253
timestamp 1745462530
transform 1 0 244 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_254
timestamp 1745462530
transform 1 0 676 0 1 4005
box -2 -2 2 2
use M2_M1  M2_M1_255
timestamp 1745462530
transform 1 0 676 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_256
timestamp 1745462530
transform 1 0 548 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_257
timestamp 1745462530
transform 1 0 548 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_258
timestamp 1745462530
transform 1 0 316 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_259
timestamp 1745462530
transform 1 0 292 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_260
timestamp 1745462530
transform 1 0 444 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_261
timestamp 1745462530
transform 1 0 404 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_262
timestamp 1745462530
transform 1 0 404 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_263
timestamp 1745462530
transform 1 0 364 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_264
timestamp 1745462530
transform 1 0 372 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_265
timestamp 1745462530
transform 1 0 300 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_266
timestamp 1745462530
transform 1 0 788 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_267
timestamp 1745462530
transform 1 0 732 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_268
timestamp 1745462530
transform 1 0 604 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_269
timestamp 1745462530
transform 1 0 780 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_270
timestamp 1745462530
transform 1 0 764 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_271
timestamp 1745462530
transform 1 0 668 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_272
timestamp 1745462530
transform 1 0 636 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_273
timestamp 1745462530
transform 1 0 2228 0 1 2625
box -2 -2 2 2
use M2_M1  M2_M1_274
timestamp 1745462530
transform 1 0 2204 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_275
timestamp 1745462530
transform 1 0 2188 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_276
timestamp 1745462530
transform 1 0 2364 0 1 2595
box -2 -2 2 2
use M2_M1  M2_M1_277
timestamp 1745462530
transform 1 0 2284 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_278
timestamp 1745462530
transform 1 0 2196 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_279
timestamp 1745462530
transform 1 0 2180 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_280
timestamp 1745462530
transform 1 0 2436 0 1 2545
box -2 -2 2 2
use M2_M1  M2_M1_281
timestamp 1745462530
transform 1 0 2372 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_282
timestamp 1745462530
transform 1 0 2364 0 1 2545
box -2 -2 2 2
use M2_M1  M2_M1_283
timestamp 1745462530
transform 1 0 2300 0 1 2635
box -2 -2 2 2
use M2_M1  M2_M1_284
timestamp 1745462530
transform 1 0 2276 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_285
timestamp 1745462530
transform 1 0 2292 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_286
timestamp 1745462530
transform 1 0 2268 0 1 2715
box -2 -2 2 2
use M2_M1  M2_M1_287
timestamp 1745462530
transform 1 0 2244 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_288
timestamp 1745462530
transform 1 0 2228 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_289
timestamp 1745462530
transform 1 0 396 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_290
timestamp 1745462530
transform 1 0 372 0 1 3515
box -2 -2 2 2
use M2_M1  M2_M1_291
timestamp 1745462530
transform 1 0 300 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_292
timestamp 1745462530
transform 1 0 268 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_293
timestamp 1745462530
transform 1 0 316 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_294
timestamp 1745462530
transform 1 0 236 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_295
timestamp 1745462530
transform 1 0 228 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_296
timestamp 1745462530
transform 1 0 204 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_297
timestamp 1745462530
transform 1 0 188 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_298
timestamp 1745462530
transform 1 0 172 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_299
timestamp 1745462530
transform 1 0 420 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_300
timestamp 1745462530
transform 1 0 396 0 1 3515
box -2 -2 2 2
use M2_M1  M2_M1_301
timestamp 1745462530
transform 1 0 268 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_302
timestamp 1745462530
transform 1 0 244 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_303
timestamp 1745462530
transform 1 0 356 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_304
timestamp 1745462530
transform 1 0 292 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_305
timestamp 1745462530
transform 1 0 212 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_306
timestamp 1745462530
transform 1 0 196 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_307
timestamp 1745462530
transform 1 0 212 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_308
timestamp 1745462530
transform 1 0 188 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_309
timestamp 1745462530
transform 1 0 132 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_310
timestamp 1745462530
transform 1 0 1588 0 1 3025
box -2 -2 2 2
use M2_M1  M2_M1_311
timestamp 1745462530
transform 1 0 1196 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_312
timestamp 1745462530
transform 1 0 1116 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_313
timestamp 1745462530
transform 1 0 1092 0 1 3225
box -2 -2 2 2
use M2_M1  M2_M1_314
timestamp 1745462530
transform 1 0 2188 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_315
timestamp 1745462530
transform 1 0 2188 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_316
timestamp 1745462530
transform 1 0 2188 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_317
timestamp 1745462530
transform 1 0 2140 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_318
timestamp 1745462530
transform 1 0 2124 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_319
timestamp 1745462530
transform 1 0 2084 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_320
timestamp 1745462530
transform 1 0 2084 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_321
timestamp 1745462530
transform 1 0 1020 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_322
timestamp 1745462530
transform 1 0 988 0 1 3235
box -2 -2 2 2
use M2_M1  M2_M1_323
timestamp 1745462530
transform 1 0 972 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_324
timestamp 1745462530
transform 1 0 2340 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_325
timestamp 1745462530
transform 1 0 2276 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_326
timestamp 1745462530
transform 1 0 2228 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_327
timestamp 1745462530
transform 1 0 2204 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_328
timestamp 1745462530
transform 1 0 2316 0 1 3315
box -2 -2 2 2
use M2_M1  M2_M1_329
timestamp 1745462530
transform 1 0 2268 0 1 3425
box -2 -2 2 2
use M2_M1  M2_M1_330
timestamp 1745462530
transform 1 0 2204 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_331
timestamp 1745462530
transform 1 0 2124 0 1 3435
box -2 -2 2 2
use M2_M1  M2_M1_332
timestamp 1745462530
transform 1 0 2100 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_333
timestamp 1745462530
transform 1 0 2228 0 1 3425
box -2 -2 2 2
use M2_M1  M2_M1_334
timestamp 1745462530
transform 1 0 2140 0 1 3425
box -2 -2 2 2
use M2_M1  M2_M1_335
timestamp 1745462530
transform 1 0 2084 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_336
timestamp 1745462530
transform 1 0 3140 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_337
timestamp 1745462530
transform 1 0 3140 0 1 3235
box -2 -2 2 2
use M2_M1  M2_M1_338
timestamp 1745462530
transform 1 0 3052 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_339
timestamp 1745462530
transform 1 0 3028 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_340
timestamp 1745462530
transform 1 0 3004 0 1 3305
box -2 -2 2 2
use M2_M1  M2_M1_341
timestamp 1745462530
transform 1 0 3004 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_342
timestamp 1745462530
transform 1 0 3108 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_343
timestamp 1745462530
transform 1 0 3076 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_344
timestamp 1745462530
transform 1 0 3060 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_345
timestamp 1745462530
transform 1 0 3028 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_346
timestamp 1745462530
transform 1 0 3012 0 1 3315
box -2 -2 2 2
use M2_M1  M2_M1_347
timestamp 1745462530
transform 1 0 3004 0 1 3225
box -2 -2 2 2
use M2_M1  M2_M1_348
timestamp 1745462530
transform 1 0 3132 0 1 3225
box -2 -2 2 2
use M2_M1  M2_M1_349
timestamp 1745462530
transform 1 0 3108 0 1 3225
box -2 -2 2 2
use M2_M1  M2_M1_350
timestamp 1745462530
transform 1 0 3004 0 1 3235
box -2 -2 2 2
use M2_M1  M2_M1_351
timestamp 1745462530
transform 1 0 2964 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_352
timestamp 1745462530
transform 1 0 2940 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_353
timestamp 1745462530
transform 1 0 1684 0 1 3115
box -2 -2 2 2
use M2_M1  M2_M1_354
timestamp 1745462530
transform 1 0 1604 0 1 3224
box -2 -2 2 2
use M2_M1  M2_M1_355
timestamp 1745462530
transform 1 0 1540 0 1 3235
box -2 -2 2 2
use M2_M1  M2_M1_356
timestamp 1745462530
transform 1 0 1516 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_357
timestamp 1745462530
transform 1 0 1492 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_358
timestamp 1745462530
transform 1 0 1380 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_359
timestamp 1745462530
transform 1 0 1324 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_360
timestamp 1745462530
transform 1 0 1300 0 1 3155
box -2 -2 2 2
use M2_M1  M2_M1_361
timestamp 1745462530
transform 1 0 1300 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_362
timestamp 1745462530
transform 1 0 1772 0 1 3225
box -2 -2 2 2
use M2_M1  M2_M1_363
timestamp 1745462530
transform 1 0 1732 0 1 3235
box -2 -2 2 2
use M2_M1  M2_M1_364
timestamp 1745462530
transform 1 0 1684 0 1 3235
box -2 -2 2 2
use M2_M1  M2_M1_365
timestamp 1745462530
transform 1 0 1660 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_366
timestamp 1745462530
transform 1 0 1572 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_367
timestamp 1745462530
transform 1 0 1340 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_368
timestamp 1745462530
transform 1 0 1332 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_369
timestamp 1745462530
transform 1 0 1860 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_370
timestamp 1745462530
transform 1 0 1828 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_371
timestamp 1745462530
transform 1 0 1748 0 1 3545
box -2 -2 2 2
use M2_M1  M2_M1_372
timestamp 1745462530
transform 1 0 1740 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_373
timestamp 1745462530
transform 1 0 1708 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_374
timestamp 1745462530
transform 1 0 1676 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_375
timestamp 1745462530
transform 1 0 1644 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_376
timestamp 1745462530
transform 1 0 1644 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_377
timestamp 1745462530
transform 1 0 1260 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_378
timestamp 1745462530
transform 1 0 724 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_379
timestamp 1745462530
transform 1 0 708 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_380
timestamp 1745462530
transform 1 0 676 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_381
timestamp 1745462530
transform 1 0 652 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_382
timestamp 1745462530
transform 1 0 2188 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_383
timestamp 1745462530
transform 1 0 2172 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_384
timestamp 1745462530
transform 1 0 2164 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_385
timestamp 1745462530
transform 1 0 2164 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_386
timestamp 1745462530
transform 1 0 2148 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_387
timestamp 1745462530
transform 1 0 2100 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_388
timestamp 1745462530
transform 1 0 2100 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_389
timestamp 1745462530
transform 1 0 2444 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_390
timestamp 1745462530
transform 1 0 2404 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_391
timestamp 1745462530
transform 1 0 2372 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_392
timestamp 1745462530
transform 1 0 2372 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_393
timestamp 1745462530
transform 1 0 2348 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_394
timestamp 1745462530
transform 1 0 2332 0 1 2625
box -2 -2 2 2
use M2_M1  M2_M1_395
timestamp 1745462530
transform 1 0 2316 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_396
timestamp 1745462530
transform 1 0 2300 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_397
timestamp 1745462530
transform 1 0 2284 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_398
timestamp 1745462530
transform 1 0 2276 0 1 2435
box -2 -2 2 2
use M2_M1  M2_M1_399
timestamp 1745462530
transform 1 0 2268 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_400
timestamp 1745462530
transform 1 0 2236 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_401
timestamp 1745462530
transform 1 0 2236 0 1 2515
box -2 -2 2 2
use M2_M1  M2_M1_402
timestamp 1745462530
transform 1 0 2212 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_403
timestamp 1745462530
transform 1 0 2068 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_404
timestamp 1745462530
transform 1 0 2324 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_405
timestamp 1745462530
transform 1 0 2316 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_406
timestamp 1745462530
transform 1 0 2308 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_407
timestamp 1745462530
transform 1 0 2308 0 1 2625
box -2 -2 2 2
use M2_M1  M2_M1_408
timestamp 1745462530
transform 1 0 2308 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_409
timestamp 1745462530
transform 1 0 2292 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_410
timestamp 1745462530
transform 1 0 2292 0 1 2515
box -2 -2 2 2
use M2_M1  M2_M1_411
timestamp 1745462530
transform 1 0 2252 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_412
timestamp 1745462530
transform 1 0 2252 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_413
timestamp 1745462530
transform 1 0 2244 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_414
timestamp 1745462530
transform 1 0 2244 0 1 2555
box -2 -2 2 2
use M2_M1  M2_M1_415
timestamp 1745462530
transform 1 0 2484 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_416
timestamp 1745462530
transform 1 0 2412 0 1 2545
box -2 -2 2 2
use M2_M1  M2_M1_417
timestamp 1745462530
transform 1 0 2660 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_418
timestamp 1745462530
transform 1 0 2252 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_419
timestamp 1745462530
transform 1 0 2228 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_420
timestamp 1745462530
transform 1 0 2132 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_421
timestamp 1745462530
transform 1 0 2604 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_422
timestamp 1745462530
transform 1 0 2220 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_423
timestamp 1745462530
transform 1 0 2092 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_424
timestamp 1745462530
transform 1 0 3364 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_425
timestamp 1745462530
transform 1 0 3324 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_426
timestamp 1745462530
transform 1 0 2596 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_427
timestamp 1745462530
transform 1 0 2564 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_428
timestamp 1745462530
transform 1 0 1532 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_429
timestamp 1745462530
transform 1 0 860 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_430
timestamp 1745462530
transform 1 0 836 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_431
timestamp 1745462530
transform 1 0 2356 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_432
timestamp 1745462530
transform 1 0 2340 0 1 2435
box -2 -2 2 2
use M2_M1  M2_M1_433
timestamp 1745462530
transform 1 0 2316 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_434
timestamp 1745462530
transform 1 0 2260 0 1 2505
box -2 -2 2 2
use M2_M1  M2_M1_435
timestamp 1745462530
transform 1 0 2260 0 1 2435
box -2 -2 2 2
use M2_M1  M2_M1_436
timestamp 1745462530
transform 1 0 2228 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_437
timestamp 1745462530
transform 1 0 3324 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_438
timestamp 1745462530
transform 1 0 3292 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_439
timestamp 1745462530
transform 1 0 2636 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_440
timestamp 1745462530
transform 1 0 2540 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_441
timestamp 1745462530
transform 1 0 1596 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_442
timestamp 1745462530
transform 1 0 948 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_443
timestamp 1745462530
transform 1 0 932 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_444
timestamp 1745462530
transform 1 0 3324 0 1 1315
box -2 -2 2 2
use M2_M1  M2_M1_445
timestamp 1745462530
transform 1 0 3236 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_446
timestamp 1745462530
transform 1 0 2676 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_447
timestamp 1745462530
transform 1 0 2220 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_448
timestamp 1745462530
transform 1 0 1596 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_449
timestamp 1745462530
transform 1 0 892 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_450
timestamp 1745462530
transform 1 0 868 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_451
timestamp 1745462530
transform 1 0 3276 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_452
timestamp 1745462530
transform 1 0 3252 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_453
timestamp 1745462530
transform 1 0 2676 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_454
timestamp 1745462530
transform 1 0 2636 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_455
timestamp 1745462530
transform 1 0 2452 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_456
timestamp 1745462530
transform 1 0 2444 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_457
timestamp 1745462530
transform 1 0 1564 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_458
timestamp 1745462530
transform 1 0 932 0 1 2515
box -2 -2 2 2
use M2_M1  M2_M1_459
timestamp 1745462530
transform 1 0 932 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_460
timestamp 1745462530
transform 1 0 1308 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_461
timestamp 1745462530
transform 1 0 1076 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_462
timestamp 1745462530
transform 1 0 1044 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_463
timestamp 1745462530
transform 1 0 1028 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_464
timestamp 1745462530
transform 1 0 2452 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_465
timestamp 1745462530
transform 1 0 2436 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_466
timestamp 1745462530
transform 1 0 2396 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_467
timestamp 1745462530
transform 1 0 2172 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_468
timestamp 1745462530
transform 1 0 2292 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_469
timestamp 1745462530
transform 1 0 2212 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_470
timestamp 1745462530
transform 1 0 2204 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_471
timestamp 1745462530
transform 1 0 2196 0 1 2625
box -2 -2 2 2
use M2_M1  M2_M1_472
timestamp 1745462530
transform 1 0 2180 0 1 2305
box -2 -2 2 2
use M2_M1  M2_M1_473
timestamp 1745462530
transform 1 0 2180 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_474
timestamp 1745462530
transform 1 0 2148 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_475
timestamp 1745462530
transform 1 0 2140 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_476
timestamp 1745462530
transform 1 0 2508 0 1 1795
box -2 -2 2 2
use M2_M1  M2_M1_477
timestamp 1745462530
transform 1 0 2508 0 1 1745
box -2 -2 2 2
use M2_M1  M2_M1_478
timestamp 1745462530
transform 1 0 2492 0 1 1795
box -2 -2 2 2
use M2_M1  M2_M1_479
timestamp 1745462530
transform 1 0 2484 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_480
timestamp 1745462530
transform 1 0 2460 0 1 1745
box -2 -2 2 2
use M2_M1  M2_M1_481
timestamp 1745462530
transform 1 0 2388 0 1 1795
box -2 -2 2 2
use M2_M1  M2_M1_482
timestamp 1745462530
transform 1 0 2372 0 1 1745
box -2 -2 2 2
use M2_M1  M2_M1_483
timestamp 1745462530
transform 1 0 2324 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_484
timestamp 1745462530
transform 1 0 2324 0 1 1745
box -2 -2 2 2
use M2_M1  M2_M1_485
timestamp 1745462530
transform 1 0 1004 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_486
timestamp 1745462530
transform 1 0 932 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_487
timestamp 1745462530
transform 1 0 908 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_488
timestamp 1745462530
transform 1 0 868 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_489
timestamp 1745462530
transform 1 0 852 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_490
timestamp 1745462530
transform 1 0 812 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_491
timestamp 1745462530
transform 1 0 1572 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_492
timestamp 1745462530
transform 1 0 1572 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_493
timestamp 1745462530
transform 1 0 1540 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_494
timestamp 1745462530
transform 1 0 1532 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_495
timestamp 1745462530
transform 1 0 1516 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_496
timestamp 1745462530
transform 1 0 3324 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_497
timestamp 1745462530
transform 1 0 3308 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_498
timestamp 1745462530
transform 1 0 3276 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_499
timestamp 1745462530
transform 1 0 3276 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_500
timestamp 1745462530
transform 1 0 3244 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_501
timestamp 1745462530
transform 1 0 3244 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_502
timestamp 1745462530
transform 1 0 2604 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_503
timestamp 1745462530
transform 1 0 2588 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_504
timestamp 1745462530
transform 1 0 2260 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_505
timestamp 1745462530
transform 1 0 2244 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_506
timestamp 1745462530
transform 1 0 2236 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_507
timestamp 1745462530
transform 1 0 2196 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_508
timestamp 1745462530
transform 1 0 2164 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_509
timestamp 1745462530
transform 1 0 2164 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_510
timestamp 1745462530
transform 1 0 2044 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_511
timestamp 1745462530
transform 1 0 3292 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_512
timestamp 1745462530
transform 1 0 3276 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_513
timestamp 1745462530
transform 1 0 3260 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_514
timestamp 1745462530
transform 1 0 3252 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_515
timestamp 1745462530
transform 1 0 3220 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_516
timestamp 1745462530
transform 1 0 3196 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_517
timestamp 1745462530
transform 1 0 1044 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_518
timestamp 1745462530
transform 1 0 996 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_519
timestamp 1745462530
transform 1 0 916 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_520
timestamp 1745462530
transform 1 0 916 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_521
timestamp 1745462530
transform 1 0 860 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_522
timestamp 1745462530
transform 1 0 844 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_523
timestamp 1745462530
transform 1 0 2676 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_524
timestamp 1745462530
transform 1 0 2652 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_525
timestamp 1745462530
transform 1 0 2652 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_526
timestamp 1745462530
transform 1 0 2636 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_527
timestamp 1745462530
transform 1 0 2596 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_528
timestamp 1745462530
transform 1 0 2580 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_529
timestamp 1745462530
transform 1 0 2148 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_530
timestamp 1745462530
transform 1 0 2132 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_531
timestamp 1745462530
transform 1 0 2108 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_532
timestamp 1745462530
transform 1 0 1340 0 1 2395
box -2 -2 2 2
use M2_M1  M2_M1_533
timestamp 1745462530
transform 1 0 2188 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_534
timestamp 1745462530
transform 1 0 2188 0 1 1745
box -2 -2 2 2
use M2_M1  M2_M1_535
timestamp 1745462530
transform 1 0 2204 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_536
timestamp 1745462530
transform 1 0 2148 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_537
timestamp 1745462530
transform 1 0 2148 0 1 1795
box -2 -2 2 2
use M2_M1  M2_M1_538
timestamp 1745462530
transform 1 0 1796 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_539
timestamp 1745462530
transform 1 0 1772 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_540
timestamp 1745462530
transform 1 0 1556 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_541
timestamp 1745462530
transform 1 0 1420 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_542
timestamp 1745462530
transform 1 0 1212 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_543
timestamp 1745462530
transform 1 0 1180 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_544
timestamp 1745462530
transform 1 0 1748 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_545
timestamp 1745462530
transform 1 0 1692 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_546
timestamp 1745462530
transform 1 0 1492 0 1 2515
box -2 -2 2 2
use M2_M1  M2_M1_547
timestamp 1745462530
transform 1 0 1436 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_548
timestamp 1745462530
transform 1 0 1412 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_549
timestamp 1745462530
transform 1 0 1292 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_550
timestamp 1745462530
transform 1 0 1228 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_551
timestamp 1745462530
transform 1 0 1180 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_552
timestamp 1745462530
transform 1 0 1764 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_553
timestamp 1745462530
transform 1 0 1716 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_554
timestamp 1745462530
transform 1 0 1540 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_555
timestamp 1745462530
transform 1 0 1492 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_556
timestamp 1745462530
transform 1 0 1340 0 1 1845
box -2 -2 2 2
use M2_M1  M2_M1_557
timestamp 1745462530
transform 1 0 1340 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_558
timestamp 1745462530
transform 1 0 1340 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_559
timestamp 1745462530
transform 1 0 1220 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_560
timestamp 1745462530
transform 1 0 1156 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_561
timestamp 1745462530
transform 1 0 812 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_562
timestamp 1745462530
transform 1 0 748 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_563
timestamp 1745462530
transform 1 0 420 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_564
timestamp 1745462530
transform 1 0 380 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_565
timestamp 1745462530
transform 1 0 364 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_566
timestamp 1745462530
transform 1 0 324 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_567
timestamp 1745462530
transform 1 0 260 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_568
timestamp 1745462530
transform 1 0 764 0 1 2655
box -2 -2 2 2
use M2_M1  M2_M1_569
timestamp 1745462530
transform 1 0 652 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_570
timestamp 1745462530
transform 1 0 564 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_571
timestamp 1745462530
transform 1 0 564 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_572
timestamp 1745462530
transform 1 0 516 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_573
timestamp 1745462530
transform 1 0 508 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_574
timestamp 1745462530
transform 1 0 428 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_575
timestamp 1745462530
transform 1 0 332 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_576
timestamp 1745462530
transform 1 0 252 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_577
timestamp 1745462530
transform 1 0 212 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_578
timestamp 1745462530
transform 1 0 212 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_579
timestamp 1745462530
transform 1 0 196 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_580
timestamp 1745462530
transform 1 0 940 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_581
timestamp 1745462530
transform 1 0 940 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_582
timestamp 1745462530
transform 1 0 932 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_583
timestamp 1745462530
transform 1 0 932 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_584
timestamp 1745462530
transform 1 0 916 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_585
timestamp 1745462530
transform 1 0 900 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_586
timestamp 1745462530
transform 1 0 380 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_587
timestamp 1745462530
transform 1 0 332 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_588
timestamp 1745462530
transform 1 0 324 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_589
timestamp 1745462530
transform 1 0 316 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_590
timestamp 1745462530
transform 1 0 244 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_591
timestamp 1745462530
transform 1 0 196 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_592
timestamp 1745462530
transform 1 0 196 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_593
timestamp 1745462530
transform 1 0 364 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_594
timestamp 1745462530
transform 1 0 364 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_595
timestamp 1745462530
transform 1 0 364 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_596
timestamp 1745462530
transform 1 0 204 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_597
timestamp 1745462530
transform 1 0 180 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_598
timestamp 1745462530
transform 1 0 180 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_599
timestamp 1745462530
transform 1 0 372 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_600
timestamp 1745462530
transform 1 0 284 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_601
timestamp 1745462530
transform 1 0 244 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_602
timestamp 1745462530
transform 1 0 220 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_603
timestamp 1745462530
transform 1 0 196 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_604
timestamp 1745462530
transform 1 0 196 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_605
timestamp 1745462530
transform 1 0 460 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_606
timestamp 1745462530
transform 1 0 460 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_607
timestamp 1745462530
transform 1 0 380 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_608
timestamp 1745462530
transform 1 0 292 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_609
timestamp 1745462530
transform 1 0 244 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_610
timestamp 1745462530
transform 1 0 188 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_611
timestamp 1745462530
transform 1 0 188 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_612
timestamp 1745462530
transform 1 0 700 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_613
timestamp 1745462530
transform 1 0 684 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_614
timestamp 1745462530
transform 1 0 684 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_615
timestamp 1745462530
transform 1 0 660 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_616
timestamp 1745462530
transform 1 0 628 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_617
timestamp 1745462530
transform 1 0 620 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_618
timestamp 1745462530
transform 1 0 532 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_619
timestamp 1745462530
transform 1 0 1892 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_620
timestamp 1745462530
transform 1 0 1804 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_621
timestamp 1745462530
transform 1 0 1668 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_622
timestamp 1745462530
transform 1 0 1468 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_623
timestamp 1745462530
transform 1 0 1388 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_624
timestamp 1745462530
transform 1 0 1124 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_625
timestamp 1745462530
transform 1 0 1020 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_626
timestamp 1745462530
transform 1 0 1876 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_627
timestamp 1745462530
transform 1 0 1764 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_628
timestamp 1745462530
transform 1 0 1652 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_629
timestamp 1745462530
transform 1 0 1540 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_630
timestamp 1745462530
transform 1 0 1436 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_631
timestamp 1745462530
transform 1 0 1340 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_632
timestamp 1745462530
transform 1 0 1316 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_633
timestamp 1745462530
transform 1 0 1868 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_634
timestamp 1745462530
transform 1 0 1812 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_635
timestamp 1745462530
transform 1 0 1708 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_636
timestamp 1745462530
transform 1 0 1604 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_637
timestamp 1745462530
transform 1 0 1380 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_638
timestamp 1745462530
transform 1 0 1324 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_639
timestamp 1745462530
transform 1 0 1244 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_640
timestamp 1745462530
transform 1 0 1884 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_641
timestamp 1745462530
transform 1 0 1876 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_642
timestamp 1745462530
transform 1 0 1700 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_643
timestamp 1745462530
transform 1 0 1532 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_644
timestamp 1745462530
transform 1 0 1468 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_645
timestamp 1745462530
transform 1 0 1404 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_646
timestamp 1745462530
transform 1 0 1300 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_647
timestamp 1745462530
transform 1 0 3068 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_648
timestamp 1745462530
transform 1 0 3020 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_649
timestamp 1745462530
transform 1 0 2716 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_650
timestamp 1745462530
transform 1 0 2268 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_651
timestamp 1745462530
transform 1 0 2188 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_652
timestamp 1745462530
transform 1 0 2188 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_653
timestamp 1745462530
transform 1 0 2772 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_654
timestamp 1745462530
transform 1 0 2676 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_655
timestamp 1745462530
transform 1 0 2660 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_656
timestamp 1745462530
transform 1 0 2580 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_657
timestamp 1745462530
transform 1 0 2508 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_658
timestamp 1745462530
transform 1 0 2284 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_659
timestamp 1745462530
transform 1 0 2220 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_660
timestamp 1745462530
transform 1 0 2972 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_661
timestamp 1745462530
transform 1 0 2900 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_662
timestamp 1745462530
transform 1 0 2764 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_663
timestamp 1745462530
transform 1 0 2700 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_664
timestamp 1745462530
transform 1 0 2268 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_665
timestamp 1745462530
transform 1 0 2268 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_666
timestamp 1745462530
transform 1 0 2228 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_667
timestamp 1745462530
transform 1 0 3068 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_668
timestamp 1745462530
transform 1 0 2996 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_669
timestamp 1745462530
transform 1 0 2940 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_670
timestamp 1745462530
transform 1 0 2644 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_671
timestamp 1745462530
transform 1 0 2596 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_672
timestamp 1745462530
transform 1 0 2492 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_673
timestamp 1745462530
transform 1 0 2436 0 1 345
box -2 -2 2 2
use M2_M1  M2_M1_674
timestamp 1745462530
transform 1 0 3844 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_675
timestamp 1745462530
transform 1 0 3796 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_676
timestamp 1745462530
transform 1 0 3796 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_677
timestamp 1745462530
transform 1 0 3708 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_678
timestamp 1745462530
transform 1 0 3508 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_679
timestamp 1745462530
transform 1 0 3500 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_680
timestamp 1745462530
transform 1 0 3348 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_681
timestamp 1745462530
transform 1 0 4212 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_682
timestamp 1745462530
transform 1 0 4212 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_683
timestamp 1745462530
transform 1 0 4124 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_684
timestamp 1745462530
transform 1 0 4068 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_685
timestamp 1745462530
transform 1 0 4044 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_686
timestamp 1745462530
transform 1 0 3988 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_687
timestamp 1745462530
transform 1 0 3740 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_688
timestamp 1745462530
transform 1 0 3956 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_689
timestamp 1745462530
transform 1 0 3948 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_690
timestamp 1745462530
transform 1 0 3748 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_691
timestamp 1745462530
transform 1 0 3716 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_692
timestamp 1745462530
transform 1 0 3636 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_693
timestamp 1745462530
transform 1 0 3484 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_694
timestamp 1745462530
transform 1 0 3364 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_695
timestamp 1745462530
transform 1 0 4308 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_696
timestamp 1745462530
transform 1 0 4252 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_697
timestamp 1745462530
transform 1 0 4204 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_698
timestamp 1745462530
transform 1 0 4140 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_699
timestamp 1745462530
transform 1 0 4124 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_700
timestamp 1745462530
transform 1 0 4084 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_701
timestamp 1745462530
transform 1 0 3804 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_702
timestamp 1745462530
transform 1 0 3796 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_703
timestamp 1745462530
transform 1 0 3676 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_704
timestamp 1745462530
transform 1 0 3660 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_705
timestamp 1745462530
transform 1 0 3660 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_706
timestamp 1745462530
transform 1 0 3660 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_707
timestamp 1745462530
transform 1 0 3500 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_708
timestamp 1745462530
transform 1 0 3468 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_709
timestamp 1745462530
transform 1 0 4212 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_710
timestamp 1745462530
transform 1 0 4204 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_711
timestamp 1745462530
transform 1 0 4204 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_712
timestamp 1745462530
transform 1 0 4188 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_713
timestamp 1745462530
transform 1 0 4172 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_714
timestamp 1745462530
transform 1 0 4148 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_715
timestamp 1745462530
transform 1 0 4108 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_716
timestamp 1745462530
transform 1 0 4052 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_717
timestamp 1745462530
transform 1 0 3844 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_718
timestamp 1745462530
transform 1 0 3844 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_719
timestamp 1745462530
transform 1 0 3796 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_720
timestamp 1745462530
transform 1 0 3772 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_721
timestamp 1745462530
transform 1 0 3676 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_722
timestamp 1745462530
transform 1 0 3636 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_723
timestamp 1745462530
transform 1 0 3564 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_724
timestamp 1745462530
transform 1 0 4300 0 1 1585
box -2 -2 2 2
use M2_M1  M2_M1_725
timestamp 1745462530
transform 1 0 4276 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_726
timestamp 1745462530
transform 1 0 4212 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_727
timestamp 1745462530
transform 1 0 4180 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_728
timestamp 1745462530
transform 1 0 4156 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_729
timestamp 1745462530
transform 1 0 4132 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_730
timestamp 1745462530
transform 1 0 3980 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_731
timestamp 1745462530
transform 1 0 4220 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_732
timestamp 1745462530
transform 1 0 4140 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_733
timestamp 1745462530
transform 1 0 3924 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_734
timestamp 1745462530
transform 1 0 3604 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_735
timestamp 1745462530
transform 1 0 3356 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_736
timestamp 1745462530
transform 1 0 3236 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_737
timestamp 1745462530
transform 1 0 4084 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_738
timestamp 1745462530
transform 1 0 4052 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_739
timestamp 1745462530
transform 1 0 3836 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_740
timestamp 1745462530
transform 1 0 3692 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_741
timestamp 1745462530
transform 1 0 3460 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_742
timestamp 1745462530
transform 1 0 3188 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_743
timestamp 1745462530
transform 1 0 3172 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_744
timestamp 1745462530
transform 1 0 1900 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_745
timestamp 1745462530
transform 1 0 1828 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_746
timestamp 1745462530
transform 1 0 1764 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_747
timestamp 1745462530
transform 1 0 1628 0 1 2835
box -2 -2 2 2
use M2_M1  M2_M1_748
timestamp 1745462530
transform 1 0 1612 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_749
timestamp 1745462530
transform 1 0 1316 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_750
timestamp 1745462530
transform 1 0 1276 0 1 2825
box -2 -2 2 2
use M2_M1  M2_M1_751
timestamp 1745462530
transform 1 0 1996 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_752
timestamp 1745462530
transform 1 0 1916 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_753
timestamp 1745462530
transform 1 0 1716 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_754
timestamp 1745462530
transform 1 0 1652 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_755
timestamp 1745462530
transform 1 0 1572 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_756
timestamp 1745462530
transform 1 0 1308 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_757
timestamp 1745462530
transform 1 0 1244 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_758
timestamp 1745462530
transform 1 0 1916 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_759
timestamp 1745462530
transform 1 0 1844 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_760
timestamp 1745462530
transform 1 0 1700 0 1 2722
box -2 -2 2 2
use M2_M1  M2_M1_761
timestamp 1745462530
transform 1 0 1692 0 1 2635
box -2 -2 2 2
use M2_M1  M2_M1_762
timestamp 1745462530
transform 1 0 1564 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_763
timestamp 1745462530
transform 1 0 1292 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_764
timestamp 1745462530
transform 1 0 1244 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_765
timestamp 1745462530
transform 1 0 484 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_766
timestamp 1745462530
transform 1 0 436 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_767
timestamp 1745462530
transform 1 0 372 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_768
timestamp 1745462530
transform 1 0 300 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_769
timestamp 1745462530
transform 1 0 244 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_770
timestamp 1745462530
transform 1 0 228 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_771
timestamp 1745462530
transform 1 0 220 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_772
timestamp 1745462530
transform 1 0 444 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_773
timestamp 1745462530
transform 1 0 436 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_774
timestamp 1745462530
transform 1 0 356 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_775
timestamp 1745462530
transform 1 0 292 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_776
timestamp 1745462530
transform 1 0 228 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_777
timestamp 1745462530
transform 1 0 212 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_778
timestamp 1745462530
transform 1 0 196 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_779
timestamp 1745462530
transform 1 0 732 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_780
timestamp 1745462530
transform 1 0 700 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_781
timestamp 1745462530
transform 1 0 676 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_782
timestamp 1745462530
transform 1 0 628 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_783
timestamp 1745462530
transform 1 0 628 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_784
timestamp 1745462530
transform 1 0 588 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_785
timestamp 1745462530
transform 1 0 532 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_786
timestamp 1745462530
transform 1 0 500 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_787
timestamp 1745462530
transform 1 0 436 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_788
timestamp 1745462530
transform 1 0 380 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_789
timestamp 1745462530
transform 1 0 372 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_790
timestamp 1745462530
transform 1 0 364 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_791
timestamp 1745462530
transform 1 0 308 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_792
timestamp 1745462530
transform 1 0 236 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_793
timestamp 1745462530
transform 1 0 932 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_794
timestamp 1745462530
transform 1 0 916 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_795
timestamp 1745462530
transform 1 0 916 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_796
timestamp 1745462530
transform 1 0 892 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_797
timestamp 1745462530
transform 1 0 860 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_798
timestamp 1745462530
transform 1 0 852 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_799
timestamp 1745462530
transform 1 0 852 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_800
timestamp 1745462530
transform 1 0 836 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_801
timestamp 1745462530
transform 1 0 500 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_802
timestamp 1745462530
transform 1 0 428 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_803
timestamp 1745462530
transform 1 0 396 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_804
timestamp 1745462530
transform 1 0 332 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_805
timestamp 1745462530
transform 1 0 228 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_806
timestamp 1745462530
transform 1 0 212 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_807
timestamp 1745462530
transform 1 0 212 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_808
timestamp 1745462530
transform 1 0 964 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_809
timestamp 1745462530
transform 1 0 876 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_810
timestamp 1745462530
transform 1 0 860 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_811
timestamp 1745462530
transform 1 0 812 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_812
timestamp 1745462530
transform 1 0 780 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_813
timestamp 1745462530
transform 1 0 716 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_814
timestamp 1745462530
transform 1 0 700 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_815
timestamp 1745462530
transform 1 0 1708 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_816
timestamp 1745462530
transform 1 0 1644 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_817
timestamp 1745462530
transform 1 0 1508 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_818
timestamp 1745462530
transform 1 0 1508 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_819
timestamp 1745462530
transform 1 0 1484 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_820
timestamp 1745462530
transform 1 0 1180 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_821
timestamp 1745462530
transform 1 0 1140 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_822
timestamp 1745462530
transform 1 0 1124 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_823
timestamp 1745462530
transform 1 0 2044 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_824
timestamp 1745462530
transform 1 0 2020 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_825
timestamp 1745462530
transform 1 0 1964 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_826
timestamp 1745462530
transform 1 0 1804 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_827
timestamp 1745462530
transform 1 0 1612 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_828
timestamp 1745462530
transform 1 0 1436 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_829
timestamp 1745462530
transform 1 0 1436 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_830
timestamp 1745462530
transform 1 0 2020 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_831
timestamp 1745462530
transform 1 0 2012 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_832
timestamp 1745462530
transform 1 0 1852 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_833
timestamp 1745462530
transform 1 0 1636 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_834
timestamp 1745462530
transform 1 0 1604 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_835
timestamp 1745462530
transform 1 0 1484 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_836
timestamp 1745462530
transform 1 0 1428 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_837
timestamp 1745462530
transform 1 0 2044 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_838
timestamp 1745462530
transform 1 0 2012 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_839
timestamp 1745462530
transform 1 0 1948 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_840
timestamp 1745462530
transform 1 0 1852 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_841
timestamp 1745462530
transform 1 0 1676 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_842
timestamp 1745462530
transform 1 0 1612 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_843
timestamp 1745462530
transform 1 0 1540 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_844
timestamp 1745462530
transform 1 0 2916 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_845
timestamp 1745462530
transform 1 0 2860 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_846
timestamp 1745462530
transform 1 0 2756 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_847
timestamp 1745462530
transform 1 0 2548 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_848
timestamp 1745462530
transform 1 0 2380 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_849
timestamp 1745462530
transform 1 0 2316 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_850
timestamp 1745462530
transform 1 0 2252 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_851
timestamp 1745462530
transform 1 0 2924 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_852
timestamp 1745462530
transform 1 0 2916 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_853
timestamp 1745462530
transform 1 0 2748 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_854
timestamp 1745462530
transform 1 0 2740 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_855
timestamp 1745462530
transform 1 0 2572 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_856
timestamp 1745462530
transform 1 0 2364 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_857
timestamp 1745462530
transform 1 0 2300 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_858
timestamp 1745462530
transform 1 0 2868 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_859
timestamp 1745462530
transform 1 0 2852 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_860
timestamp 1745462530
transform 1 0 2692 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_861
timestamp 1745462530
transform 1 0 2636 0 1 1115
box -2 -2 2 2
use M2_M1  M2_M1_862
timestamp 1745462530
transform 1 0 2620 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_863
timestamp 1745462530
transform 1 0 2380 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_864
timestamp 1745462530
transform 1 0 2316 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_865
timestamp 1745462530
transform 1 0 2860 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_866
timestamp 1745462530
transform 1 0 2820 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_867
timestamp 1745462530
transform 1 0 2692 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_868
timestamp 1745462530
transform 1 0 2652 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_869
timestamp 1745462530
transform 1 0 2620 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_870
timestamp 1745462530
transform 1 0 2412 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_871
timestamp 1745462530
transform 1 0 2388 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_872
timestamp 1745462530
transform 1 0 3452 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_873
timestamp 1745462530
transform 1 0 3396 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_874
timestamp 1745462530
transform 1 0 3340 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_875
timestamp 1745462530
transform 1 0 3340 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_876
timestamp 1745462530
transform 1 0 3324 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_877
timestamp 1745462530
transform 1 0 3284 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_878
timestamp 1745462530
transform 1 0 3228 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_879
timestamp 1745462530
transform 1 0 4324 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_880
timestamp 1745462530
transform 1 0 4260 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_881
timestamp 1745462530
transform 1 0 4244 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_882
timestamp 1745462530
transform 1 0 4204 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_883
timestamp 1745462530
transform 1 0 4164 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_884
timestamp 1745462530
transform 1 0 4076 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_885
timestamp 1745462530
transform 1 0 3972 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_886
timestamp 1745462530
transform 1 0 4236 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_887
timestamp 1745462530
transform 1 0 4172 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_888
timestamp 1745462530
transform 1 0 4148 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_889
timestamp 1745462530
transform 1 0 4084 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_890
timestamp 1745462530
transform 1 0 3820 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_891
timestamp 1745462530
transform 1 0 3468 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_892
timestamp 1745462530
transform 1 0 3404 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_893
timestamp 1745462530
transform 1 0 3940 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_894
timestamp 1745462530
transform 1 0 3892 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_895
timestamp 1745462530
transform 1 0 3812 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_896
timestamp 1745462530
transform 1 0 3796 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_897
timestamp 1745462530
transform 1 0 3628 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_898
timestamp 1745462530
transform 1 0 3476 0 1 1216
box -2 -2 2 2
use M2_M1  M2_M1_899
timestamp 1745462530
transform 1 0 3388 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_900
timestamp 1745462530
transform 1 0 4236 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_901
timestamp 1745462530
transform 1 0 4228 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_902
timestamp 1745462530
transform 1 0 4164 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_903
timestamp 1745462530
transform 1 0 4140 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_904
timestamp 1745462530
transform 1 0 4124 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_905
timestamp 1745462530
transform 1 0 4108 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_906
timestamp 1745462530
transform 1 0 4100 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_907
timestamp 1745462530
transform 1 0 3892 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_908
timestamp 1745462530
transform 1 0 3868 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_909
timestamp 1745462530
transform 1 0 3732 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_910
timestamp 1745462530
transform 1 0 3596 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_911
timestamp 1745462530
transform 1 0 3396 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_912
timestamp 1745462530
transform 1 0 3300 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_913
timestamp 1745462530
transform 1 0 3292 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_914
timestamp 1745462530
transform 1 0 3132 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_915
timestamp 1745462530
transform 1 0 2988 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_916
timestamp 1745462530
transform 1 0 2988 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_917
timestamp 1745462530
transform 1 0 2884 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_918
timestamp 1745462530
transform 1 0 2852 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_919
timestamp 1745462530
transform 1 0 2804 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_920
timestamp 1745462530
transform 1 0 2788 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_921
timestamp 1745462530
transform 1 0 2948 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_922
timestamp 1745462530
transform 1 0 2788 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_923
timestamp 1745462530
transform 1 0 2716 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_924
timestamp 1745462530
transform 1 0 2700 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_925
timestamp 1745462530
transform 1 0 2684 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_926
timestamp 1745462530
transform 1 0 2652 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_927
timestamp 1745462530
transform 1 0 2644 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_928
timestamp 1745462530
transform 1 0 4212 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_929
timestamp 1745462530
transform 1 0 4204 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_930
timestamp 1745462530
transform 1 0 3884 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_931
timestamp 1745462530
transform 1 0 3708 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_932
timestamp 1745462530
transform 1 0 3692 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_933
timestamp 1745462530
transform 1 0 3460 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_934
timestamp 1745462530
transform 1 0 3292 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_935
timestamp 1745462530
transform 1 0 3932 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_936
timestamp 1745462530
transform 1 0 3916 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_937
timestamp 1745462530
transform 1 0 3900 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_938
timestamp 1745462530
transform 1 0 3780 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_939
timestamp 1745462530
transform 1 0 3716 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_940
timestamp 1745462530
transform 1 0 3244 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_941
timestamp 1745462530
transform 1 0 3020 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_942
timestamp 1745462530
transform 1 0 4164 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_943
timestamp 1745462530
transform 1 0 4100 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_944
timestamp 1745462530
transform 1 0 3996 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_945
timestamp 1745462530
transform 1 0 3876 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_946
timestamp 1745462530
transform 1 0 3644 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_947
timestamp 1745462530
transform 1 0 3412 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_948
timestamp 1745462530
transform 1 0 3268 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_949
timestamp 1745462530
transform 1 0 4244 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_950
timestamp 1745462530
transform 1 0 4212 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_951
timestamp 1745462530
transform 1 0 4188 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_952
timestamp 1745462530
transform 1 0 3748 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_953
timestamp 1745462530
transform 1 0 3548 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_954
timestamp 1745462530
transform 1 0 3308 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_955
timestamp 1745462530
transform 1 0 3220 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_956
timestamp 1745462530
transform 1 0 4236 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_957
timestamp 1745462530
transform 1 0 4228 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_958
timestamp 1745462530
transform 1 0 3948 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_959
timestamp 1745462530
transform 1 0 3852 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_960
timestamp 1745462530
transform 1 0 3676 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_961
timestamp 1745462530
transform 1 0 3476 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_962
timestamp 1745462530
transform 1 0 3300 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_963
timestamp 1745462530
transform 1 0 3012 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_964
timestamp 1745462530
transform 1 0 2900 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_965
timestamp 1745462530
transform 1 0 2892 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_966
timestamp 1745462530
transform 1 0 2884 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_967
timestamp 1745462530
transform 1 0 2828 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_968
timestamp 1745462530
transform 1 0 2812 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_969
timestamp 1745462530
transform 1 0 2812 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_970
timestamp 1745462530
transform 1 0 2828 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_971
timestamp 1745462530
transform 1 0 2812 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_972
timestamp 1745462530
transform 1 0 2788 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_973
timestamp 1745462530
transform 1 0 2708 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_974
timestamp 1745462530
transform 1 0 2644 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_975
timestamp 1745462530
transform 1 0 2628 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_976
timestamp 1745462530
transform 1 0 2516 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_977
timestamp 1745462530
transform 1 0 1052 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_978
timestamp 1745462530
transform 1 0 1036 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_979
timestamp 1745462530
transform 1 0 1308 0 1 3025
box -2 -2 2 2
use M2_M1  M2_M1_980
timestamp 1745462530
transform 1 0 1124 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_981
timestamp 1745462530
transform 1 0 1068 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_982
timestamp 1745462530
transform 1 0 1060 0 1 3225
box -2 -2 2 2
use M2_M1  M2_M1_983
timestamp 1745462530
transform 1 0 996 0 1 3715
box -2 -2 2 2
use M2_M1  M2_M1_984
timestamp 1745462530
transform 1 0 972 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_985
timestamp 1745462530
transform 1 0 1348 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_986
timestamp 1745462530
transform 1 0 1300 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_987
timestamp 1745462530
transform 1 0 1268 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_988
timestamp 1745462530
transform 1 0 1100 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_989
timestamp 1745462530
transform 1 0 844 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_990
timestamp 1745462530
transform 1 0 1108 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_991
timestamp 1745462530
transform 1 0 1084 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_992
timestamp 1745462530
transform 1 0 1036 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_993
timestamp 1745462530
transform 1 0 1004 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_994
timestamp 1745462530
transform 1 0 956 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_995
timestamp 1745462530
transform 1 0 868 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_996
timestamp 1745462530
transform 1 0 860 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_997
timestamp 1745462530
transform 1 0 988 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_998
timestamp 1745462530
transform 1 0 820 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_999
timestamp 1745462530
transform 1 0 940 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_1000
timestamp 1745462530
transform 1 0 900 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_1001
timestamp 1745462530
transform 1 0 1692 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_1002
timestamp 1745462530
transform 1 0 1676 0 1 3115
box -2 -2 2 2
use M2_M1  M2_M1_1003
timestamp 1745462530
transform 1 0 1524 0 1 3225
box -2 -2 2 2
use M2_M1  M2_M1_1004
timestamp 1745462530
transform 1 0 1516 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_1005
timestamp 1745462530
transform 1 0 1396 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_1006
timestamp 1745462530
transform 1 0 1372 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_1007
timestamp 1745462530
transform 1 0 1356 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_1008
timestamp 1745462530
transform 1 0 1188 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_1009
timestamp 1745462530
transform 1 0 1588 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_1010
timestamp 1745462530
transform 1 0 1540 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_1011
timestamp 1745462530
transform 1 0 1740 0 1 3225
box -2 -2 2 2
use M2_M1  M2_M1_1012
timestamp 1745462530
transform 1 0 1700 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_1013
timestamp 1745462530
transform 1 0 1660 0 1 3315
box -2 -2 2 2
use M2_M1  M2_M1_1014
timestamp 1745462530
transform 1 0 1636 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_1015
timestamp 1745462530
transform 1 0 1292 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_1016
timestamp 1745462530
transform 1 0 1276 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_1017
timestamp 1745462530
transform 1 0 1100 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_1018
timestamp 1745462530
transform 1 0 1084 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_1019
timestamp 1745462530
transform 1 0 1780 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_1020
timestamp 1745462530
transform 1 0 1740 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_1021
timestamp 1745462530
transform 1 0 1732 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_1022
timestamp 1745462530
transform 1 0 1716 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_1023
timestamp 1745462530
transform 1 0 1668 0 1 3305
box -2 -2 2 2
use M2_M1  M2_M1_1024
timestamp 1745462530
transform 1 0 1620 0 1 3315
box -2 -2 2 2
use M2_M1  M2_M1_1025
timestamp 1745462530
transform 1 0 1604 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_1026
timestamp 1745462530
transform 1 0 2620 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_1027
timestamp 1745462530
transform 1 0 2588 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_1028
timestamp 1745462530
transform 1 0 2572 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_1029
timestamp 1745462530
transform 1 0 2556 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_1030
timestamp 1745462530
transform 1 0 2532 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_1031
timestamp 1745462530
transform 1 0 2468 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_1032
timestamp 1745462530
transform 1 0 2460 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_1033
timestamp 1745462530
transform 1 0 2420 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_1034
timestamp 1745462530
transform 1 0 2156 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_1035
timestamp 1745462530
transform 1 0 2124 0 1 3825
box -2 -2 2 2
use M2_M1  M2_M1_1036
timestamp 1745462530
transform 1 0 3524 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_1037
timestamp 1745462530
transform 1 0 3500 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_1038
timestamp 1745462530
transform 1 0 3460 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_1039
timestamp 1745462530
transform 1 0 3452 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_1040
timestamp 1745462530
transform 1 0 3420 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_1041
timestamp 1745462530
transform 1 0 3380 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_1042
timestamp 1745462530
transform 1 0 3316 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_1043
timestamp 1745462530
transform 1 0 3308 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_1044
timestamp 1745462530
transform 1 0 3252 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_1045
timestamp 1745462530
transform 1 0 3140 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_1046
timestamp 1745462530
transform 1 0 1972 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_1047
timestamp 1745462530
transform 1 0 1908 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_1048
timestamp 1745462530
transform 1 0 1828 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_1049
timestamp 1745462530
transform 1 0 1724 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_1050
timestamp 1745462530
transform 1 0 1556 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_1051
timestamp 1745462530
transform 1 0 1548 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_1052
timestamp 1745462530
transform 1 0 1540 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_1053
timestamp 1745462530
transform 1 0 1532 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_1054
timestamp 1745462530
transform 1 0 3580 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_1055
timestamp 1745462530
transform 1 0 3580 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_1056
timestamp 1745462530
transform 1 0 3564 0 1 3705
box -2 -2 2 2
use M2_M1  M2_M1_1057
timestamp 1745462530
transform 1 0 3524 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_1058
timestamp 1745462530
transform 1 0 3500 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_1059
timestamp 1745462530
transform 1 0 3404 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_1060
timestamp 1745462530
transform 1 0 3364 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_1061
timestamp 1745462530
transform 1 0 3276 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_1062
timestamp 1745462530
transform 1 0 3228 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_1063
timestamp 1745462530
transform 1 0 1644 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_1064
timestamp 1745462530
transform 1 0 2908 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_1065
timestamp 1745462530
transform 1 0 2900 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_1066
timestamp 1745462530
transform 1 0 2812 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_1067
timestamp 1745462530
transform 1 0 2796 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_1068
timestamp 1745462530
transform 1 0 2788 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_1069
timestamp 1745462530
transform 1 0 2780 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_1070
timestamp 1745462530
transform 1 0 2772 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_1071
timestamp 1745462530
transform 1 0 2764 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_1072
timestamp 1745462530
transform 1 0 2748 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_1073
timestamp 1745462530
transform 1 0 2748 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_1074
timestamp 1745462530
transform 1 0 2732 0 1 3555
box -2 -2 2 2
use M2_M1  M2_M1_1075
timestamp 1745462530
transform 1 0 2700 0 1 3825
box -2 -2 2 2
use M2_M1  M2_M1_1076
timestamp 1745462530
transform 1 0 1588 0 1 3515
box -2 -2 2 2
use M2_M1  M2_M1_1077
timestamp 1745462530
transform 1 0 1564 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_1078
timestamp 1745462530
transform 1 0 1668 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_1079
timestamp 1745462530
transform 1 0 1660 0 1 3715
box -2 -2 2 2
use M2_M1  M2_M1_1080
timestamp 1745462530
transform 1 0 1644 0 1 3625
box -2 -2 2 2
use M2_M1  M2_M1_1081
timestamp 1745462530
transform 1 0 1604 0 1 3635
box -2 -2 2 2
use M2_M1  M2_M1_1082
timestamp 1745462530
transform 1 0 1580 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_1083
timestamp 1745462530
transform 1 0 1548 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_1084
timestamp 1745462530
transform 1 0 1452 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_1085
timestamp 1745462530
transform 1 0 1420 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_1086
timestamp 1745462530
transform 1 0 1420 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_1087
timestamp 1745462530
transform 1 0 1812 0 1 3625
box -2 -2 2 2
use M2_M1  M2_M1_1088
timestamp 1745462530
transform 1 0 1804 0 1 3545
box -2 -2 2 2
use M2_M1  M2_M1_1089
timestamp 1745462530
transform 1 0 1804 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_1090
timestamp 1745462530
transform 1 0 1780 0 1 3515
box -2 -2 2 2
use M2_M1  M2_M1_1091
timestamp 1745462530
transform 1 0 1780 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_1092
timestamp 1745462530
transform 1 0 1836 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_1093
timestamp 1745462530
transform 1 0 1788 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_1094
timestamp 1745462530
transform 1 0 1676 0 1 3625
box -2 -2 2 2
use M2_M1  M2_M1_1095
timestamp 1745462530
transform 1 0 1660 0 1 3705
box -2 -2 2 2
use M2_M1  M2_M1_1096
timestamp 1745462530
transform 1 0 1588 0 1 3625
box -2 -2 2 2
use M2_M1  M2_M1_1097
timestamp 1745462530
transform 1 0 1428 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_1098
timestamp 1745462530
transform 1 0 1348 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_1099
timestamp 1745462530
transform 1 0 1284 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_1100
timestamp 1745462530
transform 1 0 1252 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_1101
timestamp 1745462530
transform 1 0 1252 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_1102
timestamp 1745462530
transform 1 0 1308 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_1103
timestamp 1745462530
transform 1 0 1308 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_1104
timestamp 1745462530
transform 1 0 628 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_1105
timestamp 1745462530
transform 1 0 572 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_1106
timestamp 1745462530
transform 1 0 468 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_1107
timestamp 1745462530
transform 1 0 372 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_1108
timestamp 1745462530
transform 1 0 260 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_1109
timestamp 1745462530
transform 1 0 260 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_1110
timestamp 1745462530
transform 1 0 188 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_1111
timestamp 1745462530
transform 1 0 140 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_1112
timestamp 1745462530
transform 1 0 188 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_1113
timestamp 1745462530
transform 1 0 148 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_1114
timestamp 1745462530
transform 1 0 308 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_1115
timestamp 1745462530
transform 1 0 308 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_1116
timestamp 1745462530
transform 1 0 412 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_1117
timestamp 1745462530
transform 1 0 412 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_1118
timestamp 1745462530
transform 1 0 636 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_1119
timestamp 1745462530
transform 1 0 620 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_1120
timestamp 1745462530
transform 1 0 828 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_1121
timestamp 1745462530
transform 1 0 820 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_1122
timestamp 1745462530
transform 1 0 796 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_1123
timestamp 1745462530
transform 1 0 1852 0 1 3515
box -2 -2 2 2
use M2_M1  M2_M1_1124
timestamp 1745462530
transform 1 0 1844 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_1125
timestamp 1745462530
transform 1 0 1780 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_1126
timestamp 1745462530
transform 1 0 1708 0 1 3515
box -2 -2 2 2
use M2_M1  M2_M1_1127
timestamp 1745462530
transform 1 0 1692 0 1 3395
box -2 -2 2 2
use M2_M1  M2_M1_1128
timestamp 1745462530
transform 1 0 1636 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_1129
timestamp 1745462530
transform 1 0 1628 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_1130
timestamp 1745462530
transform 1 0 1028 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_1131
timestamp 1745462530
transform 1 0 988 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_1132
timestamp 1745462530
transform 1 0 884 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_1133
timestamp 1745462530
transform 1 0 1268 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_1134
timestamp 1745462530
transform 1 0 1204 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_1135
timestamp 1745462530
transform 1 0 1164 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_1136
timestamp 1745462530
transform 1 0 1260 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_1137
timestamp 1745462530
transform 1 0 1220 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1138
timestamp 1745462530
transform 1 0 1268 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_1139
timestamp 1745462530
transform 1 0 1260 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_1140
timestamp 1745462530
transform 1 0 1220 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_1141
timestamp 1745462530
transform 1 0 1244 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_1142
timestamp 1745462530
transform 1 0 1228 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_1143
timestamp 1745462530
transform 1 0 1140 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1144
timestamp 1745462530
transform 1 0 1212 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_1145
timestamp 1745462530
transform 1 0 1164 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_1146
timestamp 1745462530
transform 1 0 1148 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_1147
timestamp 1745462530
transform 1 0 1188 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_1148
timestamp 1745462530
transform 1 0 1148 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_1149
timestamp 1745462530
transform 1 0 1132 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_1150
timestamp 1745462530
transform 1 0 868 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_1151
timestamp 1745462530
transform 1 0 868 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_1152
timestamp 1745462530
transform 1 0 860 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_1153
timestamp 1745462530
transform 1 0 828 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_1154
timestamp 1745462530
transform 1 0 812 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_1155
timestamp 1745462530
transform 1 0 804 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_1156
timestamp 1745462530
transform 1 0 900 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_1157
timestamp 1745462530
transform 1 0 868 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_1158
timestamp 1745462530
transform 1 0 244 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_1159
timestamp 1745462530
transform 1 0 188 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_1160
timestamp 1745462530
transform 1 0 228 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_1161
timestamp 1745462530
transform 1 0 172 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_1162
timestamp 1745462530
transform 1 0 236 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_1163
timestamp 1745462530
transform 1 0 196 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1164
timestamp 1745462530
transform 1 0 588 0 1 955
box -2 -2 2 2
use M2_M1  M2_M1_1165
timestamp 1745462530
transform 1 0 300 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_1166
timestamp 1745462530
transform 1 0 252 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_1167
timestamp 1745462530
transform 1 0 196 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_1168
timestamp 1745462530
transform 1 0 236 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_1169
timestamp 1745462530
transform 1 0 228 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_1170
timestamp 1745462530
transform 1 0 660 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_1171
timestamp 1745462530
transform 1 0 340 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_1172
timestamp 1745462530
transform 1 0 260 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_1173
timestamp 1745462530
transform 1 0 220 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1174
timestamp 1745462530
transform 1 0 308 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_1175
timestamp 1745462530
transform 1 0 236 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_1176
timestamp 1745462530
transform 1 0 748 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_1177
timestamp 1745462530
transform 1 0 708 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_1178
timestamp 1745462530
transform 1 0 236 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_1179
timestamp 1745462530
transform 1 0 204 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_1180
timestamp 1745462530
transform 1 0 1188 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1181
timestamp 1745462530
transform 1 0 1156 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_1182
timestamp 1745462530
transform 1 0 1100 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_1183
timestamp 1745462530
transform 1 0 1100 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_1184
timestamp 1745462530
transform 1 0 1180 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_1185
timestamp 1745462530
transform 1 0 1172 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1186
timestamp 1745462530
transform 1 0 1140 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1187
timestamp 1745462530
transform 1 0 1140 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_1188
timestamp 1745462530
transform 1 0 1348 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_1189
timestamp 1745462530
transform 1 0 1332 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_1190
timestamp 1745462530
transform 1 0 1204 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_1191
timestamp 1745462530
transform 1 0 1140 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_1192
timestamp 1745462530
transform 1 0 1372 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_1193
timestamp 1745462530
transform 1 0 1316 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_1194
timestamp 1745462530
transform 1 0 1316 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_1195
timestamp 1745462530
transform 1 0 1452 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_1196
timestamp 1745462530
transform 1 0 1412 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_1197
timestamp 1745462530
transform 1 0 1444 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_1198
timestamp 1745462530
transform 1 0 1404 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_1199
timestamp 1745462530
transform 1 0 1492 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_1200
timestamp 1745462530
transform 1 0 1420 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_1201
timestamp 1745462530
transform 1 0 1548 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_1202
timestamp 1745462530
transform 1 0 1508 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_1203
timestamp 1745462530
transform 1 0 2356 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_1204
timestamp 1745462530
transform 1 0 2340 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_1205
timestamp 1745462530
transform 1 0 2324 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_1206
timestamp 1745462530
transform 1 0 2228 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_1207
timestamp 1745462530
transform 1 0 2292 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_1208
timestamp 1745462530
transform 1 0 2276 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_1209
timestamp 1745462530
transform 1 0 2476 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1210
timestamp 1745462530
transform 1 0 2396 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_1211
timestamp 1745462530
transform 1 0 2324 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_1212
timestamp 1745462530
transform 1 0 2204 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_1213
timestamp 1745462530
transform 1 0 2428 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1214
timestamp 1745462530
transform 1 0 2348 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1215
timestamp 1745462530
transform 1 0 2628 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_1216
timestamp 1745462530
transform 1 0 2596 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_1217
timestamp 1745462530
transform 1 0 2580 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_1218
timestamp 1745462530
transform 1 0 2548 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_1219
timestamp 1745462530
transform 1 0 3468 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1220
timestamp 1745462530
transform 1 0 3428 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_1221
timestamp 1745462530
transform 1 0 3348 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_1222
timestamp 1745462530
transform 1 0 3340 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_1223
timestamp 1745462530
transform 1 0 3548 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_1224
timestamp 1745462530
transform 1 0 3452 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1225
timestamp 1745462530
transform 1 0 4036 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_1226
timestamp 1745462530
transform 1 0 3980 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1227
timestamp 1745462530
transform 1 0 3588 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_1228
timestamp 1745462530
transform 1 0 3444 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_1229
timestamp 1745462530
transform 1 0 3572 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_1230
timestamp 1745462530
transform 1 0 3572 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_1231
timestamp 1745462530
transform 1 0 4116 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_1232
timestamp 1745462530
transform 1 0 4084 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_1233
timestamp 1745462530
transform 1 0 3980 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_1234
timestamp 1745462530
transform 1 0 3940 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_1235
timestamp 1745462530
transform 1 0 3476 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_1236
timestamp 1745462530
transform 1 0 3428 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_1237
timestamp 1745462530
transform 1 0 4116 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_1238
timestamp 1745462530
transform 1 0 3948 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_1239
timestamp 1745462530
transform 1 0 3540 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_1240
timestamp 1745462530
transform 1 0 3540 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_1241
timestamp 1745462530
transform 1 0 3500 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_1242
timestamp 1745462530
transform 1 0 3492 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_1243
timestamp 1745462530
transform 1 0 3468 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_1244
timestamp 1745462530
transform 1 0 4140 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_1245
timestamp 1745462530
transform 1 0 4100 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_1246
timestamp 1745462530
transform 1 0 3668 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_1247
timestamp 1745462530
transform 1 0 3596 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_1248
timestamp 1745462530
transform 1 0 3708 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_1249
timestamp 1745462530
transform 1 0 3620 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_1250
timestamp 1745462530
transform 1 0 3620 0 1 1945
box -2 -2 2 2
use M2_M1  M2_M1_1251
timestamp 1745462530
transform 1 0 4164 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_1252
timestamp 1745462530
transform 1 0 4132 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_1253
timestamp 1745462530
transform 1 0 3404 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_1254
timestamp 1745462530
transform 1 0 3356 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1255
timestamp 1745462530
transform 1 0 2820 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_1256
timestamp 1745462530
transform 1 0 2820 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_1257
timestamp 1745462530
transform 1 0 2652 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_1258
timestamp 1745462530
transform 1 0 2612 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1259
timestamp 1745462530
transform 1 0 3260 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_1260
timestamp 1745462530
transform 1 0 3252 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_1261
timestamp 1745462530
transform 1 0 3540 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_1262
timestamp 1745462530
transform 1 0 3420 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_1263
timestamp 1745462530
transform 1 0 3380 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_1264
timestamp 1745462530
transform 1 0 3324 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_1265
timestamp 1745462530
transform 1 0 3316 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_1266
timestamp 1745462530
transform 1 0 3484 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_1267
timestamp 1745462530
transform 1 0 3452 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_1268
timestamp 1745462530
transform 1 0 3412 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_1269
timestamp 1745462530
transform 1 0 3396 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_1270
timestamp 1745462530
transform 1 0 3396 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_1271
timestamp 1745462530
transform 1 0 3380 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_1272
timestamp 1745462530
transform 1 0 3284 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_1273
timestamp 1745462530
transform 1 0 3236 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_1274
timestamp 1745462530
transform 1 0 2804 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_1275
timestamp 1745462530
transform 1 0 2788 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_1276
timestamp 1745462530
transform 1 0 3060 0 1 3105
box -2 -2 2 2
use M2_M1  M2_M1_1277
timestamp 1745462530
transform 1 0 3044 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_1278
timestamp 1745462530
transform 1 0 2964 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_1279
timestamp 1745462530
transform 1 0 2884 0 1 3115
box -2 -2 2 2
use M2_M1  M2_M1_1280
timestamp 1745462530
transform 1 0 2844 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_1281
timestamp 1745462530
transform 1 0 2716 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_1282
timestamp 1745462530
transform 1 0 2684 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_1283
timestamp 1745462530
transform 1 0 932 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_1284
timestamp 1745462530
transform 1 0 924 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_1285
timestamp 1745462530
transform 1 0 900 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_1286
timestamp 1745462530
transform 1 0 868 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_1287
timestamp 1745462530
transform 1 0 1844 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_1288
timestamp 1745462530
transform 1 0 1844 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_1289
timestamp 1745462530
transform 1 0 1836 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_1290
timestamp 1745462530
transform 1 0 1932 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1291
timestamp 1745462530
transform 1 0 1924 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_1292
timestamp 1745462530
transform 1 0 1884 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_1293
timestamp 1745462530
transform 1 0 1876 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_1294
timestamp 1745462530
transform 1 0 1900 0 1 2145
box -2 -2 2 2
use M2_M1  M2_M1_1295
timestamp 1745462530
transform 1 0 1892 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_1296
timestamp 1745462530
transform 1 0 1884 0 1 2145
box -2 -2 2 2
use M2_M1  M2_M1_1297
timestamp 1745462530
transform 1 0 1868 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_1298
timestamp 1745462530
transform 1 0 1812 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_1299
timestamp 1745462530
transform 1 0 1796 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_1300
timestamp 1745462530
transform 1 0 1764 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_1301
timestamp 1745462530
transform 1 0 1828 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_1302
timestamp 1745462530
transform 1 0 1748 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_1303
timestamp 1745462530
transform 1 0 804 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_1304
timestamp 1745462530
transform 1 0 804 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_1305
timestamp 1745462530
transform 1 0 780 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_1306
timestamp 1745462530
transform 1 0 780 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_1307
timestamp 1745462530
transform 1 0 772 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_1308
timestamp 1745462530
transform 1 0 748 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_1309
timestamp 1745462530
transform 1 0 716 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_1310
timestamp 1745462530
transform 1 0 708 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_1311
timestamp 1745462530
transform 1 0 884 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_1312
timestamp 1745462530
transform 1 0 820 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_1313
timestamp 1745462530
transform 1 0 500 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_1314
timestamp 1745462530
transform 1 0 468 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_1315
timestamp 1745462530
transform 1 0 388 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_1316
timestamp 1745462530
transform 1 0 380 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_1317
timestamp 1745462530
transform 1 0 756 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_1318
timestamp 1745462530
transform 1 0 380 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_1319
timestamp 1745462530
transform 1 0 324 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_1320
timestamp 1745462530
transform 1 0 316 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_1321
timestamp 1745462530
transform 1 0 284 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_1322
timestamp 1745462530
transform 1 0 252 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_1323
timestamp 1745462530
transform 1 0 228 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_1324
timestamp 1745462530
transform 1 0 804 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_1325
timestamp 1745462530
transform 1 0 324 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1326
timestamp 1745462530
transform 1 0 228 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_1327
timestamp 1745462530
transform 1 0 188 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_1328
timestamp 1745462530
transform 1 0 284 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_1329
timestamp 1745462530
transform 1 0 284 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_1330
timestamp 1745462530
transform 1 0 252 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_1331
timestamp 1745462530
transform 1 0 220 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_1332
timestamp 1745462530
transform 1 0 180 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_1333
timestamp 1745462530
transform 1 0 1988 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_1334
timestamp 1745462530
transform 1 0 1948 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1335
timestamp 1745462530
transform 1 0 1652 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_1336
timestamp 1745462530
transform 1 0 1612 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_1337
timestamp 1745462530
transform 1 0 2076 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1338
timestamp 1745462530
transform 1 0 1948 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_1339
timestamp 1745462530
transform 1 0 1932 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1340
timestamp 1745462530
transform 1 0 2036 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_1341
timestamp 1745462530
transform 1 0 1964 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_1342
timestamp 1745462530
transform 1 0 1964 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_1343
timestamp 1745462530
transform 1 0 1948 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_1344
timestamp 1745462530
transform 1 0 1948 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_1345
timestamp 1745462530
transform 1 0 2028 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_1346
timestamp 1745462530
transform 1 0 1972 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_1347
timestamp 1745462530
transform 1 0 2108 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_1348
timestamp 1745462530
transform 1 0 2052 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_1349
timestamp 1745462530
transform 1 0 2500 0 1 595
box -2 -2 2 2
use M2_M1  M2_M1_1350
timestamp 1745462530
transform 1 0 2484 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_1351
timestamp 1745462530
transform 1 0 2404 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_1352
timestamp 1745462530
transform 1 0 2452 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_1353
timestamp 1745462530
transform 1 0 2316 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_1354
timestamp 1745462530
transform 1 0 2572 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_1355
timestamp 1745462530
transform 1 0 2556 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_1356
timestamp 1745462530
transform 1 0 2548 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_1357
timestamp 1745462530
transform 1 0 2532 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1358
timestamp 1745462530
transform 1 0 2492 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1359
timestamp 1745462530
transform 1 0 2356 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1360
timestamp 1745462530
transform 1 0 2340 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_1361
timestamp 1745462530
transform 1 0 2548 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_1362
timestamp 1745462530
transform 1 0 2500 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_1363
timestamp 1745462530
transform 1 0 2308 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_1364
timestamp 1745462530
transform 1 0 2308 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_1365
timestamp 1745462530
transform 1 0 2628 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_1366
timestamp 1745462530
transform 1 0 2588 0 1 1115
box -2 -2 2 2
use M2_M1  M2_M1_1367
timestamp 1745462530
transform 1 0 2628 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_1368
timestamp 1745462530
transform 1 0 2588 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_1369
timestamp 1745462530
transform 1 0 3684 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_1370
timestamp 1745462530
transform 1 0 3628 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1371
timestamp 1745462530
transform 1 0 3532 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_1372
timestamp 1745462530
transform 1 0 3420 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_1373
timestamp 1745462530
transform 1 0 3764 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_1374
timestamp 1745462530
transform 1 0 3644 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1375
timestamp 1745462530
transform 1 0 3612 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1376
timestamp 1745462530
transform 1 0 4244 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_1377
timestamp 1745462530
transform 1 0 3732 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_1378
timestamp 1745462530
transform 1 0 3732 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_1379
timestamp 1745462530
transform 1 0 3804 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_1380
timestamp 1745462530
transform 1 0 3804 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_1381
timestamp 1745462530
transform 1 0 3700 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_1382
timestamp 1745462530
transform 1 0 4180 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_1383
timestamp 1745462530
transform 1 0 4132 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_1384
timestamp 1745462530
transform 1 0 3828 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_1385
timestamp 1745462530
transform 1 0 3788 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_1386
timestamp 1745462530
transform 1 0 3804 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_1387
timestamp 1745462530
transform 1 0 3764 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_1388
timestamp 1745462530
transform 1 0 4196 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_1389
timestamp 1745462530
transform 1 0 4180 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_1390
timestamp 1745462530
transform 1 0 3900 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_1391
timestamp 1745462530
transform 1 0 3748 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_1392
timestamp 1745462530
transform 1 0 4244 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_1393
timestamp 1745462530
transform 1 0 3892 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_1394
timestamp 1745462530
transform 1 0 3788 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_1395
timestamp 1745462530
transform 1 0 3876 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_1396
timestamp 1745462530
transform 1 0 3852 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_1397
timestamp 1745462530
transform 1 0 3836 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_1398
timestamp 1745462530
transform 1 0 4012 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_1399
timestamp 1745462530
transform 1 0 3940 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_1400
timestamp 1745462530
transform 1 0 2724 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_1401
timestamp 1745462530
transform 1 0 2692 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_1402
timestamp 1745462530
transform 1 0 3892 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_1403
timestamp 1745462530
transform 1 0 3804 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_1404
timestamp 1745462530
transform 1 0 3772 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_1405
timestamp 1745462530
transform 1 0 3788 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_1406
timestamp 1745462530
transform 1 0 3756 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_1407
timestamp 1745462530
transform 1 0 3884 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_1408
timestamp 1745462530
transform 1 0 3844 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_1409
timestamp 1745462530
transform 1 0 3820 0 1 2745
box -2 -2 2 2
use M2_M1  M2_M1_1410
timestamp 1745462530
transform 1 0 3772 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_1411
timestamp 1745462530
transform 1 0 3756 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_1412
timestamp 1745462530
transform 1 0 3908 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_1413
timestamp 1745462530
transform 1 0 3868 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_1414
timestamp 1745462530
transform 1 0 3820 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_1415
timestamp 1745462530
transform 1 0 3956 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_1416
timestamp 1745462530
transform 1 0 3900 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_1417
timestamp 1745462530
transform 1 0 3892 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_1418
timestamp 1745462530
transform 1 0 3868 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_1419
timestamp 1745462530
transform 1 0 3836 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_1420
timestamp 1745462530
transform 1 0 3004 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_1421
timestamp 1745462530
transform 1 0 2988 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_1422
timestamp 1745462530
transform 1 0 3012 0 1 3115
box -2 -2 2 2
use M2_M1  M2_M1_1423
timestamp 1745462530
transform 1 0 3012 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_1424
timestamp 1745462530
transform 1 0 2924 0 1 3105
box -2 -2 2 2
use M2_M1  M2_M1_1425
timestamp 1745462530
transform 1 0 2924 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_1426
timestamp 1745462530
transform 1 0 2884 0 1 3105
box -2 -2 2 2
use M2_M1  M2_M1_1427
timestamp 1745462530
transform 1 0 2844 0 1 3025
box -2 -2 2 2
use M2_M1  M2_M1_1428
timestamp 1745462530
transform 1 0 2524 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_1429
timestamp 1745462530
transform 1 0 2492 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_1430
timestamp 1745462530
transform 1 0 988 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_1431
timestamp 1745462530
transform 1 0 916 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_1432
timestamp 1745462530
transform 1 0 724 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_1433
timestamp 1745462530
transform 1 0 1772 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_1434
timestamp 1745462530
transform 1 0 1700 0 1 2825
box -2 -2 2 2
use M2_M1  M2_M1_1435
timestamp 1745462530
transform 1 0 1732 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_1436
timestamp 1745462530
transform 1 0 1668 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1437
timestamp 1745462530
transform 1 0 1708 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_1438
timestamp 1745462530
transform 1 0 1676 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_1439
timestamp 1745462530
transform 1 0 1668 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_1440
timestamp 1745462530
transform 1 0 1660 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_1441
timestamp 1745462530
transform 1 0 1620 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_1442
timestamp 1745462530
transform 1 0 1580 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_1443
timestamp 1745462530
transform 1 0 1580 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_1444
timestamp 1745462530
transform 1 0 1588 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_1445
timestamp 1745462530
transform 1 0 1564 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_1446
timestamp 1745462530
transform 1 0 1532 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_1447
timestamp 1745462530
transform 1 0 652 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_1448
timestamp 1745462530
transform 1 0 564 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_1449
timestamp 1745462530
transform 1 0 452 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_1450
timestamp 1745462530
transform 1 0 420 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_1451
timestamp 1745462530
transform 1 0 636 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_1452
timestamp 1745462530
transform 1 0 548 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_1453
timestamp 1745462530
transform 1 0 540 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_1454
timestamp 1745462530
transform 1 0 740 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_1455
timestamp 1745462530
transform 1 0 604 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_1456
timestamp 1745462530
transform 1 0 364 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_1457
timestamp 1745462530
transform 1 0 332 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_1458
timestamp 1745462530
transform 1 0 388 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_1459
timestamp 1745462530
transform 1 0 380 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_1460
timestamp 1745462530
transform 1 0 500 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1461
timestamp 1745462530
transform 1 0 492 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_1462
timestamp 1745462530
transform 1 0 460 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_1463
timestamp 1745462530
transform 1 0 452 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_1464
timestamp 1745462530
transform 1 0 476 0 1 745
box -2 -2 2 2
use M2_M1  M2_M1_1465
timestamp 1745462530
transform 1 0 444 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_1466
timestamp 1745462530
transform 1 0 428 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_1467
timestamp 1745462530
transform 1 0 428 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_1468
timestamp 1745462530
transform 1 0 412 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_1469
timestamp 1745462530
transform 1 0 412 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_1470
timestamp 1745462530
transform 1 0 556 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_1471
timestamp 1745462530
transform 1 0 380 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1472
timestamp 1745462530
transform 1 0 276 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_1473
timestamp 1745462530
transform 1 0 276 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_1474
timestamp 1745462530
transform 1 0 364 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1475
timestamp 1745462530
transform 1 0 364 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_1476
timestamp 1745462530
transform 1 0 572 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_1477
timestamp 1745462530
transform 1 0 564 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_1478
timestamp 1745462530
transform 1 0 868 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_1479
timestamp 1745462530
transform 1 0 860 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_1480
timestamp 1745462530
transform 1 0 788 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_1481
timestamp 1745462530
transform 1 0 780 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_1482
timestamp 1745462530
transform 1 0 1876 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1483
timestamp 1745462530
transform 1 0 1772 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_1484
timestamp 1745462530
transform 1 0 1748 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_1485
timestamp 1745462530
transform 1 0 1860 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1486
timestamp 1745462530
transform 1 0 1860 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_1487
timestamp 1745462530
transform 1 0 1836 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_1488
timestamp 1745462530
transform 1 0 1820 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_1489
timestamp 1745462530
transform 1 0 1788 0 1 595
box -2 -2 2 2
use M2_M1  M2_M1_1490
timestamp 1745462530
transform 1 0 1852 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_1491
timestamp 1745462530
transform 1 0 1796 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_1492
timestamp 1745462530
transform 1 0 1796 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_1493
timestamp 1745462530
transform 1 0 2052 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_1494
timestamp 1745462530
transform 1 0 2012 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_1495
timestamp 1745462530
transform 1 0 2020 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_1496
timestamp 1745462530
transform 1 0 1980 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_1497
timestamp 1745462530
transform 1 0 1956 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_1498
timestamp 1745462530
transform 1 0 1916 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_1499
timestamp 1745462530
transform 1 0 2276 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_1500
timestamp 1745462530
transform 1 0 2260 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_1501
timestamp 1745462530
transform 1 0 2212 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_1502
timestamp 1745462530
transform 1 0 2204 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_1503
timestamp 1745462530
transform 1 0 2220 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_1504
timestamp 1745462530
transform 1 0 2180 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_1505
timestamp 1745462530
transform 1 0 2412 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1506
timestamp 1745462530
transform 1 0 2332 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_1507
timestamp 1745462530
transform 1 0 2276 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_1508
timestamp 1745462530
transform 1 0 2276 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_1509
timestamp 1745462530
transform 1 0 2388 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1510
timestamp 1745462530
transform 1 0 2260 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_1511
timestamp 1745462530
transform 1 0 2220 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_1512
timestamp 1745462530
transform 1 0 2524 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_1513
timestamp 1745462530
transform 1 0 2492 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_1514
timestamp 1745462530
transform 1 0 2324 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_1515
timestamp 1745462530
transform 1 0 2284 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_1516
timestamp 1745462530
transform 1 0 2396 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_1517
timestamp 1745462530
transform 1 0 2356 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_1518
timestamp 1745462530
transform 1 0 3828 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_1519
timestamp 1745462530
transform 1 0 3828 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_1520
timestamp 1745462530
transform 1 0 3516 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_1521
timestamp 1745462530
transform 1 0 3836 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_1522
timestamp 1745462530
transform 1 0 3836 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_1523
timestamp 1745462530
transform 1 0 3812 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_1524
timestamp 1745462530
transform 1 0 4252 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_1525
timestamp 1745462530
transform 1 0 4244 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_1526
timestamp 1745462530
transform 1 0 3932 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_1527
timestamp 1745462530
transform 1 0 3908 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_1528
timestamp 1745462530
transform 1 0 4012 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_1529
timestamp 1745462530
transform 1 0 3996 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_1530
timestamp 1745462530
transform 1 0 3948 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_1531
timestamp 1745462530
transform 1 0 3916 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_1532
timestamp 1745462530
transform 1 0 4268 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_1533
timestamp 1745462530
transform 1 0 4196 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_1534
timestamp 1745462530
transform 1 0 4268 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_1535
timestamp 1745462530
transform 1 0 3596 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_1536
timestamp 1745462530
transform 1 0 3356 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_1537
timestamp 1745462530
transform 1 0 3716 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_1538
timestamp 1745462530
transform 1 0 3644 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_1539
timestamp 1745462530
transform 1 0 3572 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_1540
timestamp 1745462530
transform 1 0 4276 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_1541
timestamp 1745462530
transform 1 0 3644 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_1542
timestamp 1745462530
transform 1 0 3412 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_1543
timestamp 1745462530
transform 1 0 3684 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_1544
timestamp 1745462530
transform 1 0 3620 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_1545
timestamp 1745462530
transform 1 0 3620 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_1546
timestamp 1745462530
transform 1 0 4220 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_1547
timestamp 1745462530
transform 1 0 4156 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_1548
timestamp 1745462530
transform 1 0 4116 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_1549
timestamp 1745462530
transform 1 0 3932 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_1550
timestamp 1745462530
transform 1 0 3924 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_1551
timestamp 1745462530
transform 1 0 4172 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_1552
timestamp 1745462530
transform 1 0 4164 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_1553
timestamp 1745462530
transform 1 0 4132 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_1554
timestamp 1745462530
transform 1 0 4260 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_1555
timestamp 1745462530
transform 1 0 4252 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_1556
timestamp 1745462530
transform 1 0 4244 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_1557
timestamp 1745462530
transform 1 0 4212 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_1558
timestamp 1745462530
transform 1 0 4180 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_1559
timestamp 1745462530
transform 1 0 4164 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_1560
timestamp 1745462530
transform 1 0 4204 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_1561
timestamp 1745462530
transform 1 0 4132 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1562
timestamp 1745462530
transform 1 0 4116 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_1563
timestamp 1745462530
transform 1 0 4092 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_1564
timestamp 1745462530
transform 1 0 4084 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_1565
timestamp 1745462530
transform 1 0 2892 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_1566
timestamp 1745462530
transform 1 0 2844 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_1567
timestamp 1745462530
transform 1 0 2708 0 1 3035
box -2 -2 2 2
use M2_M1  M2_M1_1568
timestamp 1745462530
transform 1 0 2700 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_1569
timestamp 1745462530
transform 1 0 2684 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_1570
timestamp 1745462530
transform 1 0 2644 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_1571
timestamp 1745462530
transform 1 0 2612 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_1572
timestamp 1745462530
transform 1 0 2636 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_1573
timestamp 1745462530
transform 1 0 2604 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_1574
timestamp 1745462530
transform 1 0 980 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_1575
timestamp 1745462530
transform 1 0 740 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_1576
timestamp 1745462530
transform 1 0 1388 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_1577
timestamp 1745462530
transform 1 0 1364 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_1578
timestamp 1745462530
transform 1 0 1340 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_1579
timestamp 1745462530
transform 1 0 1324 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_1580
timestamp 1745462530
transform 1 0 1308 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_1581
timestamp 1745462530
transform 1 0 1300 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_1582
timestamp 1745462530
transform 1 0 1276 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_1583
timestamp 1745462530
transform 1 0 1292 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_1584
timestamp 1745462530
transform 1 0 1260 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_1585
timestamp 1745462530
transform 1 0 1276 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_1586
timestamp 1745462530
transform 1 0 1268 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_1587
timestamp 1745462530
transform 1 0 1212 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_1588
timestamp 1745462530
transform 1 0 1276 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_1589
timestamp 1745462530
transform 1 0 1260 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_1590
timestamp 1745462530
transform 1 0 1220 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_1591
timestamp 1745462530
transform 1 0 1164 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_1592
timestamp 1745462530
transform 1 0 676 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_1593
timestamp 1745462530
transform 1 0 580 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_1594
timestamp 1745462530
transform 1 0 412 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_1595
timestamp 1745462530
transform 1 0 372 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_1596
timestamp 1745462530
transform 1 0 620 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_1597
timestamp 1745462530
transform 1 0 572 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_1598
timestamp 1745462530
transform 1 0 756 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_1599
timestamp 1745462530
transform 1 0 604 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_1600
timestamp 1745462530
transform 1 0 316 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_1601
timestamp 1745462530
transform 1 0 308 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_1602
timestamp 1745462530
transform 1 0 452 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_1603
timestamp 1745462530
transform 1 0 444 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_1604
timestamp 1745462530
transform 1 0 444 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_1605
timestamp 1745462530
transform 1 0 444 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_1606
timestamp 1745462530
transform 1 0 548 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_1607
timestamp 1745462530
transform 1 0 540 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_1608
timestamp 1745462530
transform 1 0 532 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_1609
timestamp 1745462530
transform 1 0 508 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_1610
timestamp 1745462530
transform 1 0 484 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_1611
timestamp 1745462530
transform 1 0 428 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_1612
timestamp 1745462530
transform 1 0 412 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_1613
timestamp 1745462530
transform 1 0 404 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_1614
timestamp 1745462530
transform 1 0 596 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_1615
timestamp 1745462530
transform 1 0 396 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_1616
timestamp 1745462530
transform 1 0 364 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_1617
timestamp 1745462530
transform 1 0 348 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_1618
timestamp 1745462530
transform 1 0 428 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_1619
timestamp 1745462530
transform 1 0 380 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_1620
timestamp 1745462530
transform 1 0 660 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_1621
timestamp 1745462530
transform 1 0 628 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_1622
timestamp 1745462530
transform 1 0 932 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_1623
timestamp 1745462530
transform 1 0 924 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_1624
timestamp 1745462530
transform 1 0 412 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_1625
timestamp 1745462530
transform 1 0 404 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_1626
timestamp 1745462530
transform 1 0 724 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_1627
timestamp 1745462530
transform 1 0 692 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_1628
timestamp 1745462530
transform 1 0 1372 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_1629
timestamp 1745462530
transform 1 0 1372 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1630
timestamp 1745462530
transform 1 0 1188 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_1631
timestamp 1745462530
transform 1 0 1164 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_1632
timestamp 1745462530
transform 1 0 1452 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_1633
timestamp 1745462530
transform 1 0 1356 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1634
timestamp 1745462530
transform 1 0 1476 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_1635
timestamp 1745462530
transform 1 0 1444 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_1636
timestamp 1745462530
transform 1 0 1444 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_1637
timestamp 1745462530
transform 1 0 1412 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_1638
timestamp 1745462530
transform 1 0 1444 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_1639
timestamp 1745462530
transform 1 0 1428 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_1640
timestamp 1745462530
transform 1 0 1620 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_1641
timestamp 1745462530
transform 1 0 1572 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_1642
timestamp 1745462530
transform 1 0 1612 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_1643
timestamp 1745462530
transform 1 0 1548 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_1644
timestamp 1745462530
transform 1 0 1692 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_1645
timestamp 1745462530
transform 1 0 1692 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_1646
timestamp 1745462530
transform 1 0 2948 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_1647
timestamp 1745462530
transform 1 0 2884 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_1648
timestamp 1745462530
transform 1 0 2884 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_1649
timestamp 1745462530
transform 1 0 3108 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_1650
timestamp 1745462530
transform 1 0 2924 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_1651
timestamp 1745462530
transform 1 0 2900 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_1652
timestamp 1745462530
transform 1 0 2852 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1653
timestamp 1745462530
transform 1 0 2828 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_1654
timestamp 1745462530
transform 1 0 2700 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_1655
timestamp 1745462530
transform 1 0 3028 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_1656
timestamp 1745462530
transform 1 0 2836 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1657
timestamp 1745462530
transform 1 0 2996 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_1658
timestamp 1745462530
transform 1 0 2988 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_1659
timestamp 1745462530
transform 1 0 2924 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_1660
timestamp 1745462530
transform 1 0 2892 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_1661
timestamp 1745462530
transform 1 0 2868 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_1662
timestamp 1745462530
transform 1 0 2860 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_1663
timestamp 1745462530
transform 1 0 3292 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1664
timestamp 1745462530
transform 1 0 3292 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_1665
timestamp 1745462530
transform 1 0 3236 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_1666
timestamp 1745462530
transform 1 0 3212 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_1667
timestamp 1745462530
transform 1 0 3396 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_1668
timestamp 1745462530
transform 1 0 3244 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1669
timestamp 1745462530
transform 1 0 3196 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1670
timestamp 1745462530
transform 1 0 4100 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1671
timestamp 1745462530
transform 1 0 4100 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_1672
timestamp 1745462530
transform 1 0 3388 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1673
timestamp 1745462530
transform 1 0 3228 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_1674
timestamp 1745462530
transform 1 0 3396 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_1675
timestamp 1745462530
transform 1 0 3364 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1676
timestamp 1745462530
transform 1 0 3348 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_1677
timestamp 1745462530
transform 1 0 4172 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_1678
timestamp 1745462530
transform 1 0 4116 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_1679
timestamp 1745462530
transform 1 0 4084 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_1680
timestamp 1745462530
transform 1 0 4036 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_1681
timestamp 1745462530
transform 1 0 3420 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_1682
timestamp 1745462530
transform 1 0 3300 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_1683
timestamp 1745462530
transform 1 0 3396 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_1684
timestamp 1745462530
transform 1 0 3340 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_1685
timestamp 1745462530
transform 1 0 4108 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_1686
timestamp 1745462530
transform 1 0 4036 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_1687
timestamp 1745462530
transform 1 0 3428 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_1688
timestamp 1745462530
transform 1 0 3316 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_1689
timestamp 1745462530
transform 1 0 3540 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_1690
timestamp 1745462530
transform 1 0 3444 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_1691
timestamp 1745462530
transform 1 0 3412 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_1692
timestamp 1745462530
transform 1 0 4092 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_1693
timestamp 1745462530
transform 1 0 4044 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_1694
timestamp 1745462530
transform 1 0 3492 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_1695
timestamp 1745462530
transform 1 0 3356 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_1696
timestamp 1745462530
transform 1 0 3596 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_1697
timestamp 1745462530
transform 1 0 3468 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_1698
timestamp 1745462530
transform 1 0 3428 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_1699
timestamp 1745462530
transform 1 0 4188 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_1700
timestamp 1745462530
transform 1 0 4156 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_1701
timestamp 1745462530
transform 1 0 3308 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_1702
timestamp 1745462530
transform 1 0 3268 0 1 1755
box -2 -2 2 2
use M2_M1  M2_M1_1703
timestamp 1745462530
transform 1 0 3300 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_1704
timestamp 1745462530
transform 1 0 3204 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_1705
timestamp 1745462530
transform 1 0 3028 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_1706
timestamp 1745462530
transform 1 0 2988 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_1707
timestamp 1745462530
transform 1 0 3276 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_1708
timestamp 1745462530
transform 1 0 3260 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_1709
timestamp 1745462530
transform 1 0 3180 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_1710
timestamp 1745462530
transform 1 0 3228 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_1711
timestamp 1745462530
transform 1 0 3196 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_1712
timestamp 1745462530
transform 1 0 3308 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_1713
timestamp 1745462530
transform 1 0 3260 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_1714
timestamp 1745462530
transform 1 0 3220 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_1715
timestamp 1745462530
transform 1 0 3268 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_1716
timestamp 1745462530
transform 1 0 3204 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_1717
timestamp 1745462530
transform 1 0 3204 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_1718
timestamp 1745462530
transform 1 0 3172 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_1719
timestamp 1745462530
transform 1 0 2772 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_1720
timestamp 1745462530
transform 1 0 2748 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_1721
timestamp 1745462530
transform 1 0 2820 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_1722
timestamp 1745462530
transform 1 0 2764 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_1723
timestamp 1745462530
transform 1 0 2676 0 1 3115
box -2 -2 2 2
use M2_M1  M2_M1_1724
timestamp 1745462530
transform 1 0 2620 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_1725
timestamp 1745462530
transform 1 0 2604 0 1 3115
box -2 -2 2 2
use M2_M1  M2_M1_1726
timestamp 1745462530
transform 1 0 2820 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_1727
timestamp 1745462530
transform 1 0 2788 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_1728
timestamp 1745462530
transform 1 0 1620 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_1729
timestamp 1745462530
transform 1 0 1580 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_1730
timestamp 1745462530
transform 1 0 1580 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_1731
timestamp 1745462530
transform 1 0 1540 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1732
timestamp 1745462530
transform 1 0 1572 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_1733
timestamp 1745462530
transform 1 0 1532 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_1734
timestamp 1745462530
transform 1 0 1468 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_1735
timestamp 1745462530
transform 1 0 1460 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_1736
timestamp 1745462530
transform 1 0 1452 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_1737
timestamp 1745462530
transform 1 0 1444 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_1738
timestamp 1745462530
transform 1 0 1404 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_1739
timestamp 1745462530
transform 1 0 1388 0 1 2585
box -2 -2 2 2
use M2_M1  M2_M1_1740
timestamp 1745462530
transform 1 0 1388 0 1 2395
box -2 -2 2 2
use M2_M1  M2_M1_1741
timestamp 1745462530
transform 1 0 1372 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_1742
timestamp 1745462530
transform 1 0 1372 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_1743
timestamp 1745462530
transform 1 0 1420 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_1744
timestamp 1745462530
transform 1 0 1340 0 1 2285
box -2 -2 2 2
use M2_M1  M2_M1_1745
timestamp 1745462530
transform 1 0 740 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_1746
timestamp 1745462530
transform 1 0 652 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_1747
timestamp 1745462530
transform 1 0 292 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_1748
timestamp 1745462530
transform 1 0 204 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_1749
timestamp 1745462530
transform 1 0 612 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_1750
timestamp 1745462530
transform 1 0 604 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_1751
timestamp 1745462530
transform 1 0 772 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_1752
timestamp 1745462530
transform 1 0 724 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_1753
timestamp 1745462530
transform 1 0 244 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_1754
timestamp 1745462530
transform 1 0 204 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_1755
timestamp 1745462530
transform 1 0 956 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_1756
timestamp 1745462530
transform 1 0 948 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_1757
timestamp 1745462530
transform 1 0 700 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_1758
timestamp 1745462530
transform 1 0 228 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_1759
timestamp 1745462530
transform 1 0 196 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_1760
timestamp 1745462530
transform 1 0 204 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_1761
timestamp 1745462530
transform 1 0 204 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_1762
timestamp 1745462530
transform 1 0 556 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_1763
timestamp 1745462530
transform 1 0 484 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_1764
timestamp 1745462530
transform 1 0 316 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_1765
timestamp 1745462530
transform 1 0 204 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_1766
timestamp 1745462530
transform 1 0 444 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_1767
timestamp 1745462530
transform 1 0 420 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_1768
timestamp 1745462530
transform 1 0 596 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_1769
timestamp 1745462530
transform 1 0 564 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_1770
timestamp 1745462530
transform 1 0 532 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_1771
timestamp 1745462530
transform 1 0 444 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_1772
timestamp 1745462530
transform 1 0 516 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_1773
timestamp 1745462530
transform 1 0 516 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_1774
timestamp 1745462530
transform 1 0 844 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_1775
timestamp 1745462530
transform 1 0 804 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_1776
timestamp 1745462530
transform 1 0 1132 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_1777
timestamp 1745462530
transform 1 0 1116 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1778
timestamp 1745462530
transform 1 0 1076 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_1779
timestamp 1745462530
transform 1 0 1068 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_1780
timestamp 1745462530
transform 1 0 1060 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_1781
timestamp 1745462530
transform 1 0 1004 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1782
timestamp 1745462530
transform 1 0 1388 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_1783
timestamp 1745462530
transform 1 0 1268 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_1784
timestamp 1745462530
transform 1 0 1220 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_1785
timestamp 1745462530
transform 1 0 1084 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_1786
timestamp 1745462530
transform 1 0 1284 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_1787
timestamp 1745462530
transform 1 0 1252 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_1788
timestamp 1745462530
transform 1 0 1252 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_1789
timestamp 1745462530
transform 1 0 1340 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_1790
timestamp 1745462530
transform 1 0 1308 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_1791
timestamp 1745462530
transform 1 0 1444 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_1792
timestamp 1745462530
transform 1 0 1404 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_1793
timestamp 1745462530
transform 1 0 1436 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_1794
timestamp 1745462530
transform 1 0 1396 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_1795
timestamp 1745462530
transform 1 0 2052 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_1796
timestamp 1745462530
transform 1 0 2012 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_1797
timestamp 1745462530
transform 1 0 2788 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_1798
timestamp 1745462530
transform 1 0 2764 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_1799
timestamp 1745462530
transform 1 0 2756 0 1 585
box -2 -2 2 2
use M2_M1  M2_M1_1800
timestamp 1745462530
transform 1 0 2740 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_1801
timestamp 1745462530
transform 1 0 2732 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_1802
timestamp 1745462530
transform 1 0 2708 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_1803
timestamp 1745462530
transform 1 0 2772 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_1804
timestamp 1745462530
transform 1 0 2772 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_1805
timestamp 1745462530
transform 1 0 2740 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_1806
timestamp 1745462530
transform 1 0 2716 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1807
timestamp 1745462530
transform 1 0 2660 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_1808
timestamp 1745462530
transform 1 0 2652 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_1809
timestamp 1745462530
transform 1 0 2796 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_1810
timestamp 1745462530
transform 1 0 2732 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1811
timestamp 1745462530
transform 1 0 2700 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1812
timestamp 1745462530
transform 1 0 3060 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_1813
timestamp 1745462530
transform 1 0 3028 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_1814
timestamp 1745462530
transform 1 0 2756 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_1815
timestamp 1745462530
transform 1 0 2748 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_1816
timestamp 1745462530
transform 1 0 3612 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_1817
timestamp 1745462530
transform 1 0 3588 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_1818
timestamp 1745462530
transform 1 0 3292 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_1819
timestamp 1745462530
transform 1 0 3612 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_1820
timestamp 1745462530
transform 1 0 3564 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_1821
timestamp 1745462530
transform 1 0 3564 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_1822
timestamp 1745462530
transform 1 0 3772 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_1823
timestamp 1745462530
transform 1 0 3692 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_1824
timestamp 1745462530
transform 1 0 3692 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_1825
timestamp 1745462530
transform 1 0 3676 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_1826
timestamp 1745462530
transform 1 0 3676 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_1827
timestamp 1745462530
transform 1 0 3676 0 1 345
box -2 -2 2 2
use M2_M1  M2_M1_1828
timestamp 1745462530
transform 1 0 4348 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_1829
timestamp 1745462530
transform 1 0 4268 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_1830
timestamp 1745462530
transform 1 0 4252 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_1831
timestamp 1745462530
transform 1 0 4212 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_1832
timestamp 1745462530
transform 1 0 4180 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_1833
timestamp 1745462530
transform 1 0 4140 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_1834
timestamp 1745462530
transform 1 0 3636 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_1835
timestamp 1745462530
transform 1 0 3596 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_1836
timestamp 1745462530
transform 1 0 4244 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_1837
timestamp 1745462530
transform 1 0 3780 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_1838
timestamp 1745462530
transform 1 0 3588 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_1839
timestamp 1745462530
transform 1 0 3708 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_1840
timestamp 1745462530
transform 1 0 3676 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_1841
timestamp 1745462530
transform 1 0 4244 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_1842
timestamp 1745462530
transform 1 0 3788 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_1843
timestamp 1745462530
transform 1 0 3620 0 1 1885
box -2 -2 2 2
use M2_M1  M2_M1_1844
timestamp 1745462530
transform 1 0 3804 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_1845
timestamp 1745462530
transform 1 0 3740 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_1846
timestamp 1745462530
transform 1 0 3740 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_1847
timestamp 1745462530
transform 1 0 4324 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_1848
timestamp 1745462530
transform 1 0 4316 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_1849
timestamp 1745462530
transform 1 0 3604 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_1850
timestamp 1745462530
transform 1 0 3572 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1851
timestamp 1745462530
transform 1 0 3700 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_1852
timestamp 1745462530
transform 1 0 3620 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_1853
timestamp 1745462530
transform 1 0 3588 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_1854
timestamp 1745462530
transform 1 0 3724 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_1855
timestamp 1745462530
transform 1 0 3692 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_1856
timestamp 1745462530
transform 1 0 3652 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_1857
timestamp 1745462530
transform 1 0 3612 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_1858
timestamp 1745462530
transform 1 0 3612 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_1859
timestamp 1745462530
transform 1 0 3564 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_1860
timestamp 1745462530
transform 1 0 3556 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_1861
timestamp 1745462530
transform 1 0 3684 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_1862
timestamp 1745462530
transform 1 0 3612 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_1863
timestamp 1745462530
transform 1 0 3548 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_1864
timestamp 1745462530
transform 1 0 3644 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_1865
timestamp 1745462530
transform 1 0 3572 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_1866
timestamp 1745462530
transform 1 0 3532 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_1867
timestamp 1745462530
transform 1 0 3500 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_1868
timestamp 1745462530
transform 1 0 3492 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_1869
timestamp 1745462530
transform 1 0 3556 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_1870
timestamp 1745462530
transform 1 0 3524 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_1871
timestamp 1745462530
transform 1 0 3508 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_1872
timestamp 1745462530
transform 1 0 3460 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_1873
timestamp 1745462530
transform 1 0 3452 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_1874
timestamp 1745462530
transform 1 0 3332 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_1875
timestamp 1745462530
transform 1 0 3268 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_1876
timestamp 1745462530
transform 1 0 3244 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_1877
timestamp 1745462530
transform 1 0 3164 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_1878
timestamp 1745462530
transform 1 0 3164 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_1879
timestamp 1745462530
transform 1 0 3508 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_1880
timestamp 1745462530
transform 1 0 3476 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_1881
timestamp 1745462530
transform 1 0 3420 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_1882
timestamp 1745462530
transform 1 0 3404 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_1883
timestamp 1745462530
transform 1 0 3356 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_1884
timestamp 1745462530
transform 1 0 3284 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_1885
timestamp 1745462530
transform 1 0 3284 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_1886
timestamp 1745462530
transform 1 0 3268 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_1887
timestamp 1745462530
transform 1 0 3220 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_1888
timestamp 1745462530
transform 1 0 3204 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_1889
timestamp 1745462530
transform 1 0 2796 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_1890
timestamp 1745462530
transform 1 0 2636 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_1891
timestamp 1745462530
transform 1 0 2588 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_1892
timestamp 1745462530
transform 1 0 2524 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_1893
timestamp 1745462530
transform 1 0 2476 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_1894
timestamp 1745462530
transform 1 0 2476 0 1 3345
box -2 -2 2 2
use M2_M1  M2_M1_1895
timestamp 1745462530
transform 1 0 2468 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_1896
timestamp 1745462530
transform 1 0 2468 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_1897
timestamp 1745462530
transform 1 0 2420 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_1898
timestamp 1745462530
transform 1 0 2868 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_1899
timestamp 1745462530
transform 1 0 2868 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_1900
timestamp 1745462530
transform 1 0 2860 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_1901
timestamp 1745462530
transform 1 0 2796 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_1902
timestamp 1745462530
transform 1 0 2772 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_1903
timestamp 1745462530
transform 1 0 2764 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_1904
timestamp 1745462530
transform 1 0 2740 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_1905
timestamp 1745462530
transform 1 0 2716 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_1906
timestamp 1745462530
transform 1 0 2700 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_1907
timestamp 1745462530
transform 1 0 2692 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_1908
timestamp 1745462530
transform 1 0 3076 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_1909
timestamp 1745462530
transform 1 0 3036 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_1910
timestamp 1745462530
transform 1 0 2988 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_1911
timestamp 1745462530
transform 1 0 2988 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_1912
timestamp 1745462530
transform 1 0 2916 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_1913
timestamp 1745462530
transform 1 0 3044 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_1914
timestamp 1745462530
transform 1 0 3036 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_1915
timestamp 1745462530
transform 1 0 3012 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_1916
timestamp 1745462530
transform 1 0 2972 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_1917
timestamp 1745462530
transform 1 0 2940 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_1918
timestamp 1745462530
transform 1 0 2900 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_1919
timestamp 1745462530
transform 1 0 2892 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_1920
timestamp 1745462530
transform 1 0 2884 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_1921
timestamp 1745462530
transform 1 0 2868 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_1922
timestamp 1745462530
transform 1 0 2852 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_1923
timestamp 1745462530
transform 1 0 3564 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_1924
timestamp 1745462530
transform 1 0 3548 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_1925
timestamp 1745462530
transform 1 0 3500 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_1926
timestamp 1745462530
transform 1 0 3484 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_1927
timestamp 1745462530
transform 1 0 3484 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_1928
timestamp 1745462530
transform 1 0 3364 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_1929
timestamp 1745462530
transform 1 0 3324 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_1930
timestamp 1745462530
transform 1 0 3228 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_1931
timestamp 1745462530
transform 1 0 3212 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_1932
timestamp 1745462530
transform 1 0 3196 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_1933
timestamp 1745462530
transform 1 0 3468 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_1934
timestamp 1745462530
transform 1 0 3436 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_1935
timestamp 1745462530
transform 1 0 3380 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_1936
timestamp 1745462530
transform 1 0 3356 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_1937
timestamp 1745462530
transform 1 0 3196 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_1938
timestamp 1745462530
transform 1 0 3188 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_1939
timestamp 1745462530
transform 1 0 3124 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_1940
timestamp 1745462530
transform 1 0 3108 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_1941
timestamp 1745462530
transform 1 0 3108 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_1942
timestamp 1745462530
transform 1 0 2812 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_1943
timestamp 1745462530
transform 1 0 2572 0 1 3395
box -2 -2 2 2
use M2_M1  M2_M1_1944
timestamp 1745462530
transform 1 0 2572 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_1945
timestamp 1745462530
transform 1 0 2540 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_1946
timestamp 1745462530
transform 1 0 2540 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_1947
timestamp 1745462530
transform 1 0 2532 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_1948
timestamp 1745462530
transform 1 0 2516 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_1949
timestamp 1745462530
transform 1 0 2444 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_1950
timestamp 1745462530
transform 1 0 2436 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_1951
timestamp 1745462530
transform 1 0 2396 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_1952
timestamp 1745462530
transform 1 0 2652 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_1953
timestamp 1745462530
transform 1 0 2564 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_1954
timestamp 1745462530
transform 1 0 1876 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_1955
timestamp 1745462530
transform 1 0 1868 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_1956
timestamp 1745462530
transform 1 0 1828 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_1957
timestamp 1745462530
transform 1 0 1772 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_1958
timestamp 1745462530
transform 1 0 1724 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_1959
timestamp 1745462530
transform 1 0 1700 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_1960
timestamp 1745462530
transform 1 0 1860 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_1961
timestamp 1745462530
transform 1 0 1812 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_1962
timestamp 1745462530
transform 1 0 1772 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_1963
timestamp 1745462530
transform 1 0 1772 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_1964
timestamp 1745462530
transform 1 0 1756 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_1965
timestamp 1745462530
transform 1 0 1748 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_1966
timestamp 1745462530
transform 1 0 2620 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_1967
timestamp 1745462530
transform 1 0 2580 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_1968
timestamp 1745462530
transform 1 0 2532 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_1969
timestamp 1745462530
transform 1 0 2500 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_1970
timestamp 1745462530
transform 1 0 2052 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_1971
timestamp 1745462530
transform 1 0 2020 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_1972
timestamp 1745462530
transform 1 0 2652 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_1973
timestamp 1745462530
transform 1 0 2612 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_1974
timestamp 1745462530
transform 1 0 2588 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_1975
timestamp 1745462530
transform 1 0 2476 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_1976
timestamp 1745462530
transform 1 0 2084 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_1977
timestamp 1745462530
transform 1 0 2060 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_1978
timestamp 1745462530
transform 1 0 1932 0 1 2625
box -2 -2 2 2
use M2_M1  M2_M1_1979
timestamp 1745462530
transform 1 0 1892 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_1980
timestamp 1745462530
transform 1 0 1612 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_1981
timestamp 1745462530
transform 1 0 1596 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_1982
timestamp 1745462530
transform 1 0 1556 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_1983
timestamp 1745462530
transform 1 0 1508 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_1984
timestamp 1745462530
transform 1 0 1484 0 1 3595
box -2 -2 2 2
use M2_M1  M2_M1_1985
timestamp 1745462530
transform 1 0 3580 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_1986
timestamp 1745462530
transform 1 0 3580 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_1987
timestamp 1745462530
transform 1 0 3556 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_1988
timestamp 1745462530
transform 1 0 3460 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_1989
timestamp 1745462530
transform 1 0 3076 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_1990
timestamp 1745462530
transform 1 0 2700 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_1991
timestamp 1745462530
transform 1 0 2636 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_1992
timestamp 1745462530
transform 1 0 2372 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_1993
timestamp 1745462530
transform 1 0 2260 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_1994
timestamp 1745462530
transform 1 0 2100 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_1995
timestamp 1745462530
transform 1 0 3524 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_1996
timestamp 1745462530
transform 1 0 3476 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_1997
timestamp 1745462530
transform 1 0 3460 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_1998
timestamp 1745462530
transform 1 0 3244 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_1999
timestamp 1745462530
transform 1 0 3036 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_2000
timestamp 1745462530
transform 1 0 2764 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_2001
timestamp 1745462530
transform 1 0 2668 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_2002
timestamp 1745462530
transform 1 0 2324 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_2003
timestamp 1745462530
transform 1 0 2156 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_2004
timestamp 1745462530
transform 1 0 1828 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_2005
timestamp 1745462530
transform 1 0 1988 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_2006
timestamp 1745462530
transform 1 0 1980 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_2007
timestamp 1745462530
transform 1 0 1924 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_2008
timestamp 1745462530
transform 1 0 2020 0 1 2505
box -2 -2 2 2
use M2_M1  M2_M1_2009
timestamp 1745462530
transform 1 0 2020 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_2010
timestamp 1745462530
transform 1 0 1988 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_2011
timestamp 1745462530
transform 1 0 1924 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_2012
timestamp 1745462530
transform 1 0 2004 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_2013
timestamp 1745462530
transform 1 0 1980 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_2014
timestamp 1745462530
transform 1 0 1836 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_2015
timestamp 1745462530
transform 1 0 1828 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_2016
timestamp 1745462530
transform 1 0 1820 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_2017
timestamp 1745462530
transform 1 0 1732 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_2018
timestamp 1745462530
transform 1 0 1852 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_2019
timestamp 1745462530
transform 1 0 1748 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_2020
timestamp 1745462530
transform 1 0 1716 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_2021
timestamp 1745462530
transform 1 0 700 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_2022
timestamp 1745462530
transform 1 0 628 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_2023
timestamp 1745462530
transform 1 0 396 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_2024
timestamp 1745462530
transform 1 0 364 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_2025
timestamp 1745462530
transform 1 0 660 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_2026
timestamp 1745462530
transform 1 0 604 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_2027
timestamp 1745462530
transform 1 0 572 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_2028
timestamp 1745462530
transform 1 0 716 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_2029
timestamp 1745462530
transform 1 0 644 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_2030
timestamp 1745462530
transform 1 0 236 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_2031
timestamp 1745462530
transform 1 0 204 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_2032
timestamp 1745462530
transform 1 0 988 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_2033
timestamp 1745462530
transform 1 0 908 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_2034
timestamp 1745462530
transform 1 0 844 0 1 2435
box -2 -2 2 2
use M2_M1  M2_M1_2035
timestamp 1745462530
transform 1 0 820 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_2036
timestamp 1745462530
transform 1 0 700 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_2037
timestamp 1745462530
transform 1 0 308 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_2038
timestamp 1745462530
transform 1 0 300 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_2039
timestamp 1745462530
transform 1 0 316 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_2040
timestamp 1745462530
transform 1 0 308 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_2041
timestamp 1745462530
transform 1 0 308 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_2042
timestamp 1745462530
transform 1 0 308 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_2043
timestamp 1745462530
transform 1 0 556 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_2044
timestamp 1745462530
transform 1 0 372 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_2045
timestamp 1745462530
transform 1 0 340 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_2046
timestamp 1745462530
transform 1 0 316 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2047
timestamp 1745462530
transform 1 0 596 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_2048
timestamp 1745462530
transform 1 0 492 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_2049
timestamp 1745462530
transform 1 0 284 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_2050
timestamp 1745462530
transform 1 0 276 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_2051
timestamp 1745462530
transform 1 0 620 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_2052
timestamp 1745462530
transform 1 0 492 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_2053
timestamp 1745462530
transform 1 0 476 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_2054
timestamp 1745462530
transform 1 0 732 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_2055
timestamp 1745462530
transform 1 0 700 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_2056
timestamp 1745462530
transform 1 0 876 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_2057
timestamp 1745462530
transform 1 0 868 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_2058
timestamp 1745462530
transform 1 0 516 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_2059
timestamp 1745462530
transform 1 0 508 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_2060
timestamp 1745462530
transform 1 0 708 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_2061
timestamp 1745462530
transform 1 0 676 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_2062
timestamp 1745462530
transform 1 0 1628 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_2063
timestamp 1745462530
transform 1 0 1628 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_2064
timestamp 1745462530
transform 1 0 1516 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_2065
timestamp 1745462530
transform 1 0 1508 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_2066
timestamp 1745462530
transform 1 0 1700 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_2067
timestamp 1745462530
transform 1 0 1612 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_2068
timestamp 1745462530
transform 1 0 1708 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_2069
timestamp 1745462530
transform 1 0 1700 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_2070
timestamp 1745462530
transform 1 0 1660 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_2071
timestamp 1745462530
transform 1 0 1652 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_2072
timestamp 1745462530
transform 1 0 1756 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_2073
timestamp 1745462530
transform 1 0 1700 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_2074
timestamp 1745462530
transform 1 0 1684 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_2075
timestamp 1745462530
transform 1 0 1748 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_2076
timestamp 1745462530
transform 1 0 1716 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_2077
timestamp 1745462530
transform 1 0 1812 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_2078
timestamp 1745462530
transform 1 0 1764 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_2079
timestamp 1745462530
transform 1 0 1860 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_2080
timestamp 1745462530
transform 1 0 1820 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2081
timestamp 1745462530
transform 1 0 1860 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_2082
timestamp 1745462530
transform 1 0 1764 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_2083
timestamp 1745462530
transform 1 0 2964 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_2084
timestamp 1745462530
transform 1 0 2924 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_2085
timestamp 1745462530
transform 1 0 2892 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_2086
timestamp 1745462530
transform 1 0 3060 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_2087
timestamp 1745462530
transform 1 0 2876 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_2088
timestamp 1745462530
transform 1 0 2988 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_2089
timestamp 1745462530
transform 1 0 2956 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_2090
timestamp 1745462530
transform 1 0 2892 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_2091
timestamp 1745462530
transform 1 0 2956 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_2092
timestamp 1745462530
transform 1 0 2940 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_2093
timestamp 1745462530
transform 1 0 3916 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_2094
timestamp 1745462530
transform 1 0 3780 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_2095
timestamp 1745462530
transform 1 0 3380 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_2096
timestamp 1745462530
transform 1 0 3356 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_2097
timestamp 1745462530
transform 1 0 3908 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_2098
timestamp 1745462530
transform 1 0 3764 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_2099
timestamp 1745462530
transform 1 0 4172 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_2100
timestamp 1745462530
transform 1 0 4100 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_2101
timestamp 1745462530
transform 1 0 3932 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_2102
timestamp 1745462530
transform 1 0 3932 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_2103
timestamp 1745462530
transform 1 0 4020 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_2104
timestamp 1745462530
transform 1 0 3916 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_2105
timestamp 1745462530
transform 1 0 4180 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_2106
timestamp 1745462530
transform 1 0 4148 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_2107
timestamp 1745462530
transform 1 0 4156 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_2108
timestamp 1745462530
transform 1 0 4124 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_2109
timestamp 1745462530
transform 1 0 3900 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_2110
timestamp 1745462530
transform 1 0 3868 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2111
timestamp 1745462530
transform 1 0 4260 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_2112
timestamp 1745462530
transform 1 0 4132 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_2113
timestamp 1745462530
transform 1 0 4052 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_2114
timestamp 1745462530
transform 1 0 3900 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_2115
timestamp 1745462530
transform 1 0 3916 0 1 1785
box -2 -2 2 2
use M2_M1  M2_M1_2116
timestamp 1745462530
transform 1 0 3884 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_2117
timestamp 1745462530
transform 1 0 4268 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_2118
timestamp 1745462530
transform 1 0 4204 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_2119
timestamp 1745462530
transform 1 0 4068 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_2120
timestamp 1745462530
transform 1 0 3932 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_2121
timestamp 1745462530
transform 1 0 3916 0 1 1985
box -2 -2 2 2
use M2_M1  M2_M1_2122
timestamp 1745462530
transform 1 0 3916 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_2123
timestamp 1745462530
transform 1 0 4244 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_2124
timestamp 1745462530
transform 1 0 4212 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_2125
timestamp 1745462530
transform 1 0 4212 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_2126
timestamp 1745462530
transform 1 0 4148 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_2127
timestamp 1745462530
transform 1 0 4116 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_2128
timestamp 1745462530
transform 1 0 4132 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_2129
timestamp 1745462530
transform 1 0 4108 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_2130
timestamp 1745462530
transform 1 0 4100 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_2131
timestamp 1745462530
transform 1 0 4204 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_2132
timestamp 1745462530
transform 1 0 4196 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_2133
timestamp 1745462530
transform 1 0 4244 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_2134
timestamp 1745462530
transform 1 0 4236 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_2135
timestamp 1745462530
transform 1 0 4180 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_2136
timestamp 1745462530
transform 1 0 4260 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_2137
timestamp 1745462530
transform 1 0 4252 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_2138
timestamp 1745462530
transform 1 0 4164 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_2139
timestamp 1745462530
transform 1 0 4132 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_2140
timestamp 1745462530
transform 1 0 4124 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_2141
timestamp 1745462530
transform 1 0 2908 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_2142
timestamp 1745462530
transform 1 0 2892 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_2143
timestamp 1745462530
transform 1 0 1124 0 1 3825
box -2 -2 2 2
use M2_M1  M2_M1_2144
timestamp 1745462530
transform 1 0 1124 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_2145
timestamp 1745462530
transform 1 0 1124 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_2146
timestamp 1745462530
transform 1 0 3380 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_2147
timestamp 1745462530
transform 1 0 3356 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2148
timestamp 1745462530
transform 1 0 3332 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_2149
timestamp 1745462530
transform 1 0 3100 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_2150
timestamp 1745462530
transform 1 0 3052 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_2151
timestamp 1745462530
transform 1 0 2884 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_2152
timestamp 1745462530
transform 1 0 2492 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_2153
timestamp 1745462530
transform 1 0 2484 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_2154
timestamp 1745462530
transform 1 0 2436 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_2155
timestamp 1745462530
transform 1 0 2876 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_2156
timestamp 1745462530
transform 1 0 2868 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_2157
timestamp 1745462530
transform 1 0 3124 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_2158
timestamp 1745462530
transform 1 0 3116 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_2159
timestamp 1745462530
transform 1 0 3660 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_2160
timestamp 1745462530
transform 1 0 3628 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_2161
timestamp 1745462530
transform 1 0 3636 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_2162
timestamp 1745462530
transform 1 0 3628 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_2163
timestamp 1745462530
transform 1 0 3628 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_2164
timestamp 1745462530
transform 1 0 3620 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_2165
timestamp 1745462530
transform 1 0 3276 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_2166
timestamp 1745462530
transform 1 0 3260 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_2167
timestamp 1745462530
transform 1 0 2420 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_2168
timestamp 1745462530
transform 1 0 2404 0 1 4005
box -2 -2 2 2
use M2_M1  M2_M1_2169
timestamp 1745462530
transform 1 0 2260 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_2170
timestamp 1745462530
transform 1 0 2244 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_2171
timestamp 1745462530
transform 1 0 3268 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2172
timestamp 1745462530
transform 1 0 3260 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_2173
timestamp 1745462530
transform 1 0 3252 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2174
timestamp 1745462530
transform 1 0 3164 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_2175
timestamp 1745462530
transform 1 0 3004 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_2176
timestamp 1745462530
transform 1 0 2788 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_2177
timestamp 1745462530
transform 1 0 2444 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2178
timestamp 1745462530
transform 1 0 2396 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_2179
timestamp 1745462530
transform 1 0 2356 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_2180
timestamp 1745462530
transform 1 0 2772 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_2181
timestamp 1745462530
transform 1 0 2740 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_2182
timestamp 1745462530
transform 1 0 3052 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_2183
timestamp 1745462530
transform 1 0 3044 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_2184
timestamp 1745462530
transform 1 0 3516 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_2185
timestamp 1745462530
transform 1 0 3476 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_2186
timestamp 1745462530
transform 1 0 3412 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_2187
timestamp 1745462530
transform 1 0 3380 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_2188
timestamp 1745462530
transform 1 0 3532 0 1 4005
box -2 -2 2 2
use M2_M1  M2_M1_2189
timestamp 1745462530
transform 1 0 3500 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_2190
timestamp 1745462530
transform 1 0 3220 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_2191
timestamp 1745462530
transform 1 0 3204 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_2192
timestamp 1745462530
transform 1 0 2444 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_2193
timestamp 1745462530
transform 1 0 2436 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_2194
timestamp 1745462530
transform 1 0 2212 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_2195
timestamp 1745462530
transform 1 0 2204 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_2196
timestamp 1745462530
transform 1 0 3556 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2197
timestamp 1745462530
transform 1 0 3516 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2198
timestamp 1745462530
transform 1 0 3476 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2199
timestamp 1745462530
transform 1 0 3428 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2200
timestamp 1745462530
transform 1 0 2892 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2201
timestamp 1745462530
transform 1 0 2724 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2202
timestamp 1745462530
transform 1 0 2580 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_2203
timestamp 1745462530
transform 1 0 2532 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2204
timestamp 1745462530
transform 1 0 2484 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2205
timestamp 1745462530
transform 1 0 2964 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_2206
timestamp 1745462530
transform 1 0 2948 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_2207
timestamp 1745462530
transform 1 0 4332 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_2208
timestamp 1745462530
transform 1 0 4292 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_2209
timestamp 1745462530
transform 1 0 4244 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_2210
timestamp 1745462530
transform 1 0 4204 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_2211
timestamp 1745462530
transform 1 0 4260 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_2212
timestamp 1745462530
transform 1 0 4220 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2213
timestamp 1745462530
transform 1 0 3988 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_2214
timestamp 1745462530
transform 1 0 3956 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_2215
timestamp 1745462530
transform 1 0 2012 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_2216
timestamp 1745462530
transform 1 0 1980 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_2217
timestamp 1745462530
transform 1 0 2044 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_2218
timestamp 1745462530
transform 1 0 2012 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_2219
timestamp 1745462530
transform 1 0 3332 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_2220
timestamp 1745462530
transform 1 0 3292 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_2221
timestamp 1745462530
transform 1 0 3268 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_2222
timestamp 1745462530
transform 1 0 3212 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_2223
timestamp 1745462530
transform 1 0 2876 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_2224
timestamp 1745462530
transform 1 0 2860 0 1 3235
box -2 -2 2 2
use M2_M1  M2_M1_2225
timestamp 1745462530
transform 1 0 2684 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_2226
timestamp 1745462530
transform 1 0 2596 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_2227
timestamp 1745462530
transform 1 0 2412 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_2228
timestamp 1745462530
transform 1 0 2412 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_2229
timestamp 1745462530
transform 1 0 1748 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_2230
timestamp 1745462530
transform 1 0 1740 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_2231
timestamp 1745462530
transform 1 0 4236 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_2232
timestamp 1745462530
transform 1 0 4196 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_2233
timestamp 1745462530
transform 1 0 4252 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_2234
timestamp 1745462530
transform 1 0 4204 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_2235
timestamp 1745462530
transform 1 0 4076 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_2236
timestamp 1745462530
transform 1 0 4060 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_2237
timestamp 1745462530
transform 1 0 3852 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_2238
timestamp 1745462530
transform 1 0 3812 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_2239
timestamp 1745462530
transform 1 0 1596 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_2240
timestamp 1745462530
transform 1 0 1588 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_2241
timestamp 1745462530
transform 1 0 1628 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_2242
timestamp 1745462530
transform 1 0 1620 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_2243
timestamp 1745462530
transform 1 0 2756 0 1 3025
box -2 -2 2 2
use M2_M1  M2_M1_2244
timestamp 1745462530
transform 1 0 2708 0 1 3025
box -2 -2 2 2
use M2_M1  M2_M1_2245
timestamp 1745462530
transform 1 0 2676 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_2246
timestamp 1745462530
transform 1 0 2556 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_2247
timestamp 1745462530
transform 1 0 3492 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_2248
timestamp 1745462530
transform 1 0 3444 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_2249
timestamp 1745462530
transform 1 0 3388 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_2250
timestamp 1745462530
transform 1 0 3348 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_2251
timestamp 1745462530
transform 1 0 2916 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_2252
timestamp 1745462530
transform 1 0 2756 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_2253
timestamp 1745462530
transform 1 0 2748 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_2254
timestamp 1745462530
transform 1 0 2564 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_2255
timestamp 1745462530
transform 1 0 2500 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_2256
timestamp 1745462530
transform 1 0 2716 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_2257
timestamp 1745462530
transform 1 0 2708 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_2258
timestamp 1745462530
transform 1 0 2892 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_2259
timestamp 1745462530
transform 1 0 2884 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_2260
timestamp 1745462530
transform 1 0 4100 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_2261
timestamp 1745462530
transform 1 0 4060 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_2262
timestamp 1745462530
transform 1 0 4076 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_2263
timestamp 1745462530
transform 1 0 4036 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2264
timestamp 1745462530
transform 1 0 4172 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2265
timestamp 1745462530
transform 1 0 4164 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_2266
timestamp 1745462530
transform 1 0 3996 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_2267
timestamp 1745462530
transform 1 0 3956 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2268
timestamp 1745462530
transform 1 0 2052 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2269
timestamp 1745462530
transform 1 0 2044 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_2270
timestamp 1745462530
transform 1 0 1972 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_2271
timestamp 1745462530
transform 1 0 1956 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_2272
timestamp 1745462530
transform 1 0 3468 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_2273
timestamp 1745462530
transform 1 0 3468 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_2274
timestamp 1745462530
transform 1 0 3412 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_2275
timestamp 1745462530
transform 1 0 3348 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_2276
timestamp 1745462530
transform 1 0 2844 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_2277
timestamp 1745462530
transform 1 0 2756 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_2278
timestamp 1745462530
transform 1 0 2748 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_2279
timestamp 1745462530
transform 1 0 2540 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_2280
timestamp 1745462530
transform 1 0 2508 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_2281
timestamp 1745462530
transform 1 0 2500 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_2282
timestamp 1745462530
transform 1 0 1908 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_2283
timestamp 1745462530
transform 1 0 1892 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_2284
timestamp 1745462530
transform 1 0 1820 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_2285
timestamp 1745462530
transform 1 0 1812 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_2286
timestamp 1745462530
transform 1 0 4252 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_2287
timestamp 1745462530
transform 1 0 4212 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_2288
timestamp 1745462530
transform 1 0 4252 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_2289
timestamp 1745462530
transform 1 0 4204 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2290
timestamp 1745462530
transform 1 0 4060 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_2291
timestamp 1745462530
transform 1 0 4020 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_2292
timestamp 1745462530
transform 1 0 3980 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_2293
timestamp 1745462530
transform 1 0 3948 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_2294
timestamp 1745462530
transform 1 0 1700 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_2295
timestamp 1745462530
transform 1 0 1692 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_2296
timestamp 1745462530
transform 1 0 1684 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_2297
timestamp 1745462530
transform 1 0 1676 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_2298
timestamp 1745462530
transform 1 0 3556 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2299
timestamp 1745462530
transform 1 0 3540 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_2300
timestamp 1745462530
transform 1 0 3500 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_2301
timestamp 1745462530
transform 1 0 3444 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_2302
timestamp 1745462530
transform 1 0 2956 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_2303
timestamp 1745462530
transform 1 0 2732 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_2304
timestamp 1745462530
transform 1 0 2692 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_2305
timestamp 1745462530
transform 1 0 2604 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_2306
timestamp 1745462530
transform 1 0 2548 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_2307
timestamp 1745462530
transform 1 0 2700 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_2308
timestamp 1745462530
transform 1 0 2676 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_2309
timestamp 1745462530
transform 1 0 3012 0 1 4005
box -2 -2 2 2
use M2_M1  M2_M1_2310
timestamp 1745462530
transform 1 0 2972 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_2311
timestamp 1745462530
transform 1 0 3788 0 1 4005
box -2 -2 2 2
use M2_M1  M2_M1_2312
timestamp 1745462530
transform 1 0 3756 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_2313
timestamp 1745462530
transform 1 0 3892 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_2314
timestamp 1745462530
transform 1 0 3884 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_2315
timestamp 1745462530
transform 1 0 3716 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_2316
timestamp 1745462530
transform 1 0 3660 0 1 3945
box -2 -2 2 2
use M2_M1  M2_M1_2317
timestamp 1745462530
transform 1 0 3740 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_2318
timestamp 1745462530
transform 1 0 3700 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_2319
timestamp 1745462530
transform 1 0 2524 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_2320
timestamp 1745462530
transform 1 0 2516 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_2321
timestamp 1745462530
transform 1 0 2324 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_2322
timestamp 1745462530
transform 1 0 2316 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_2323
timestamp 1745462530
transform 1 0 3220 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_2324
timestamp 1745462530
transform 1 0 3204 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_2325
timestamp 1745462530
transform 1 0 3164 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_2326
timestamp 1745462530
transform 1 0 3116 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_2327
timestamp 1745462530
transform 1 0 3036 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_2328
timestamp 1745462530
transform 1 0 2852 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_2329
timestamp 1745462530
transform 1 0 2644 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_2330
timestamp 1745462530
transform 1 0 2620 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_2331
timestamp 1745462530
transform 1 0 2596 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_2332
timestamp 1745462530
transform 1 0 3156 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_2333
timestamp 1745462530
transform 1 0 3148 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_2334
timestamp 1745462530
transform 1 0 3404 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_2335
timestamp 1745462530
transform 1 0 3396 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_2336
timestamp 1745462530
transform 1 0 3332 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_2337
timestamp 1745462530
transform 1 0 3324 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_2338
timestamp 1745462530
transform 1 0 3388 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_2339
timestamp 1745462530
transform 1 0 3380 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_2340
timestamp 1745462530
transform 1 0 3196 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_2341
timestamp 1745462530
transform 1 0 3188 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_2342
timestamp 1745462530
transform 1 0 2420 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_2343
timestamp 1745462530
transform 1 0 2412 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_2344
timestamp 1745462530
transform 1 0 2108 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_2345
timestamp 1745462530
transform 1 0 2100 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_2346
timestamp 1745462530
transform 1 0 2828 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_2347
timestamp 1745462530
transform 1 0 2812 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_2348
timestamp 1745462530
transform 1 0 2796 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_2349
timestamp 1745462530
transform 1 0 2764 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_2350
timestamp 1745462530
transform 1 0 3140 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_2351
timestamp 1745462530
transform 1 0 3044 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_2352
timestamp 1745462530
transform 1 0 3028 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_2353
timestamp 1745462530
transform 1 0 1748 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_2354
timestamp 1745462530
transform 1 0 1612 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_2355
timestamp 1745462530
transform 1 0 1588 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_2356
timestamp 1745462530
transform 1 0 2804 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_2357
timestamp 1745462530
transform 1 0 2804 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_2358
timestamp 1745462530
transform 1 0 2772 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_2359
timestamp 1745462530
transform 1 0 1724 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_2360
timestamp 1745462530
transform 1 0 1580 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_2361
timestamp 1745462530
transform 1 0 1556 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_2362
timestamp 1745462530
transform 1 0 3860 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_2363
timestamp 1745462530
transform 1 0 3844 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_2364
timestamp 1745462530
transform 1 0 4084 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_2365
timestamp 1745462530
transform 1 0 4052 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_2366
timestamp 1745462530
transform 1 0 4252 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_2367
timestamp 1745462530
transform 1 0 4236 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_2368
timestamp 1745462530
transform 1 0 4244 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_2369
timestamp 1745462530
transform 1 0 4228 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_2370
timestamp 1745462530
transform 1 0 1820 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_2371
timestamp 1745462530
transform 1 0 1708 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_2372
timestamp 1745462530
transform 1 0 1684 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_2373
timestamp 1745462530
transform 1 0 1860 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_2374
timestamp 1745462530
transform 1 0 1756 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_2375
timestamp 1745462530
transform 1 0 1732 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_2376
timestamp 1745462530
transform 1 0 1716 0 1 3835
box -2 -2 2 2
use M2_M1  M2_M1_2377
timestamp 1745462530
transform 1 0 1668 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_2378
timestamp 1745462530
transform 1 0 1500 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_2379
timestamp 1745462530
transform 1 0 1692 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_2380
timestamp 1745462530
transform 1 0 1684 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_2381
timestamp 1745462530
transform 1 0 1612 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_2382
timestamp 1745462530
transform 1 0 4012 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_2383
timestamp 1745462530
transform 1 0 3972 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_2384
timestamp 1745462530
transform 1 0 4068 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_2385
timestamp 1745462530
transform 1 0 4052 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_2386
timestamp 1745462530
transform 1 0 4252 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2387
timestamp 1745462530
transform 1 0 4236 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2388
timestamp 1745462530
transform 1 0 4260 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_2389
timestamp 1745462530
transform 1 0 4244 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_2390
timestamp 1745462530
transform 1 0 1804 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_2391
timestamp 1745462530
transform 1 0 1804 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_2392
timestamp 1745462530
transform 1 0 1788 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_2393
timestamp 1745462530
transform 1 0 1884 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_2394
timestamp 1745462530
transform 1 0 1836 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_2395
timestamp 1745462530
transform 1 0 1836 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_2396
timestamp 1745462530
transform 1 0 2044 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_2397
timestamp 1745462530
transform 1 0 1948 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_2398
timestamp 1745462530
transform 1 0 1948 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_2399
timestamp 1745462530
transform 1 0 2076 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_2400
timestamp 1745462530
transform 1 0 2036 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_2401
timestamp 1745462530
transform 1 0 2036 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2402
timestamp 1745462530
transform 1 0 4004 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2403
timestamp 1745462530
transform 1 0 3988 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2404
timestamp 1745462530
transform 1 0 4156 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2405
timestamp 1745462530
transform 1 0 4148 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_2406
timestamp 1745462530
transform 1 0 4084 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2407
timestamp 1745462530
transform 1 0 4068 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2408
timestamp 1745462530
transform 1 0 4108 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_2409
timestamp 1745462530
transform 1 0 4092 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_2410
timestamp 1745462530
transform 1 0 2876 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_2411
timestamp 1745462530
transform 1 0 2876 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_2412
timestamp 1745462530
transform 1 0 2660 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_2413
timestamp 1745462530
transform 1 0 2700 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_2414
timestamp 1745462530
transform 1 0 2564 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_2415
timestamp 1745462530
transform 1 0 2564 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_2416
timestamp 1745462530
transform 1 0 2068 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_2417
timestamp 1745462530
transform 1 0 2036 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_2418
timestamp 1745462530
transform 1 0 2020 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_2419
timestamp 1745462530
transform 1 0 2044 0 1 3745
box -2 -2 2 2
use M2_M1  M2_M1_2420
timestamp 1745462530
transform 1 0 2012 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_2421
timestamp 1745462530
transform 1 0 2004 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_2422
timestamp 1745462530
transform 1 0 3980 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_2423
timestamp 1745462530
transform 1 0 3916 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2424
timestamp 1745462530
transform 1 0 4268 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2425
timestamp 1745462530
transform 1 0 4252 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2426
timestamp 1745462530
transform 1 0 4252 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_2427
timestamp 1745462530
transform 1 0 4236 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_2428
timestamp 1745462530
transform 1 0 4340 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_2429
timestamp 1745462530
transform 1 0 4324 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_2430
timestamp 1745462530
transform 1 0 2940 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_2431
timestamp 1745462530
transform 1 0 2900 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_2432
timestamp 1745462530
transform 1 0 2628 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_2433
timestamp 1745462530
transform 1 0 2612 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_2434
timestamp 1745462530
transform 1 0 2556 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_2435
timestamp 1745462530
transform 1 0 2524 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_2436
timestamp 1745462530
transform 1 0 2308 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_2437
timestamp 1745462530
transform 1 0 2276 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_2438
timestamp 1745462530
transform 1 0 2252 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_2439
timestamp 1745462530
transform 1 0 2508 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_2440
timestamp 1745462530
transform 1 0 2460 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_2441
timestamp 1745462530
transform 1 0 2364 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_2442
timestamp 1745462530
transform 1 0 3748 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_2443
timestamp 1745462530
transform 1 0 3732 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_2444
timestamp 1745462530
transform 1 0 3452 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_2445
timestamp 1745462530
transform 1 0 3724 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_2446
timestamp 1745462530
transform 1 0 3708 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_2447
timestamp 1745462530
transform 1 0 3588 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_2448
timestamp 1745462530
transform 1 0 3908 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_2449
timestamp 1745462530
transform 1 0 3876 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_2450
timestamp 1745462530
transform 1 0 3556 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_2451
timestamp 1745462530
transform 1 0 3796 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_2452
timestamp 1745462530
transform 1 0 3780 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_2453
timestamp 1745462530
transform 1 0 3572 0 1 4005
box -2 -2 2 2
use M2_M1  M2_M1_2454
timestamp 1745462530
transform 1 0 3068 0 1 4005
box -2 -2 2 2
use M2_M1  M2_M1_2455
timestamp 1745462530
transform 1 0 3004 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_2456
timestamp 1745462530
transform 1 0 3004 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_2457
timestamp 1745462530
transform 1 0 2692 0 1 4005
box -2 -2 2 2
use M2_M1  M2_M1_2458
timestamp 1745462530
transform 1 0 2684 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_2459
timestamp 1745462530
transform 1 0 2668 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_2460
timestamp 1745462530
transform 1 0 2228 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_2461
timestamp 1745462530
transform 1 0 2196 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_2462
timestamp 1745462530
transform 1 0 2172 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_2463
timestamp 1745462530
transform 1 0 2428 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_2464
timestamp 1745462530
transform 1 0 2388 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_2465
timestamp 1745462530
transform 1 0 2348 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_2466
timestamp 1745462530
transform 1 0 3420 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_2467
timestamp 1745462530
transform 1 0 3308 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_2468
timestamp 1745462530
transform 1 0 3196 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_2469
timestamp 1745462530
transform 1 0 3596 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_2470
timestamp 1745462530
transform 1 0 3540 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_2471
timestamp 1745462530
transform 1 0 3524 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_2472
timestamp 1745462530
transform 1 0 3532 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_2473
timestamp 1745462530
transform 1 0 3492 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_2474
timestamp 1745462530
transform 1 0 3404 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_2475
timestamp 1745462530
transform 1 0 3564 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_2476
timestamp 1745462530
transform 1 0 3556 0 1 4005
box -2 -2 2 2
use M2_M1  M2_M1_2477
timestamp 1745462530
transform 1 0 3508 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_2478
timestamp 1745462530
transform 1 0 3084 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_2479
timestamp 1745462530
transform 1 0 3036 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_2480
timestamp 1745462530
transform 1 0 3028 0 1 4005
box -2 -2 2 2
use M2_M1  M2_M1_2481
timestamp 1745462530
transform 1 0 2780 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_2482
timestamp 1745462530
transform 1 0 2764 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_2483
timestamp 1745462530
transform 1 0 2660 0 1 4005
box -2 -2 2 2
use M2_M1  M2_M1_2484
timestamp 1745462530
transform 1 0 2236 0 1 4005
box -2 -2 2 2
use M2_M1  M2_M1_2485
timestamp 1745462530
transform 1 0 2236 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_2486
timestamp 1745462530
transform 1 0 2396 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_2487
timestamp 1745462530
transform 1 0 2348 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_2488
timestamp 1745462530
transform 1 0 2348 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_2489
timestamp 1745462530
transform 1 0 3284 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_2490
timestamp 1745462530
transform 1 0 3268 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_2491
timestamp 1745462530
transform 1 0 3252 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_2492
timestamp 1745462530
transform 1 0 3692 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_2493
timestamp 1745462530
transform 1 0 3612 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_2494
timestamp 1745462530
transform 1 0 3564 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_2495
timestamp 1745462530
transform 1 0 3628 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_2496
timestamp 1745462530
transform 1 0 3620 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_2497
timestamp 1745462530
transform 1 0 3484 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_2498
timestamp 1745462530
transform 1 0 3668 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_2499
timestamp 1745462530
transform 1 0 3652 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_2500
timestamp 1745462530
transform 1 0 3508 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_2501
timestamp 1745462530
transform 1 0 3108 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_2502
timestamp 1745462530
transform 1 0 3092 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_2503
timestamp 1745462530
transform 1 0 3076 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_2504
timestamp 1745462530
transform 1 0 2860 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_2505
timestamp 1745462530
transform 1 0 2788 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_2506
timestamp 1745462530
transform 1 0 2708 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_2507
timestamp 1745462530
transform 1 0 2124 0 1 4005
box -2 -2 2 2
use M2_M1  M2_M1_2508
timestamp 1745462530
transform 1 0 2100 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_2509
timestamp 1745462530
transform 1 0 2092 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_2510
timestamp 1745462530
transform 1 0 2404 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_2511
timestamp 1745462530
transform 1 0 2372 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_2512
timestamp 1745462530
transform 1 0 2332 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_2513
timestamp 1745462530
transform 1 0 3244 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_2514
timestamp 1745462530
transform 1 0 3228 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_2515
timestamp 1745462530
transform 1 0 3180 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_2516
timestamp 1745462530
transform 1 0 3516 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_2517
timestamp 1745462530
transform 1 0 3404 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_2518
timestamp 1745462530
transform 1 0 3372 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_2519
timestamp 1745462530
transform 1 0 3468 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_2520
timestamp 1745462530
transform 1 0 3468 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_2521
timestamp 1745462530
transform 1 0 3316 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_2522
timestamp 1745462530
transform 1 0 3484 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_2523
timestamp 1745462530
transform 1 0 3420 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_2524
timestamp 1745462530
transform 1 0 3388 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_2525
timestamp 1745462530
transform 1 0 2268 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_2526
timestamp 1745462530
transform 1 0 2236 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_2527
timestamp 1745462530
transform 1 0 2180 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_2528
timestamp 1745462530
transform 1 0 2180 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_2529
timestamp 1745462530
transform 1 0 2156 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_2530
timestamp 1745462530
transform 1 0 2140 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_2531
timestamp 1745462530
transform 1 0 2132 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_2532
timestamp 1745462530
transform 1 0 452 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_2533
timestamp 1745462530
transform 1 0 428 0 1 4005
box -2 -2 2 2
use M2_M1  M2_M1_2534
timestamp 1745462530
transform 1 0 484 0 1 3915
box -2 -2 2 2
use M2_M1  M2_M1_2535
timestamp 1745462530
transform 1 0 420 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_2536
timestamp 1745462530
transform 1 0 340 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_2537
timestamp 1745462530
transform 1 0 340 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_2538
timestamp 1745462530
transform 1 0 300 0 1 4025
box -2 -2 2 2
use M2_M1  M2_M1_2539
timestamp 1745462530
transform 1 0 476 0 1 3995
box -2 -2 2 2
use M2_M1  M2_M1_2540
timestamp 1745462530
transform 1 0 452 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_2541
timestamp 1745462530
transform 1 0 452 0 1 4025
box -2 -2 2 2
use M2_M1  M2_M1_2542
timestamp 1745462530
transform 1 0 316 0 1 4025
box -2 -2 2 2
use M2_M1  M2_M1_2543
timestamp 1745462530
transform 1 0 1292 0 1 3825
box -2 -2 2 2
use M2_M1  M2_M1_2544
timestamp 1745462530
transform 1 0 1228 0 1 3825
box -2 -2 2 2
use M2_M1  M2_M1_2545
timestamp 1745462530
transform 1 0 468 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_2546
timestamp 1745462530
transform 1 0 204 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_2547
timestamp 1745462530
transform 1 0 164 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_2548
timestamp 1745462530
transform 1 0 1580 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2549
timestamp 1745462530
transform 1 0 1540 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_2550
timestamp 1745462530
transform 1 0 1404 0 1 3625
box -2 -2 2 2
use M2_M1  M2_M1_2551
timestamp 1745462530
transform 1 0 1372 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_2552
timestamp 1745462530
transform 1 0 1372 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2553
timestamp 1745462530
transform 1 0 1316 0 1 3825
box -2 -2 2 2
use M2_M1  M2_M1_2554
timestamp 1745462530
transform 1 0 1276 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_2555
timestamp 1745462530
transform 1 0 1556 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_2556
timestamp 1745462530
transform 1 0 1556 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_2557
timestamp 1745462530
transform 1 0 1508 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_2558
timestamp 1745462530
transform 1 0 1500 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_2559
timestamp 1745462530
transform 1 0 1476 0 1 3745
box -2 -2 2 2
use M2_M1  M2_M1_2560
timestamp 1745462530
transform 1 0 1444 0 1 3625
box -2 -2 2 2
use M2_M1  M2_M1_2561
timestamp 1745462530
transform 1 0 1340 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2562
timestamp 1745462530
transform 1 0 1460 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2563
timestamp 1745462530
transform 1 0 1444 0 1 3435
box -2 -2 2 2
use M2_M1  M2_M1_2564
timestamp 1745462530
transform 1 0 588 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_2565
timestamp 1745462530
transform 1 0 572 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_2566
timestamp 1745462530
transform 1 0 564 0 1 4005
box -2 -2 2 2
use M2_M1  M2_M1_2567
timestamp 1745462530
transform 1 0 1020 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_2568
timestamp 1745462530
transform 1 0 940 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_2569
timestamp 1745462530
transform 1 0 908 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_2570
timestamp 1745462530
transform 1 0 3884 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_2571
timestamp 1745462530
transform 1 0 3844 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_2572
timestamp 1745462530
transform 1 0 3836 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_2573
timestamp 1745462530
transform 1 0 3796 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_2574
timestamp 1745462530
transform 1 0 3668 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_2575
timestamp 1745462530
transform 1 0 3612 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_2576
timestamp 1745462530
transform 1 0 3516 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_2577
timestamp 1745462530
transform 1 0 3348 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_2578
timestamp 1745462530
transform 1 0 3060 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_2579
timestamp 1745462530
transform 1 0 3020 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_2580
timestamp 1745462530
transform 1 0 2836 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_2581
timestamp 1745462530
transform 1 0 2700 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_2582
timestamp 1745462530
transform 1 0 2324 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_2583
timestamp 1745462530
transform 1 0 2188 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_2584
timestamp 1745462530
transform 1 0 2148 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_2585
timestamp 1745462530
transform 1 0 2044 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_2586
timestamp 1745462530
transform 1 0 1540 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_2587
timestamp 1745462530
transform 1 0 3860 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_2588
timestamp 1745462530
transform 1 0 3828 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_2589
timestamp 1745462530
transform 1 0 3820 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_2590
timestamp 1745462530
transform 1 0 3780 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_2591
timestamp 1745462530
transform 1 0 3652 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_2592
timestamp 1745462530
transform 1 0 3580 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_2593
timestamp 1745462530
transform 1 0 3500 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_2594
timestamp 1745462530
transform 1 0 3332 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_2595
timestamp 1745462530
transform 1 0 3044 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_2596
timestamp 1745462530
transform 1 0 3004 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_2597
timestamp 1745462530
transform 1 0 2820 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_2598
timestamp 1745462530
transform 1 0 2684 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_2599
timestamp 1745462530
transform 1 0 2308 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_2600
timestamp 1745462530
transform 1 0 2172 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_2601
timestamp 1745462530
transform 1 0 2132 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_2602
timestamp 1745462530
transform 1 0 2028 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_2603
timestamp 1745462530
transform 1 0 1388 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_2604
timestamp 1745462530
transform 1 0 1356 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_2605
timestamp 1745462530
transform 1 0 1108 0 1 3995
box -2 -2 2 2
use M2_M1  M2_M1_2606
timestamp 1745462530
transform 1 0 1044 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_2607
timestamp 1745462530
transform 1 0 980 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_2608
timestamp 1745462530
transform 1 0 4148 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_2609
timestamp 1745462530
transform 1 0 4140 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_2610
timestamp 1745462530
transform 1 0 4124 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_2611
timestamp 1745462530
transform 1 0 4124 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_2612
timestamp 1745462530
transform 1 0 4116 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_2613
timestamp 1745462530
transform 1 0 4092 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_2614
timestamp 1745462530
transform 1 0 4004 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_2615
timestamp 1745462530
transform 1 0 3940 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_2616
timestamp 1745462530
transform 1 0 2956 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_2617
timestamp 1745462530
transform 1 0 2932 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_2618
timestamp 1745462530
transform 1 0 2636 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_2619
timestamp 1745462530
transform 1 0 2580 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_2620
timestamp 1745462530
transform 1 0 1988 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_2621
timestamp 1745462530
transform 1 0 1964 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_2622
timestamp 1745462530
transform 1 0 1916 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_2623
timestamp 1745462530
transform 1 0 1876 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_2624
timestamp 1745462530
transform 1 0 1412 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_2625
timestamp 1745462530
transform 1 0 1372 0 1 4115
box -2 -2 2 2
use M2_M1  M2_M1_2626
timestamp 1745462530
transform 1 0 1372 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_2627
timestamp 1745462530
transform 1 0 724 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_2628
timestamp 1745462530
transform 1 0 708 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_2629
timestamp 1745462530
transform 1 0 644 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_2630
timestamp 1745462530
transform 1 0 612 0 1 4115
box -2 -2 2 2
use M2_M1  M2_M1_2631
timestamp 1745462530
transform 1 0 620 0 1 4145
box -2 -2 2 2
use M2_M1  M2_M1_2632
timestamp 1745462530
transform 1 0 580 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_2633
timestamp 1745462530
transform 1 0 580 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_2634
timestamp 1745462530
transform 1 0 772 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_2635
timestamp 1745462530
transform 1 0 764 0 1 3945
box -2 -2 2 2
use M2_M1  M2_M1_2636
timestamp 1745462530
transform 1 0 748 0 1 3945
box -2 -2 2 2
use M2_M1  M2_M1_2637
timestamp 1745462530
transform 1 0 132 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_2638
timestamp 1745462530
transform 1 0 116 0 1 4115
box -2 -2 2 2
use M2_M1  M2_M1_2639
timestamp 1745462530
transform 1 0 116 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_2640
timestamp 1745462530
transform 1 0 92 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_2641
timestamp 1745462530
transform 1 0 92 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_2642
timestamp 1745462530
transform 1 0 204 0 1 4235
box -2 -2 2 2
use M2_M1  M2_M1_2643
timestamp 1745462530
transform 1 0 180 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_2644
timestamp 1745462530
transform 1 0 124 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_2645
timestamp 1745462530
transform 1 0 212 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_2646
timestamp 1745462530
transform 1 0 196 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_2647
timestamp 1745462530
transform 1 0 188 0 1 4225
box -2 -2 2 2
use M2_M1  M2_M1_2648
timestamp 1745462530
transform 1 0 132 0 1 3795
box -2 -2 2 2
use M2_M1  M2_M1_2649
timestamp 1745462530
transform 1 0 100 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_2650
timestamp 1745462530
transform 1 0 196 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_2651
timestamp 1745462530
transform 1 0 172 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_2652
timestamp 1745462530
transform 1 0 196 0 1 4005
box -2 -2 2 2
use M2_M1  M2_M1_2653
timestamp 1745462530
transform 1 0 132 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_2654
timestamp 1745462530
transform 1 0 116 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_2655
timestamp 1745462530
transform 1 0 836 0 1 4005
box -2 -2 2 2
use M2_M1  M2_M1_2656
timestamp 1745462530
transform 1 0 780 0 1 4115
box -2 -2 2 2
use M2_M1  M2_M1_2657
timestamp 1745462530
transform 1 0 700 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_2658
timestamp 1745462530
transform 1 0 396 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_2659
timestamp 1745462530
transform 1 0 316 0 1 4005
box -2 -2 2 2
use M2_M1  M2_M1_2660
timestamp 1745462530
transform 1 0 308 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_2661
timestamp 1745462530
transform 1 0 228 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_2662
timestamp 1745462530
transform 1 0 324 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_2663
timestamp 1745462530
transform 1 0 284 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_2664
timestamp 1745462530
transform 1 0 676 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_2665
timestamp 1745462530
transform 1 0 644 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_2666
timestamp 1745462530
transform 1 0 628 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_2667
timestamp 1745462530
transform 1 0 964 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_2668
timestamp 1745462530
transform 1 0 892 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_2669
timestamp 1745462530
transform 1 0 1004 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_2670
timestamp 1745462530
transform 1 0 932 0 1 4115
box -2 -2 2 2
use M2_M1  M2_M1_2671
timestamp 1745462530
transform 1 0 828 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_2672
timestamp 1745462530
transform 1 0 724 0 1 4115
box -2 -2 2 2
use M2_M1  M2_M1_2673
timestamp 1745462530
transform 1 0 700 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_2674
timestamp 1745462530
transform 1 0 684 0 1 4195
box -2 -2 2 2
use M2_M1  M2_M1_2675
timestamp 1745462530
transform 1 0 700 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_2676
timestamp 1745462530
transform 1 0 684 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_2677
timestamp 1745462530
transform 1 0 1292 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_2678
timestamp 1745462530
transform 1 0 1276 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_2679
timestamp 1745462530
transform 1 0 1180 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_2680
timestamp 1745462530
transform 1 0 1164 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_2681
timestamp 1745462530
transform 1 0 956 0 1 4005
box -2 -2 2 2
use M2_M1  M2_M1_2682
timestamp 1745462530
transform 1 0 924 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_2683
timestamp 1745462530
transform 1 0 828 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_2684
timestamp 1745462530
transform 1 0 708 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_2685
timestamp 1745462530
transform 1 0 524 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_2686
timestamp 1745462530
transform 1 0 500 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_2687
timestamp 1745462530
transform 1 0 364 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_2688
timestamp 1745462530
transform 1 0 260 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_2689
timestamp 1745462530
transform 1 0 236 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_2690
timestamp 1745462530
transform 1 0 204 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_2691
timestamp 1745462530
transform 1 0 1172 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_2692
timestamp 1745462530
transform 1 0 1172 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_2693
timestamp 1745462530
transform 1 0 852 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_2694
timestamp 1745462530
transform 1 0 740 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_2695
timestamp 1745462530
transform 1 0 700 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_2696
timestamp 1745462530
transform 1 0 636 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_2697
timestamp 1745462530
transform 1 0 604 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_2698
timestamp 1745462530
transform 1 0 580 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_2699
timestamp 1745462530
transform 1 0 516 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_2700
timestamp 1745462530
transform 1 0 500 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_2701
timestamp 1745462530
transform 1 0 500 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_2702
timestamp 1745462530
transform 1 0 460 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_2703
timestamp 1745462530
transform 1 0 428 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_2704
timestamp 1745462530
transform 1 0 380 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_2705
timestamp 1745462530
transform 1 0 1004 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_2706
timestamp 1745462530
transform 1 0 972 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_2707
timestamp 1745462530
transform 1 0 948 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_2708
timestamp 1745462530
transform 1 0 2164 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_2709
timestamp 1745462530
transform 1 0 2164 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_2710
timestamp 1745462530
transform 1 0 908 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_2711
timestamp 1745462530
transform 1 0 2252 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_2712
timestamp 1745462530
transform 1 0 2132 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_2713
timestamp 1745462530
transform 1 0 2084 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_2714
timestamp 1745462530
transform 1 0 1612 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_2715
timestamp 1745462530
transform 1 0 2580 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_2716
timestamp 1745462530
transform 1 0 2556 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_2717
timestamp 1745462530
transform 1 0 2228 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_2718
timestamp 1745462530
transform 1 0 2220 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_2719
timestamp 1745462530
transform 1 0 2012 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_2720
timestamp 1745462530
transform 1 0 1972 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_2721
timestamp 1745462530
transform 1 0 1948 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_2722
timestamp 1745462530
transform 1 0 1948 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_2723
timestamp 1745462530
transform 1 0 2276 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_2724
timestamp 1745462530
transform 1 0 2244 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_2725
timestamp 1745462530
transform 1 0 2004 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_2726
timestamp 1745462530
transform 1 0 1948 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_2727
timestamp 1745462530
transform 1 0 2204 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2728
timestamp 1745462530
transform 1 0 2124 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_2729
timestamp 1745462530
transform 1 0 2100 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_2730
timestamp 1745462530
transform 1 0 1572 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_2731
timestamp 1745462530
transform 1 0 1980 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_2732
timestamp 1745462530
transform 1 0 1436 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2733
timestamp 1745462530
transform 1 0 1332 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_2734
timestamp 1745462530
transform 1 0 1332 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_2735
timestamp 1745462530
transform 1 0 2268 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_2736
timestamp 1745462530
transform 1 0 2188 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_2737
timestamp 1745462530
transform 1 0 2180 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2738
timestamp 1745462530
transform 1 0 2164 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_2739
timestamp 1745462530
transform 1 0 2124 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_2740
timestamp 1745462530
transform 1 0 1804 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_2741
timestamp 1745462530
transform 1 0 1796 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_2742
timestamp 1745462530
transform 1 0 4028 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_2743
timestamp 1745462530
transform 1 0 4004 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_2744
timestamp 1745462530
transform 1 0 3956 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_2745
timestamp 1745462530
transform 1 0 3948 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_2746
timestamp 1745462530
transform 1 0 3956 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_2747
timestamp 1745462530
transform 1 0 3948 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_2748
timestamp 1745462530
transform 1 0 3892 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_2749
timestamp 1745462530
transform 1 0 3868 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_2750
timestamp 1745462530
transform 1 0 1636 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_2751
timestamp 1745462530
transform 1 0 1612 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_2752
timestamp 1745462530
transform 1 0 1348 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_2753
timestamp 1745462530
transform 1 0 1324 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_2754
timestamp 1745462530
transform 1 0 4292 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_2755
timestamp 1745462530
transform 1 0 4284 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_2756
timestamp 1745462530
transform 1 0 4284 0 1 4005
box -2 -2 2 2
use M2_M1  M2_M1_2757
timestamp 1745462530
transform 1 0 4180 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_2758
timestamp 1745462530
transform 1 0 1652 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_2759
timestamp 1745462530
transform 1 0 1628 0 1 4005
box -2 -2 2 2
use M2_M1  M2_M1_2760
timestamp 1745462530
transform 1 0 1556 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_2761
timestamp 1745462530
transform 1 0 1404 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_2762
timestamp 1745462530
transform 1 0 1364 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_2763
timestamp 1745462530
transform 1 0 1308 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_2764
timestamp 1745462530
transform 1 0 1260 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_2765
timestamp 1745462530
transform 1 0 1220 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_2766
timestamp 1745462530
transform 1 0 1212 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_2767
timestamp 1745462530
transform 1 0 1116 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_2768
timestamp 1745462530
transform 1 0 1108 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_2769
timestamp 1745462530
transform 1 0 1020 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_2770
timestamp 1745462530
transform 1 0 940 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_2771
timestamp 1745462530
transform 1 0 820 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_2772
timestamp 1745462530
transform 1 0 748 0 1 4005
box -2 -2 2 2
use M2_M1  M2_M1_2773
timestamp 1745462530
transform 1 0 732 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_2774
timestamp 1745462530
transform 1 0 644 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_2775
timestamp 1745462530
transform 1 0 3356 0 1 4005
box -2 -2 2 2
use M2_M1  M2_M1_2776
timestamp 1745462530
transform 1 0 3252 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_2777
timestamp 1745462530
transform 1 0 3244 0 1 4005
box -2 -2 2 2
use M2_M1  M2_M1_2778
timestamp 1745462530
transform 1 0 3124 0 1 4005
box -2 -2 2 2
use M2_M1  M2_M1_2779
timestamp 1745462530
transform 1 0 2460 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_2780
timestamp 1745462530
transform 1 0 2068 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_2781
timestamp 1745462530
transform 1 0 1340 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_2782
timestamp 1745462530
transform 1 0 996 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_2783
timestamp 1745462530
transform 1 0 868 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_2784
timestamp 1745462530
transform 1 0 556 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_2785
timestamp 1745462530
transform 1 0 380 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_2786
timestamp 1745462530
transform 1 0 356 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_2787
timestamp 1745462530
transform 1 0 348 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_2788
timestamp 1745462530
transform 1 0 244 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_2789
timestamp 1745462530
transform 1 0 3884 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_2790
timestamp 1745462530
transform 1 0 3836 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_2791
timestamp 1745462530
transform 1 0 3724 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_2792
timestamp 1745462530
transform 1 0 3636 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_2793
timestamp 1745462530
transform 1 0 3636 0 1 4005
box -2 -2 2 2
use M2_M1  M2_M1_2794
timestamp 1745462530
transform 1 0 3540 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_2795
timestamp 1745462530
transform 1 0 3388 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_2796
timestamp 1745462530
transform 1 0 3292 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_2797
timestamp 1745462530
transform 1 0 3100 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_2798
timestamp 1745462530
transform 1 0 3084 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_2799
timestamp 1745462530
transform 1 0 2812 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_2800
timestamp 1745462530
transform 1 0 2748 0 1 4005
box -2 -2 2 2
use M2_M1  M2_M1_2801
timestamp 1745462530
transform 1 0 2460 0 1 4005
box -2 -2 2 2
use M2_M1  M2_M1_2802
timestamp 1745462530
transform 1 0 2252 0 1 4005
box -2 -2 2 2
use M2_M1  M2_M1_2803
timestamp 1745462530
transform 1 0 3924 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_2804
timestamp 1745462530
transform 1 0 3908 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_2805
timestamp 1745462530
transform 1 0 3844 0 1 4005
box -2 -2 2 2
use M2_M1  M2_M1_2806
timestamp 1745462530
transform 1 0 3764 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_2807
timestamp 1745462530
transform 1 0 3732 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_2808
timestamp 1745462530
transform 1 0 3196 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_2809
timestamp 1745462530
transform 1 0 2908 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_2810
timestamp 1745462530
transform 1 0 2868 0 1 4005
box -2 -2 2 2
use M2_M1  M2_M1_2811
timestamp 1745462530
transform 1 0 2724 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_2812
timestamp 1745462530
transform 1 0 2556 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_2813
timestamp 1745462530
transform 1 0 2444 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_2814
timestamp 1745462530
transform 1 0 2348 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_2815
timestamp 1745462530
transform 1 0 2212 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_2816
timestamp 1745462530
transform 1 0 2036 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_2817
timestamp 1745462530
transform 1 0 4292 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_2818
timestamp 1745462530
transform 1 0 4292 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_2819
timestamp 1745462530
transform 1 0 4284 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_2820
timestamp 1745462530
transform 1 0 4284 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_2821
timestamp 1745462530
transform 1 0 4164 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_2822
timestamp 1745462530
transform 1 0 4116 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_2823
timestamp 1745462530
transform 1 0 4044 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_2824
timestamp 1745462530
transform 1 0 3988 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_2825
timestamp 1745462530
transform 1 0 3932 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_2826
timestamp 1745462530
transform 1 0 2916 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_2827
timestamp 1745462530
transform 1 0 2580 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_2828
timestamp 1745462530
transform 1 0 1980 0 1 4005
box -2 -2 2 2
use M2_M1  M2_M1_2829
timestamp 1745462530
transform 1 0 1916 0 1 3955
box -2 -2 2 2
use M2_M1  M2_M1_2830
timestamp 1745462530
transform 1 0 1916 0 1 3905
box -2 -2 2 2
use M2_M1  M2_M1_2831
timestamp 1745462530
transform 1 0 1916 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_2832
timestamp 1745462530
transform 1 0 1908 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_2833
timestamp 1745462530
transform 1 0 4292 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_2834
timestamp 1745462530
transform 1 0 4292 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_2835
timestamp 1745462530
transform 1 0 4284 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_2836
timestamp 1745462530
transform 1 0 4284 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_2837
timestamp 1745462530
transform 1 0 4100 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_2838
timestamp 1745462530
transform 1 0 4020 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_2839
timestamp 1745462530
transform 1 0 3924 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_2840
timestamp 1745462530
transform 1 0 1932 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_2841
timestamp 1745462530
transform 1 0 1828 0 1 4005
box -2 -2 2 2
use M2_M1  M2_M1_2842
timestamp 1745462530
transform 1 0 1748 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_2843
timestamp 1745462530
transform 1 0 1620 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_2844
timestamp 1745462530
transform 1 0 1516 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_2845
timestamp 1745462530
transform 1 0 1500 0 1 4005
box -2 -2 2 2
use M2_M1  M2_M1_2846
timestamp 1745462530
transform 1 0 1388 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_2847
timestamp 1745462530
transform 1 0 4292 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_2848
timestamp 1745462530
transform 1 0 4284 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_2849
timestamp 1745462530
transform 1 0 4252 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_2850
timestamp 1745462530
transform 1 0 4188 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_2851
timestamp 1745462530
transform 1 0 4116 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_2852
timestamp 1745462530
transform 1 0 4084 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_2853
timestamp 1745462530
transform 1 0 4068 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_2854
timestamp 1745462530
transform 1 0 3908 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_2855
timestamp 1745462530
transform 1 0 3020 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_2856
timestamp 1745462530
transform 1 0 2892 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_2857
timestamp 1745462530
transform 1 0 2788 0 1 3807
box -2 -2 2 2
use M2_M1  M2_M1_2858
timestamp 1745462530
transform 1 0 2772 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_2859
timestamp 1745462530
transform 1 0 1460 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_2860
timestamp 1745462530
transform 1 0 1348 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_2861
timestamp 1745462530
transform 1 0 4284 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_2862
timestamp 1745462530
transform 1 0 4284 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_2863
timestamp 1745462530
transform 1 0 4244 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_2864
timestamp 1745462530
transform 1 0 4196 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_2865
timestamp 1745462530
transform 1 0 4188 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_2866
timestamp 1745462530
transform 1 0 4164 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_2867
timestamp 1745462530
transform 1 0 4092 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_2868
timestamp 1745462530
transform 1 0 4012 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_2869
timestamp 1745462530
transform 1 0 3996 0 1 3115
box -2 -2 2 2
use M2_M1  M2_M1_2870
timestamp 1745462530
transform 1 0 3996 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_2871
timestamp 1745462530
transform 1 0 3964 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_2872
timestamp 1745462530
transform 1 0 3956 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_2873
timestamp 1745462530
transform 1 0 3196 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_2874
timestamp 1745462530
transform 1 0 3004 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_2875
timestamp 1745462530
transform 1 0 4164 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_2876
timestamp 1745462530
transform 1 0 4140 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_2877
timestamp 1745462530
transform 1 0 4036 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_2878
timestamp 1745462530
transform 1 0 3916 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_2879
timestamp 1745462530
transform 1 0 3348 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_2880
timestamp 1745462530
transform 1 0 3124 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_2881
timestamp 1745462530
transform 1 0 3100 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_2882
timestamp 1745462530
transform 1 0 3004 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_2883
timestamp 1745462530
transform 1 0 2996 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_2884
timestamp 1745462530
transform 1 0 2956 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_2885
timestamp 1745462530
transform 1 0 2908 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_2886
timestamp 1745462530
transform 1 0 2892 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_2887
timestamp 1745462530
transform 1 0 2796 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_2888
timestamp 1745462530
transform 1 0 2156 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_2889
timestamp 1745462530
transform 1 0 1852 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_2890
timestamp 1745462530
transform 1 0 1748 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_2891
timestamp 1745462530
transform 1 0 1748 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_2892
timestamp 1745462530
transform 1 0 1716 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_2893
timestamp 1745462530
transform 1 0 1716 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_2894
timestamp 1745462530
transform 1 0 1708 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_2895
timestamp 1745462530
transform 1 0 1676 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_2896
timestamp 1745462530
transform 1 0 1524 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_2897
timestamp 1745462530
transform 1 0 1356 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_2898
timestamp 1745462530
transform 1 0 732 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_2899
timestamp 1745462530
transform 1 0 692 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_2900
timestamp 1745462530
transform 1 0 572 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_2901
timestamp 1745462530
transform 1 0 572 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_2902
timestamp 1745462530
transform 1 0 548 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_2903
timestamp 1745462530
transform 1 0 1828 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_2904
timestamp 1745462530
transform 1 0 1732 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_2905
timestamp 1745462530
transform 1 0 1724 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_2906
timestamp 1745462530
transform 1 0 1636 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_2907
timestamp 1745462530
transform 1 0 1620 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_2908
timestamp 1745462530
transform 1 0 908 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_2909
timestamp 1745462530
transform 1 0 532 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_2910
timestamp 1745462530
transform 1 0 508 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_2911
timestamp 1745462530
transform 1 0 284 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_2912
timestamp 1745462530
transform 1 0 260 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_2913
timestamp 1745462530
transform 1 0 220 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_2914
timestamp 1745462530
transform 1 0 212 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_2915
timestamp 1745462530
transform 1 0 204 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_2916
timestamp 1745462530
transform 1 0 148 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_2917
timestamp 1745462530
transform 1 0 100 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_2918
timestamp 1745462530
transform 1 0 92 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_2919
timestamp 1745462530
transform 1 0 3716 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_2920
timestamp 1745462530
transform 1 0 3684 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_2921
timestamp 1745462530
transform 1 0 3668 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_2922
timestamp 1745462530
transform 1 0 3604 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_2923
timestamp 1745462530
transform 1 0 3572 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_2924
timestamp 1745462530
transform 1 0 3468 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_2925
timestamp 1745462530
transform 1 0 2964 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_2926
timestamp 1745462530
transform 1 0 2524 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_2927
timestamp 1745462530
transform 1 0 2204 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_2928
timestamp 1745462530
transform 1 0 2084 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_2929
timestamp 1745462530
transform 1 0 2052 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_2930
timestamp 1745462530
transform 1 0 2012 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_2931
timestamp 1745462530
transform 1 0 1940 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_2932
timestamp 1745462530
transform 1 0 1916 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_2933
timestamp 1745462530
transform 1 0 4292 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_2934
timestamp 1745462530
transform 1 0 4292 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_2935
timestamp 1745462530
transform 1 0 4284 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_2936
timestamp 1745462530
transform 1 0 4284 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_2937
timestamp 1745462530
transform 1 0 4284 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_2938
timestamp 1745462530
transform 1 0 4092 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_2939
timestamp 1745462530
transform 1 0 3716 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_2940
timestamp 1745462530
transform 1 0 3644 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_2941
timestamp 1745462530
transform 1 0 3636 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_2942
timestamp 1745462530
transform 1 0 3596 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_2943
timestamp 1745462530
transform 1 0 3548 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_2944
timestamp 1745462530
transform 1 0 2820 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_2945
timestamp 1745462530
transform 1 0 2620 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_2946
timestamp 1745462530
transform 1 0 2292 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_2947
timestamp 1745462530
transform 1 0 3684 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_2948
timestamp 1745462530
transform 1 0 3604 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_2949
timestamp 1745462530
transform 1 0 3572 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_2950
timestamp 1745462530
transform 1 0 3236 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_2951
timestamp 1745462530
transform 1 0 3012 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_2952
timestamp 1745462530
transform 1 0 2820 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_2953
timestamp 1745462530
transform 1 0 2724 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_2954
timestamp 1745462530
transform 1 0 2716 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_2955
timestamp 1745462530
transform 1 0 2708 0 1 995
box -2 -2 2 2
use M2_M1  M2_M1_2956
timestamp 1745462530
transform 1 0 2692 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_2957
timestamp 1745462530
transform 1 0 2684 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_2958
timestamp 1745462530
transform 1 0 2676 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_2959
timestamp 1745462530
transform 1 0 2668 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_2960
timestamp 1745462530
transform 1 0 2556 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_2961
timestamp 1745462530
transform 1 0 2196 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_2962
timestamp 1745462530
transform 1 0 2020 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_2963
timestamp 1745462530
transform 1 0 1356 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_2964
timestamp 1745462530
transform 1 0 1292 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_2965
timestamp 1745462530
transform 1 0 1284 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_2966
timestamp 1745462530
transform 1 0 1252 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_2967
timestamp 1745462530
transform 1 0 1180 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_2968
timestamp 1745462530
transform 1 0 1116 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_2969
timestamp 1745462530
transform 1 0 980 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_2970
timestamp 1745462530
transform 1 0 964 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_2971
timestamp 1745462530
transform 1 0 748 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_2972
timestamp 1745462530
transform 1 0 724 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_2973
timestamp 1745462530
transform 1 0 596 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_2974
timestamp 1745462530
transform 1 0 508 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_2975
timestamp 1745462530
transform 1 0 460 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_2976
timestamp 1745462530
transform 1 0 372 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_2977
timestamp 1745462530
transform 1 0 1380 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_2978
timestamp 1745462530
transform 1 0 1380 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_2979
timestamp 1745462530
transform 1 0 1348 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_2980
timestamp 1745462530
transform 1 0 1340 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_2981
timestamp 1745462530
transform 1 0 980 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_2982
timestamp 1745462530
transform 1 0 484 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_2983
timestamp 1745462530
transform 1 0 476 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_2984
timestamp 1745462530
transform 1 0 268 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_2985
timestamp 1745462530
transform 1 0 92 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_2986
timestamp 1745462530
transform 1 0 92 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_2987
timestamp 1745462530
transform 1 0 92 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_2988
timestamp 1745462530
transform 1 0 92 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_2989
timestamp 1745462530
transform 1 0 84 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_2990
timestamp 1745462530
transform 1 0 84 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_2991
timestamp 1745462530
transform 1 0 3268 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_2992
timestamp 1745462530
transform 1 0 3164 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_2993
timestamp 1745462530
transform 1 0 3132 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_2994
timestamp 1745462530
transform 1 0 3084 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_2995
timestamp 1745462530
transform 1 0 3068 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_2996
timestamp 1745462530
transform 1 0 3060 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_2997
timestamp 1745462530
transform 1 0 2884 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_2998
timestamp 1745462530
transform 1 0 2748 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_2999
timestamp 1745462530
transform 1 0 2684 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_3000
timestamp 1745462530
transform 1 0 2684 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_3001
timestamp 1745462530
transform 1 0 1548 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3002
timestamp 1745462530
transform 1 0 1548 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_3003
timestamp 1745462530
transform 1 0 1524 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_3004
timestamp 1745462530
transform 1 0 1524 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_3005
timestamp 1745462530
transform 1 0 1524 0 1 2395
box -2 -2 2 2
use M2_M1  M2_M1_3006
timestamp 1745462530
transform 1 0 1460 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_3007
timestamp 1745462530
transform 1 0 4212 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_3008
timestamp 1745462530
transform 1 0 4204 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_3009
timestamp 1745462530
transform 1 0 4116 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_3010
timestamp 1745462530
transform 1 0 4116 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3011
timestamp 1745462530
transform 1 0 4076 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_3012
timestamp 1745462530
transform 1 0 3988 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_3013
timestamp 1745462530
transform 1 0 3508 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_3014
timestamp 1745462530
transform 1 0 3452 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_3015
timestamp 1745462530
transform 1 0 3348 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_3016
timestamp 1745462530
transform 1 0 3260 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_3017
timestamp 1745462530
transform 1 0 3260 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_3018
timestamp 1745462530
transform 1 0 3236 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_3019
timestamp 1745462530
transform 1 0 2788 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_3020
timestamp 1745462530
transform 1 0 2228 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_3021
timestamp 1745462530
transform 1 0 3148 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_3022
timestamp 1745462530
transform 1 0 3140 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_3023
timestamp 1745462530
transform 1 0 3116 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_3024
timestamp 1745462530
transform 1 0 3076 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3025
timestamp 1745462530
transform 1 0 3036 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_3026
timestamp 1745462530
transform 1 0 2924 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_3027
timestamp 1745462530
transform 1 0 2908 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_3028
timestamp 1745462530
transform 1 0 2892 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_3029
timestamp 1745462530
transform 1 0 2852 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_3030
timestamp 1745462530
transform 1 0 2724 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_3031
timestamp 1745462530
transform 1 0 2140 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_3032
timestamp 1745462530
transform 1 0 1580 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_3033
timestamp 1745462530
transform 1 0 1556 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_3034
timestamp 1745462530
transform 1 0 1524 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_3035
timestamp 1745462530
transform 1 0 1596 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_3036
timestamp 1745462530
transform 1 0 1572 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_3037
timestamp 1745462530
transform 1 0 1500 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3038
timestamp 1745462530
transform 1 0 1380 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_3039
timestamp 1745462530
transform 1 0 1292 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_3040
timestamp 1745462530
transform 1 0 1036 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_3041
timestamp 1745462530
transform 1 0 924 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_3042
timestamp 1745462530
transform 1 0 692 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_3043
timestamp 1745462530
transform 1 0 572 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_3044
timestamp 1745462530
transform 1 0 468 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_3045
timestamp 1745462530
transform 1 0 452 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_3046
timestamp 1745462530
transform 1 0 444 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_3047
timestamp 1745462530
transform 1 0 388 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_3048
timestamp 1745462530
transform 1 0 308 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_3049
timestamp 1745462530
transform 1 0 1988 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_3050
timestamp 1745462530
transform 1 0 1340 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3051
timestamp 1745462530
transform 1 0 1308 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_3052
timestamp 1745462530
transform 1 0 1284 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_3053
timestamp 1745462530
transform 1 0 1236 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_3054
timestamp 1745462530
transform 1 0 1228 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3055
timestamp 1745462530
transform 1 0 1212 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_3056
timestamp 1745462530
transform 1 0 804 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_3057
timestamp 1745462530
transform 1 0 564 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3058
timestamp 1745462530
transform 1 0 476 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_3059
timestamp 1745462530
transform 1 0 420 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_3060
timestamp 1745462530
transform 1 0 348 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_3061
timestamp 1745462530
transform 1 0 332 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3062
timestamp 1745462530
transform 1 0 188 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3063
timestamp 1745462530
transform 1 0 4292 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3064
timestamp 1745462530
transform 1 0 4292 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_3065
timestamp 1745462530
transform 1 0 4276 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_3066
timestamp 1745462530
transform 1 0 4252 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_3067
timestamp 1745462530
transform 1 0 4164 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_3068
timestamp 1745462530
transform 1 0 4116 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3069
timestamp 1745462530
transform 1 0 3964 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3070
timestamp 1745462530
transform 1 0 3292 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_3071
timestamp 1745462530
transform 1 0 2852 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_3072
timestamp 1745462530
transform 1 0 2788 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_3073
timestamp 1745462530
transform 1 0 2556 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_3074
timestamp 1745462530
transform 1 0 2508 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3075
timestamp 1745462530
transform 1 0 2308 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_3076
timestamp 1745462530
transform 1 0 1124 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3077
timestamp 1745462530
transform 1 0 4292 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_3078
timestamp 1745462530
transform 1 0 4292 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_3079
timestamp 1745462530
transform 1 0 4292 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_3080
timestamp 1745462530
transform 1 0 4292 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_3081
timestamp 1745462530
transform 1 0 4284 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_3082
timestamp 1745462530
transform 1 0 4284 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_3083
timestamp 1745462530
transform 1 0 4276 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_3084
timestamp 1745462530
transform 1 0 4052 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_3085
timestamp 1745462530
transform 1 0 3996 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_3086
timestamp 1745462530
transform 1 0 3804 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_3087
timestamp 1745462530
transform 1 0 3628 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_3088
timestamp 1745462530
transform 1 0 3604 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_3089
timestamp 1745462530
transform 1 0 3460 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_3090
timestamp 1745462530
transform 1 0 2276 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_3091
timestamp 1745462530
transform 1 0 2356 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_3092
timestamp 1745462530
transform 1 0 2228 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_3093
timestamp 1745462530
transform 1 0 2228 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_3094
timestamp 1745462530
transform 1 0 2188 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_3095
timestamp 1745462530
transform 1 0 2172 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_3096
timestamp 1745462530
transform 1 0 2100 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_3097
timestamp 1745462530
transform 1 0 2092 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_3098
timestamp 1745462530
transform 1 0 2068 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_3099
timestamp 1745462530
transform 1 0 1988 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_3100
timestamp 1745462530
transform 1 0 1980 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_3101
timestamp 1745462530
transform 1 0 1900 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_3102
timestamp 1745462530
transform 1 0 1892 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_3103
timestamp 1745462530
transform 1 0 1868 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_3104
timestamp 1745462530
transform 1 0 1820 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_3105
timestamp 1745462530
transform 1 0 1964 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_3106
timestamp 1745462530
transform 1 0 1788 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_3107
timestamp 1745462530
transform 1 0 1788 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_3108
timestamp 1745462530
transform 1 0 1676 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_3109
timestamp 1745462530
transform 1 0 812 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_3110
timestamp 1745462530
transform 1 0 668 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_3111
timestamp 1745462530
transform 1 0 548 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_3112
timestamp 1745462530
transform 1 0 436 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_3113
timestamp 1745462530
transform 1 0 428 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_3114
timestamp 1745462530
transform 1 0 332 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_3115
timestamp 1745462530
transform 1 0 268 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_3116
timestamp 1745462530
transform 1 0 268 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_3117
timestamp 1745462530
transform 1 0 260 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_3118
timestamp 1745462530
transform 1 0 172 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_3119
timestamp 1745462530
transform 1 0 2396 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3120
timestamp 1745462530
transform 1 0 1972 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_3121
timestamp 1745462530
transform 1 0 1724 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_3122
timestamp 1745462530
transform 1 0 1708 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3123
timestamp 1745462530
transform 1 0 1676 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_3124
timestamp 1745462530
transform 1 0 1652 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_3125
timestamp 1745462530
transform 1 0 1644 0 1 2455
box -2 -2 2 2
use M2_M1  M2_M1_3126
timestamp 1745462530
transform 1 0 1628 0 1 2455
box -2 -2 2 2
use M2_M1  M2_M1_3127
timestamp 1745462530
transform 1 0 1604 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_3128
timestamp 1745462530
transform 1 0 1548 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_3129
timestamp 1745462530
transform 1 0 1012 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_3130
timestamp 1745462530
transform 1 0 428 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_3131
timestamp 1745462530
transform 1 0 404 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_3132
timestamp 1745462530
transform 1 0 404 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_3133
timestamp 1745462530
transform 1 0 308 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_3134
timestamp 1745462530
transform 1 0 212 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_3135
timestamp 1745462530
transform 1 0 3988 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_3136
timestamp 1745462530
transform 1 0 3980 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_3137
timestamp 1745462530
transform 1 0 3948 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_3138
timestamp 1745462530
transform 1 0 3908 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_3139
timestamp 1745462530
transform 1 0 3892 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_3140
timestamp 1745462530
transform 1 0 3876 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_3141
timestamp 1745462530
transform 1 0 3876 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_3142
timestamp 1745462530
transform 1 0 3820 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3143
timestamp 1745462530
transform 1 0 3796 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3144
timestamp 1745462530
transform 1 0 3652 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3145
timestamp 1745462530
transform 1 0 3060 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_3146
timestamp 1745462530
transform 1 0 3060 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_3147
timestamp 1745462530
transform 1 0 2572 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_3148
timestamp 1745462530
transform 1 0 2540 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_3149
timestamp 1745462530
transform 1 0 4292 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3150
timestamp 1745462530
transform 1 0 4284 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_3151
timestamp 1745462530
transform 1 0 4284 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_3152
timestamp 1745462530
transform 1 0 4188 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_3153
timestamp 1745462530
transform 1 0 4132 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_3154
timestamp 1745462530
transform 1 0 3844 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_3155
timestamp 1745462530
transform 1 0 3756 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_3156
timestamp 1745462530
transform 1 0 3756 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_3157
timestamp 1745462530
transform 1 0 3708 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_3158
timestamp 1745462530
transform 1 0 3692 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3159
timestamp 1745462530
transform 1 0 3436 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_3160
timestamp 1745462530
transform 1 0 2604 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_3161
timestamp 1745462530
transform 1 0 2572 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_3162
timestamp 1745462530
transform 1 0 2564 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_3163
timestamp 1745462530
transform 1 0 2468 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_3164
timestamp 1745462530
transform 1 0 2460 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_3165
timestamp 1745462530
transform 1 0 2356 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_3166
timestamp 1745462530
transform 1 0 2356 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_3167
timestamp 1745462530
transform 1 0 2340 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_3168
timestamp 1745462530
transform 1 0 2244 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_3169
timestamp 1745462530
transform 1 0 2156 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_3170
timestamp 1745462530
transform 1 0 2156 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_3171
timestamp 1745462530
transform 1 0 2076 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_3172
timestamp 1745462530
transform 1 0 2060 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_3173
timestamp 1745462530
transform 1 0 1988 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_3174
timestamp 1745462530
transform 1 0 1988 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_3175
timestamp 1745462530
transform 1 0 1980 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_3176
timestamp 1745462530
transform 1 0 1972 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_3177
timestamp 1745462530
transform 1 0 1636 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_3178
timestamp 1745462530
transform 1 0 1572 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_3179
timestamp 1745462530
transform 1 0 892 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_3180
timestamp 1745462530
transform 1 0 804 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_3181
timestamp 1745462530
transform 1 0 772 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_3182
timestamp 1745462530
transform 1 0 764 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_3183
timestamp 1745462530
transform 1 0 356 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_3184
timestamp 1745462530
transform 1 0 308 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_3185
timestamp 1745462530
transform 1 0 252 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_3186
timestamp 1745462530
transform 1 0 212 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_3187
timestamp 1745462530
transform 1 0 116 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_3188
timestamp 1745462530
transform 1 0 100 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_3189
timestamp 1745462530
transform 1 0 100 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_3190
timestamp 1745462530
transform 1 0 92 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_3191
timestamp 1745462530
transform 1 0 2844 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_3192
timestamp 1745462530
transform 1 0 2740 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_3193
timestamp 1745462530
transform 1 0 2660 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3194
timestamp 1745462530
transform 1 0 2108 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_3195
timestamp 1745462530
transform 1 0 1980 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_3196
timestamp 1745462530
transform 1 0 1916 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_3197
timestamp 1745462530
transform 1 0 1900 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_3198
timestamp 1745462530
transform 1 0 1884 0 1 2435
box -2 -2 2 2
use M2_M1  M2_M1_3199
timestamp 1745462530
transform 1 0 1884 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_3200
timestamp 1745462530
transform 1 0 1876 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_3201
timestamp 1745462530
transform 1 0 1820 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3202
timestamp 1745462530
transform 1 0 1716 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_3203
timestamp 1745462530
transform 1 0 1012 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3204
timestamp 1745462530
transform 1 0 756 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_3205
timestamp 1745462530
transform 1 0 652 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_3206
timestamp 1745462530
transform 1 0 444 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3207
timestamp 1745462530
transform 1 0 4100 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_3208
timestamp 1745462530
transform 1 0 4076 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_3209
timestamp 1745462530
transform 1 0 3612 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_3210
timestamp 1745462530
transform 1 0 3452 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_3211
timestamp 1745462530
transform 1 0 3436 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_3212
timestamp 1745462530
transform 1 0 3428 0 1 2385
box -2 -2 2 2
use M2_M1  M2_M1_3213
timestamp 1745462530
transform 1 0 3420 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_3214
timestamp 1745462530
transform 1 0 3412 0 1 2385
box -2 -2 2 2
use M2_M1  M2_M1_3215
timestamp 1745462530
transform 1 0 3388 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_3216
timestamp 1745462530
transform 1 0 3372 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3217
timestamp 1745462530
transform 1 0 3364 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_3218
timestamp 1745462530
transform 1 0 3364 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_3219
timestamp 1745462530
transform 1 0 3252 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_3220
timestamp 1745462530
transform 1 0 2676 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_3221
timestamp 1745462530
transform 1 0 2492 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_3222
timestamp 1745462530
transform 1 0 2276 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_3223
timestamp 1745462530
transform 1 0 3996 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3224
timestamp 1745462530
transform 1 0 3956 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_3225
timestamp 1745462530
transform 1 0 3948 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_3226
timestamp 1745462530
transform 1 0 3860 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_3227
timestamp 1745462530
transform 1 0 3484 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_3228
timestamp 1745462530
transform 1 0 3476 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_3229
timestamp 1745462530
transform 1 0 3468 0 1 785
box -2 -2 2 2
use M2_M1  M2_M1_3230
timestamp 1745462530
transform 1 0 3468 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_3231
timestamp 1745462530
transform 1 0 3436 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_3232
timestamp 1745462530
transform 1 0 3412 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_3233
timestamp 1745462530
transform 1 0 3228 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_3234
timestamp 1745462530
transform 1 0 2612 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_3235
timestamp 1745462530
transform 1 0 2596 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_3236
timestamp 1745462530
transform 1 0 2340 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_3237
timestamp 1745462530
transform 1 0 2332 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_3238
timestamp 1745462530
transform 1 0 2204 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_3239
timestamp 1745462530
transform 1 0 2196 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_3240
timestamp 1745462530
transform 1 0 2108 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3241
timestamp 1745462530
transform 1 0 2100 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_3242
timestamp 1745462530
transform 1 0 2092 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_3243
timestamp 1745462530
transform 1 0 2084 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_3244
timestamp 1745462530
transform 1 0 1380 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_3245
timestamp 1745462530
transform 1 0 1316 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_3246
timestamp 1745462530
transform 1 0 1284 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_3247
timestamp 1745462530
transform 1 0 1244 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_3248
timestamp 1745462530
transform 1 0 1196 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_3249
timestamp 1745462530
transform 1 0 1188 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_3250
timestamp 1745462530
transform 1 0 1020 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_3251
timestamp 1745462530
transform 1 0 1012 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_3252
timestamp 1745462530
transform 1 0 980 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_3253
timestamp 1745462530
transform 1 0 924 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_3254
timestamp 1745462530
transform 1 0 860 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_3255
timestamp 1745462530
transform 1 0 812 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_3256
timestamp 1745462530
transform 1 0 796 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_3257
timestamp 1745462530
transform 1 0 652 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_3258
timestamp 1745462530
transform 1 0 132 0 1 1855
box -2 -2 2 2
use M2_M1  M2_M1_3259
timestamp 1745462530
transform 1 0 100 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3260
timestamp 1745462530
transform 1 0 92 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_3261
timestamp 1745462530
transform 1 0 92 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_3262
timestamp 1745462530
transform 1 0 92 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_3263
timestamp 1745462530
transform 1 0 92 0 1 1855
box -2 -2 2 2
use M2_M1  M2_M1_3264
timestamp 1745462530
transform 1 0 92 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_3265
timestamp 1745462530
transform 1 0 92 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_3266
timestamp 1745462530
transform 1 0 92 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_3267
timestamp 1745462530
transform 1 0 92 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_3268
timestamp 1745462530
transform 1 0 92 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_3269
timestamp 1745462530
transform 1 0 1468 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3270
timestamp 1745462530
transform 1 0 1412 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_3271
timestamp 1745462530
transform 1 0 1404 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_3272
timestamp 1745462530
transform 1 0 1148 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_3273
timestamp 1745462530
transform 1 0 1108 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_3274
timestamp 1745462530
transform 1 0 1084 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_3275
timestamp 1745462530
transform 1 0 1052 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_3276
timestamp 1745462530
transform 1 0 1052 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_3277
timestamp 1745462530
transform 1 0 1020 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_3278
timestamp 1745462530
transform 1 0 996 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3279
timestamp 1745462530
transform 1 0 980 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_3280
timestamp 1745462530
transform 1 0 980 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_3281
timestamp 1745462530
transform 1 0 868 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_3282
timestamp 1745462530
transform 1 0 852 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_3283
timestamp 1745462530
transform 1 0 2364 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_3284
timestamp 1745462530
transform 1 0 2284 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3285
timestamp 1745462530
transform 1 0 2268 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_3286
timestamp 1745462530
transform 1 0 2196 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_3287
timestamp 1745462530
transform 1 0 2100 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_3288
timestamp 1745462530
transform 1 0 1996 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_3289
timestamp 1745462530
transform 1 0 1044 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3290
timestamp 1745462530
transform 1 0 1036 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_3291
timestamp 1745462530
transform 1 0 1028 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3292
timestamp 1745462530
transform 1 0 900 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_3293
timestamp 1745462530
transform 1 0 764 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_3294
timestamp 1745462530
transform 1 0 732 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_3295
timestamp 1745462530
transform 1 0 716 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_3296
timestamp 1745462530
transform 1 0 692 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_3297
timestamp 1745462530
transform 1 0 1180 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3298
timestamp 1745462530
transform 1 0 964 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3299
timestamp 1745462530
transform 1 0 692 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3300
timestamp 1745462530
transform 1 0 612 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_3301
timestamp 1745462530
transform 1 0 404 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_3302
timestamp 1745462530
transform 1 0 380 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_3303
timestamp 1745462530
transform 1 0 292 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_3304
timestamp 1745462530
transform 1 0 268 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_3305
timestamp 1745462530
transform 1 0 156 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_3306
timestamp 1745462530
transform 1 0 148 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_3307
timestamp 1745462530
transform 1 0 100 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3308
timestamp 1745462530
transform 1 0 92 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_3309
timestamp 1745462530
transform 1 0 92 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_3310
timestamp 1745462530
transform 1 0 92 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_3311
timestamp 1745462530
transform 1 0 916 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_3312
timestamp 1745462530
transform 1 0 908 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3313
timestamp 1745462530
transform 1 0 2212 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_3314
timestamp 1745462530
transform 1 0 2148 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_3315
timestamp 1745462530
transform 1 0 2124 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_3316
timestamp 1745462530
transform 1 0 2116 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_3317
timestamp 1745462530
transform 1 0 2060 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_3318
timestamp 1745462530
transform 1 0 2028 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_3319
timestamp 1745462530
transform 1 0 1988 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_3320
timestamp 1745462530
transform 1 0 1988 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_3321
timestamp 1745462530
transform 1 0 2132 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_3322
timestamp 1745462530
transform 1 0 2132 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_3323
timestamp 1745462530
transform 1 0 2052 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_3324
timestamp 1745462530
transform 1 0 1956 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_3325
timestamp 1745462530
transform 1 0 4372 0 1 4255
box -2 -2 2 2
use M2_M1  M2_M1_3326
timestamp 1745462530
transform 1 0 3932 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_3327
timestamp 1745462530
transform 1 0 3908 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_3328
timestamp 1745462530
transform 1 0 1860 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3329
timestamp 1745462530
transform 1 0 1708 0 1 4332
box -2 -2 2 2
use M2_M1  M2_M1_3330
timestamp 1745462530
transform 1 0 1620 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_3331
timestamp 1745462530
transform 1 0 1588 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_3332
timestamp 1745462530
transform 1 0 1556 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_3333
timestamp 1745462530
transform 1 0 1548 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_3334
timestamp 1745462530
transform 1 0 1548 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_3335
timestamp 1745462530
transform 1 0 1524 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_3336
timestamp 1745462530
transform 1 0 1524 0 1 2105
box -2 -2 2 2
use M2_M1  M2_M1_3337
timestamp 1745462530
transform 1 0 1396 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_3338
timestamp 1745462530
transform 1 0 1356 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_3339
timestamp 1745462530
transform 1 0 1324 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_3340
timestamp 1745462530
transform 1 0 1324 0 1 1785
box -2 -2 2 2
use M2_M1  M2_M1_3341
timestamp 1745462530
transform 1 0 1316 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_3342
timestamp 1745462530
transform 1 0 924 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_3343
timestamp 1745462530
transform 1 0 580 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_3344
timestamp 1745462530
transform 1 0 484 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_3345
timestamp 1745462530
transform 1 0 276 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_3346
timestamp 1745462530
transform 1 0 252 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_3347
timestamp 1745462530
transform 1 0 220 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_3348
timestamp 1745462530
transform 1 0 212 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_3349
timestamp 1745462530
transform 1 0 204 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_3350
timestamp 1745462530
transform 1 0 172 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_3351
timestamp 1745462530
transform 1 0 1348 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_3352
timestamp 1745462530
transform 1 0 1324 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_3353
timestamp 1745462530
transform 1 0 1316 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_3354
timestamp 1745462530
transform 1 0 1260 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_3355
timestamp 1745462530
transform 1 0 1084 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_3356
timestamp 1745462530
transform 1 0 1028 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_3357
timestamp 1745462530
transform 1 0 844 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_3358
timestamp 1745462530
transform 1 0 820 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_3359
timestamp 1745462530
transform 1 0 612 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_3360
timestamp 1745462530
transform 1 0 476 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_3361
timestamp 1745462530
transform 1 0 412 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_3362
timestamp 1745462530
transform 1 0 396 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_3363
timestamp 1745462530
transform 1 0 372 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_3364
timestamp 1745462530
transform 1 0 3172 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_3365
timestamp 1745462530
transform 1 0 3036 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_3366
timestamp 1745462530
transform 1 0 2772 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_3367
timestamp 1745462530
transform 1 0 2748 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_3368
timestamp 1745462530
transform 1 0 2740 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_3369
timestamp 1745462530
transform 1 0 2724 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_3370
timestamp 1745462530
transform 1 0 2676 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_3371
timestamp 1745462530
transform 1 0 2636 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_3372
timestamp 1745462530
transform 1 0 2612 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_3373
timestamp 1745462530
transform 1 0 2228 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_3374
timestamp 1745462530
transform 1 0 2028 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_3375
timestamp 1745462530
transform 1 0 1412 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_3376
timestamp 1745462530
transform 1 0 1412 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_3377
timestamp 1745462530
transform 1 0 4324 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_3378
timestamp 1745462530
transform 1 0 4308 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_3379
timestamp 1745462530
transform 1 0 4252 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_3380
timestamp 1745462530
transform 1 0 4228 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_3381
timestamp 1745462530
transform 1 0 4220 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_3382
timestamp 1745462530
transform 1 0 4204 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_3383
timestamp 1745462530
transform 1 0 4148 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_3384
timestamp 1745462530
transform 1 0 3780 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_3385
timestamp 1745462530
transform 1 0 3724 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_3386
timestamp 1745462530
transform 1 0 3684 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_3387
timestamp 1745462530
transform 1 0 3628 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_3388
timestamp 1745462530
transform 1 0 3612 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_3389
timestamp 1745462530
transform 1 0 3540 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_3390
timestamp 1745462530
transform 1 0 2604 0 1 1985
box -2 -2 2 2
use M2_M1  M2_M1_3391
timestamp 1745462530
transform 1 0 3700 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_3392
timestamp 1745462530
transform 1 0 3652 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_3393
timestamp 1745462530
transform 1 0 3636 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_3394
timestamp 1745462530
transform 1 0 3628 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_3395
timestamp 1745462530
transform 1 0 3620 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_3396
timestamp 1745462530
transform 1 0 3588 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_3397
timestamp 1745462530
transform 1 0 3580 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_3398
timestamp 1745462530
transform 1 0 3532 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3399
timestamp 1745462530
transform 1 0 3468 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3400
timestamp 1745462530
transform 1 0 2868 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_3401
timestamp 1745462530
transform 1 0 2852 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_3402
timestamp 1745462530
transform 1 0 2828 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_3403
timestamp 1745462530
transform 1 0 2612 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_3404
timestamp 1745462530
transform 1 0 2604 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_3405
timestamp 1745462530
transform 1 0 2572 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_3406
timestamp 1745462530
transform 1 0 1532 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_3407
timestamp 1745462530
transform 1 0 1524 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_3408
timestamp 1745462530
transform 1 0 1308 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_3409
timestamp 1745462530
transform 1 0 1292 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_3410
timestamp 1745462530
transform 1 0 2580 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_3411
timestamp 1745462530
transform 1 0 2556 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_3412
timestamp 1745462530
transform 1 0 2228 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_3413
timestamp 1745462530
transform 1 0 2212 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_3414
timestamp 1745462530
transform 1 0 1228 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_3415
timestamp 1745462530
transform 1 0 1228 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_3416
timestamp 1745462530
transform 1 0 1228 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_3417
timestamp 1745462530
transform 1 0 1180 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_3418
timestamp 1745462530
transform 1 0 1204 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_3419
timestamp 1745462530
transform 1 0 1188 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_3420
timestamp 1745462530
transform 1 0 1188 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_3421
timestamp 1745462530
transform 1 0 1164 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_3422
timestamp 1745462530
transform 1 0 1148 0 1 1835
box -2 -2 2 2
use M2_M1  M2_M1_3423
timestamp 1745462530
transform 1 0 1132 0 1 1835
box -2 -2 2 2
use M2_M1  M2_M1_3424
timestamp 1745462530
transform 1 0 1124 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_3425
timestamp 1745462530
transform 1 0 956 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3426
timestamp 1745462530
transform 1 0 836 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3427
timestamp 1745462530
transform 1 0 780 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_3428
timestamp 1745462530
transform 1 0 660 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_3429
timestamp 1745462530
transform 1 0 220 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_3430
timestamp 1745462530
transform 1 0 220 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_3431
timestamp 1745462530
transform 1 0 212 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_3432
timestamp 1745462530
transform 1 0 204 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_3433
timestamp 1745462530
transform 1 0 196 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_3434
timestamp 1745462530
transform 1 0 1420 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_3435
timestamp 1745462530
transform 1 0 1348 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_3436
timestamp 1745462530
transform 1 0 1292 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_3437
timestamp 1745462530
transform 1 0 1156 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_3438
timestamp 1745462530
transform 1 0 1132 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_3439
timestamp 1745462530
transform 1 0 1124 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_3440
timestamp 1745462530
transform 1 0 932 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_3441
timestamp 1745462530
transform 1 0 916 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_3442
timestamp 1745462530
transform 1 0 668 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_3443
timestamp 1745462530
transform 1 0 236 0 1 1255
box -2 -2 2 2
use M2_M1  M2_M1_3444
timestamp 1745462530
transform 1 0 236 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_3445
timestamp 1745462530
transform 1 0 212 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_3446
timestamp 1745462530
transform 1 0 212 0 1 1255
box -2 -2 2 2
use M2_M1  M2_M1_3447
timestamp 1745462530
transform 1 0 196 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_3448
timestamp 1745462530
transform 1 0 196 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_3449
timestamp 1745462530
transform 1 0 3308 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_3450
timestamp 1745462530
transform 1 0 2604 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_3451
timestamp 1745462530
transform 1 0 2556 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_3452
timestamp 1745462530
transform 1 0 2436 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_3453
timestamp 1745462530
transform 1 0 2396 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_3454
timestamp 1745462530
transform 1 0 2356 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_3455
timestamp 1745462530
transform 1 0 2356 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_3456
timestamp 1745462530
transform 1 0 2292 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_3457
timestamp 1745462530
transform 1 0 2292 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_3458
timestamp 1745462530
transform 1 0 2292 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_3459
timestamp 1745462530
transform 1 0 2196 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_3460
timestamp 1745462530
transform 1 0 1516 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_3461
timestamp 1745462530
transform 1 0 1452 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_3462
timestamp 1745462530
transform 1 0 1420 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_3463
timestamp 1745462530
transform 1 0 4140 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_3464
timestamp 1745462530
transform 1 0 4116 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_3465
timestamp 1745462530
transform 1 0 4092 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_3466
timestamp 1745462530
transform 1 0 4076 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_3467
timestamp 1745462530
transform 1 0 4004 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_3468
timestamp 1745462530
transform 1 0 3956 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_3469
timestamp 1745462530
transform 1 0 3668 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_3470
timestamp 1745462530
transform 1 0 3516 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_3471
timestamp 1745462530
transform 1 0 3508 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_3472
timestamp 1745462530
transform 1 0 3468 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_3473
timestamp 1745462530
transform 1 0 3452 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_3474
timestamp 1745462530
transform 1 0 3452 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_3475
timestamp 1745462530
transform 1 0 3292 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_3476
timestamp 1745462530
transform 1 0 3460 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_3477
timestamp 1745462530
transform 1 0 3428 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_3478
timestamp 1745462530
transform 1 0 3428 0 1 2395
box -2 -2 2 2
use M2_M1  M2_M1_3479
timestamp 1745462530
transform 1 0 3412 0 1 2395
box -2 -2 2 2
use M2_M1  M2_M1_3480
timestamp 1745462530
transform 1 0 3388 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_3481
timestamp 1745462530
transform 1 0 3372 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_3482
timestamp 1745462530
transform 1 0 3372 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_3483
timestamp 1745462530
transform 1 0 3276 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3484
timestamp 1745462530
transform 1 0 3212 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3485
timestamp 1745462530
transform 1 0 3196 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_3486
timestamp 1745462530
transform 1 0 2860 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_3487
timestamp 1745462530
transform 1 0 2772 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_3488
timestamp 1745462530
transform 1 0 2764 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_3489
timestamp 1745462530
transform 1 0 2732 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_3490
timestamp 1745462530
transform 1 0 2692 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_3491
timestamp 1745462530
transform 1 0 2628 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_3492
timestamp 1745462530
transform 1 0 1164 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_3493
timestamp 1745462530
transform 1 0 1164 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_3494
timestamp 1745462530
transform 1 0 1116 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_3495
timestamp 1745462530
transform 1 0 1108 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_3496
timestamp 1745462530
transform 1 0 3252 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_3497
timestamp 1745462530
transform 1 0 2836 0 1 2195
box -2 -2 2 2
use M2_M1  M2_M1_3498
timestamp 1745462530
transform 1 0 2420 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_3499
timestamp 1745462530
transform 1 0 2388 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_3500
timestamp 1745462530
transform 1 0 1876 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_3501
timestamp 1745462530
transform 1 0 1876 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_3502
timestamp 1745462530
transform 1 0 1828 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_3503
timestamp 1745462530
transform 1 0 1812 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_3504
timestamp 1745462530
transform 1 0 1836 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_3505
timestamp 1745462530
transform 1 0 1804 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_3506
timestamp 1745462530
transform 1 0 1788 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_3507
timestamp 1745462530
transform 1 0 1708 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_3508
timestamp 1745462530
transform 1 0 884 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3509
timestamp 1745462530
transform 1 0 756 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3510
timestamp 1745462530
transform 1 0 660 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3511
timestamp 1745462530
transform 1 0 660 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_3512
timestamp 1745462530
transform 1 0 444 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_3513
timestamp 1745462530
transform 1 0 356 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_3514
timestamp 1745462530
transform 1 0 340 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_3515
timestamp 1745462530
transform 1 0 332 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_3516
timestamp 1745462530
transform 1 0 324 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_3517
timestamp 1745462530
transform 1 0 1916 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_3518
timestamp 1745462530
transform 1 0 1900 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_3519
timestamp 1745462530
transform 1 0 1892 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_3520
timestamp 1745462530
transform 1 0 1884 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_3521
timestamp 1745462530
transform 1 0 1884 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_3522
timestamp 1745462530
transform 1 0 1812 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_3523
timestamp 1745462530
transform 1 0 1620 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_3524
timestamp 1745462530
transform 1 0 900 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_3525
timestamp 1745462530
transform 1 0 844 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_3526
timestamp 1745462530
transform 1 0 692 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_3527
timestamp 1745462530
transform 1 0 204 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_3528
timestamp 1745462530
transform 1 0 204 0 1 905
box -2 -2 2 2
use M2_M1  M2_M1_3529
timestamp 1745462530
transform 1 0 204 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_3530
timestamp 1745462530
transform 1 0 204 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_3531
timestamp 1745462530
transform 1 0 204 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_3532
timestamp 1745462530
transform 1 0 196 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_3533
timestamp 1745462530
transform 1 0 3364 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_3534
timestamp 1745462530
transform 1 0 2604 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_3535
timestamp 1745462530
transform 1 0 2588 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_3536
timestamp 1745462530
transform 1 0 2484 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_3537
timestamp 1745462530
transform 1 0 2452 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_3538
timestamp 1745462530
transform 1 0 2348 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_3539
timestamp 1745462530
transform 1 0 2284 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_3540
timestamp 1745462530
transform 1 0 2284 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_3541
timestamp 1745462530
transform 1 0 2284 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_3542
timestamp 1745462530
transform 1 0 2204 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_3543
timestamp 1745462530
transform 1 0 1996 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_3544
timestamp 1745462530
transform 1 0 1988 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_3545
timestamp 1745462530
transform 1 0 1980 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_3546
timestamp 1745462530
transform 1 0 4204 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_3547
timestamp 1745462530
transform 1 0 4188 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_3548
timestamp 1745462530
transform 1 0 4180 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_3549
timestamp 1745462530
transform 1 0 4148 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_3550
timestamp 1745462530
transform 1 0 4132 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_3551
timestamp 1745462530
transform 1 0 3980 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_3552
timestamp 1745462530
transform 1 0 3804 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_3553
timestamp 1745462530
transform 1 0 3788 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_3554
timestamp 1745462530
transform 1 0 3780 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_3555
timestamp 1745462530
transform 1 0 3780 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_3556
timestamp 1745462530
transform 1 0 3780 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_3557
timestamp 1745462530
transform 1 0 3756 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_3558
timestamp 1745462530
transform 1 0 3740 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_3559
timestamp 1745462530
transform 1 0 2764 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_3560
timestamp 1745462530
transform 1 0 3948 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_3561
timestamp 1745462530
transform 1 0 3948 0 1 1895
box -2 -2 2 2
use M2_M1  M2_M1_3562
timestamp 1745462530
transform 1 0 3932 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_3563
timestamp 1745462530
transform 1 0 3876 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_3564
timestamp 1745462530
transform 1 0 3868 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_3565
timestamp 1745462530
transform 1 0 3852 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_3566
timestamp 1745462530
transform 1 0 3844 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_3567
timestamp 1745462530
transform 1 0 3844 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_3568
timestamp 1745462530
transform 1 0 3836 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_3569
timestamp 1745462530
transform 1 0 3764 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_3570
timestamp 1745462530
transform 1 0 3732 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3571
timestamp 1745462530
transform 1 0 2972 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_3572
timestamp 1745462530
transform 1 0 2972 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_3573
timestamp 1745462530
transform 1 0 2940 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_3574
timestamp 1745462530
transform 1 0 2940 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_3575
timestamp 1745462530
transform 1 0 2924 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_3576
timestamp 1745462530
transform 1 0 2716 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_3577
timestamp 1745462530
transform 1 0 2700 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_3578
timestamp 1745462530
transform 1 0 2500 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_3579
timestamp 1745462530
transform 1 0 1860 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_3580
timestamp 1745462530
transform 1 0 1860 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_3581
timestamp 1745462530
transform 1 0 1788 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_3582
timestamp 1745462530
transform 1 0 1788 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_3583
timestamp 1745462530
transform 1 0 2732 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_3584
timestamp 1745462530
transform 1 0 2700 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_3585
timestamp 1745462530
transform 1 0 2188 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_3586
timestamp 1745462530
transform 1 0 2156 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_3587
timestamp 1745462530
transform 1 0 1740 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_3588
timestamp 1745462530
transform 1 0 1700 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_3589
timestamp 1745462530
transform 1 0 1700 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_3590
timestamp 1745462530
transform 1 0 1684 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_3591
timestamp 1745462530
transform 1 0 1724 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_3592
timestamp 1745462530
transform 1 0 1564 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_3593
timestamp 1745462530
transform 1 0 1564 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_3594
timestamp 1745462530
transform 1 0 1532 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_3595
timestamp 1745462530
transform 1 0 1532 0 1 2185
box -2 -2 2 2
use M2_M1  M2_M1_3596
timestamp 1745462530
transform 1 0 1516 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_3597
timestamp 1745462530
transform 1 0 956 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_3598
timestamp 1745462530
transform 1 0 556 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_3599
timestamp 1745462530
transform 1 0 532 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_3600
timestamp 1745462530
transform 1 0 492 0 1 2595
box -2 -2 2 2
use M2_M1  M2_M1_3601
timestamp 1745462530
transform 1 0 452 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_3602
timestamp 1745462530
transform 1 0 428 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_3603
timestamp 1745462530
transform 1 0 420 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_3604
timestamp 1745462530
transform 1 0 420 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_3605
timestamp 1745462530
transform 1 0 348 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_3606
timestamp 1745462530
transform 1 0 340 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_3607
timestamp 1745462530
transform 1 0 1876 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_3608
timestamp 1745462530
transform 1 0 1836 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_3609
timestamp 1745462530
transform 1 0 1828 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_3610
timestamp 1745462530
transform 1 0 1820 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_3611
timestamp 1745462530
transform 1 0 1780 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_3612
timestamp 1745462530
transform 1 0 1692 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_3613
timestamp 1745462530
transform 1 0 1684 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_3614
timestamp 1745462530
transform 1 0 812 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_3615
timestamp 1745462530
transform 1 0 740 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_3616
timestamp 1745462530
transform 1 0 540 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_3617
timestamp 1745462530
transform 1 0 372 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_3618
timestamp 1745462530
transform 1 0 316 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_3619
timestamp 1745462530
transform 1 0 308 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_3620
timestamp 1745462530
transform 1 0 292 0 1 435
box -2 -2 2 2
use M2_M1  M2_M1_3621
timestamp 1745462530
transform 1 0 284 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_3622
timestamp 1745462530
transform 1 0 252 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_3623
timestamp 1745462530
transform 1 0 3404 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_3624
timestamp 1745462530
transform 1 0 2500 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_3625
timestamp 1745462530
transform 1 0 2364 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_3626
timestamp 1745462530
transform 1 0 2348 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_3627
timestamp 1745462530
transform 1 0 2348 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_3628
timestamp 1745462530
transform 1 0 2292 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_3629
timestamp 1745462530
transform 1 0 2236 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_3630
timestamp 1745462530
transform 1 0 2236 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_3631
timestamp 1745462530
transform 1 0 2228 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_3632
timestamp 1745462530
transform 1 0 2196 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_3633
timestamp 1745462530
transform 1 0 2020 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_3634
timestamp 1745462530
transform 1 0 1996 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_3635
timestamp 1745462530
transform 1 0 1924 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_3636
timestamp 1745462530
transform 1 0 4308 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_3637
timestamp 1745462530
transform 1 0 4308 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_3638
timestamp 1745462530
transform 1 0 4220 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_3639
timestamp 1745462530
transform 1 0 4220 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_3640
timestamp 1745462530
transform 1 0 4220 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_3641
timestamp 1745462530
transform 1 0 4212 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_3642
timestamp 1745462530
transform 1 0 4180 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_3643
timestamp 1745462530
transform 1 0 3964 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_3644
timestamp 1745462530
transform 1 0 3916 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_3645
timestamp 1745462530
transform 1 0 3812 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_3646
timestamp 1745462530
transform 1 0 3668 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_3647
timestamp 1745462530
transform 1 0 3636 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_3648
timestamp 1745462530
transform 1 0 2724 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_3649
timestamp 1745462530
transform 1 0 4220 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3650
timestamp 1745462530
transform 1 0 4220 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_3651
timestamp 1745462530
transform 1 0 4196 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_3652
timestamp 1745462530
transform 1 0 4180 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_3653
timestamp 1745462530
transform 1 0 4140 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_3654
timestamp 1745462530
transform 1 0 4052 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3655
timestamp 1745462530
transform 1 0 3900 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3656
timestamp 1745462530
transform 1 0 3244 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_3657
timestamp 1745462530
transform 1 0 2868 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_3658
timestamp 1745462530
transform 1 0 2836 0 1 2505
box -2 -2 2 2
use M2_M1  M2_M1_3659
timestamp 1745462530
transform 1 0 2836 0 1 2485
box -2 -2 2 2
use M2_M1  M2_M1_3660
timestamp 1745462530
transform 1 0 2828 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_3661
timestamp 1745462530
transform 1 0 2740 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_3662
timestamp 1745462530
transform 1 0 2668 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_3663
timestamp 1745462530
transform 1 0 2612 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_3664
timestamp 1745462530
transform 1 0 1708 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_3665
timestamp 1745462530
transform 1 0 1708 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_3666
timestamp 1745462530
transform 1 0 1684 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_3667
timestamp 1745462530
transform 1 0 1676 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_3668
timestamp 1745462530
transform 1 0 1676 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_3669
timestamp 1745462530
transform 1 0 2724 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_3670
timestamp 1745462530
transform 1 0 2692 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_3671
timestamp 1745462530
transform 1 0 2292 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_3672
timestamp 1745462530
transform 1 0 2188 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_3673
timestamp 1745462530
transform 1 0 1316 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_3674
timestamp 1745462530
transform 1 0 1308 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_3675
timestamp 1745462530
transform 1 0 1292 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_3676
timestamp 1745462530
transform 1 0 1284 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_3677
timestamp 1745462530
transform 1 0 1284 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_3678
timestamp 1745462530
transform 1 0 1276 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_3679
timestamp 1745462530
transform 1 0 1236 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_3680
timestamp 1745462530
transform 1 0 1228 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_3681
timestamp 1745462530
transform 1 0 1228 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_3682
timestamp 1745462530
transform 1 0 1220 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_3683
timestamp 1745462530
transform 1 0 1204 0 1 1885
box -2 -2 2 2
use M2_M1  M2_M1_3684
timestamp 1745462530
transform 1 0 956 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_3685
timestamp 1745462530
transform 1 0 684 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_3686
timestamp 1745462530
transform 1 0 532 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_3687
timestamp 1745462530
transform 1 0 476 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_3688
timestamp 1745462530
transform 1 0 420 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_3689
timestamp 1745462530
transform 1 0 420 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_3690
timestamp 1745462530
transform 1 0 404 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_3691
timestamp 1745462530
transform 1 0 388 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_3692
timestamp 1745462530
transform 1 0 372 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_3693
timestamp 1745462530
transform 1 0 292 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_3694
timestamp 1745462530
transform 1 0 1476 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_3695
timestamp 1745462530
transform 1 0 1452 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_3696
timestamp 1745462530
transform 1 0 1396 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_3697
timestamp 1745462530
transform 1 0 1388 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_3698
timestamp 1745462530
transform 1 0 1292 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_3699
timestamp 1745462530
transform 1 0 1140 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_3700
timestamp 1745462530
transform 1 0 900 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_3701
timestamp 1745462530
transform 1 0 700 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_3702
timestamp 1745462530
transform 1 0 636 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_3703
timestamp 1745462530
transform 1 0 404 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_3704
timestamp 1745462530
transform 1 0 380 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_3705
timestamp 1745462530
transform 1 0 380 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_3706
timestamp 1745462530
transform 1 0 324 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_3707
timestamp 1745462530
transform 1 0 3252 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_3708
timestamp 1745462530
transform 1 0 3076 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_3709
timestamp 1745462530
transform 1 0 2980 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_3710
timestamp 1745462530
transform 1 0 2964 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_3711
timestamp 1745462530
transform 1 0 2900 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_3712
timestamp 1745462530
transform 1 0 2884 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_3713
timestamp 1745462530
transform 1 0 2844 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_3714
timestamp 1745462530
transform 1 0 2836 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_3715
timestamp 1745462530
transform 1 0 2836 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_3716
timestamp 1745462530
transform 1 0 2820 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_3717
timestamp 1745462530
transform 1 0 2636 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_3718
timestamp 1745462530
transform 1 0 2596 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_3719
timestamp 1745462530
transform 1 0 1660 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_3720
timestamp 1745462530
transform 1 0 1636 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_3721
timestamp 1745462530
transform 1 0 1596 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_3722
timestamp 1745462530
transform 1 0 1588 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_3723
timestamp 1745462530
transform 1 0 4164 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_3724
timestamp 1745462530
transform 1 0 4124 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_3725
timestamp 1745462530
transform 1 0 4076 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_3726
timestamp 1745462530
transform 1 0 4068 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_3727
timestamp 1745462530
transform 1 0 4068 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_3728
timestamp 1745462530
transform 1 0 4060 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_3729
timestamp 1745462530
transform 1 0 4060 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_3730
timestamp 1745462530
transform 1 0 3548 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_3731
timestamp 1745462530
transform 1 0 3484 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_3732
timestamp 1745462530
transform 1 0 3372 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_3733
timestamp 1745462530
transform 1 0 3364 0 1 1035
box -2 -2 2 2
use M2_M1  M2_M1_3734
timestamp 1745462530
transform 1 0 3356 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_3735
timestamp 1745462530
transform 1 0 3356 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_3736
timestamp 1745462530
transform 1 0 2908 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_3737
timestamp 1745462530
transform 1 0 3284 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_3738
timestamp 1745462530
transform 1 0 3276 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_3739
timestamp 1745462530
transform 1 0 3252 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_3740
timestamp 1745462530
transform 1 0 3252 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_3741
timestamp 1745462530
transform 1 0 3236 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_3742
timestamp 1745462530
transform 1 0 3228 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_3743
timestamp 1745462530
transform 1 0 3204 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_3744
timestamp 1745462530
transform 1 0 3180 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3745
timestamp 1745462530
transform 1 0 3004 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3746
timestamp 1745462530
transform 1 0 2884 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_3747
timestamp 1745462530
transform 1 0 2796 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_3748
timestamp 1745462530
transform 1 0 2772 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_3749
timestamp 1745462530
transform 1 0 2772 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_3750
timestamp 1745462530
transform 1 0 2756 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_3751
timestamp 1745462530
transform 1 0 1644 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_3752
timestamp 1745462530
transform 1 0 1284 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_3753
timestamp 1745462530
transform 1 0 1276 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_3754
timestamp 1745462530
transform 1 0 1220 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_3755
timestamp 1745462530
transform 1 0 2892 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_3756
timestamp 1745462530
transform 1 0 2868 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_3757
timestamp 1745462530
transform 1 0 2844 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_3758
timestamp 1745462530
transform 1 0 2588 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_3759
timestamp 1745462530
transform 1 0 2580 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_3760
timestamp 1745462530
transform 1 0 1948 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_3761
timestamp 1745462530
transform 1 0 1892 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_3762
timestamp 1745462530
transform 1 0 1884 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_3763
timestamp 1745462530
transform 1 0 1884 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_3764
timestamp 1745462530
transform 1 0 1788 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_3765
timestamp 1745462530
transform 1 0 1788 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_3766
timestamp 1745462530
transform 1 0 1780 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_3767
timestamp 1745462530
transform 1 0 1724 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_3768
timestamp 1745462530
transform 1 0 964 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_3769
timestamp 1745462530
transform 1 0 588 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_3770
timestamp 1745462530
transform 1 0 580 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_3771
timestamp 1745462530
transform 1 0 372 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_3772
timestamp 1745462530
transform 1 0 332 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_3773
timestamp 1745462530
transform 1 0 276 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_3774
timestamp 1745462530
transform 1 0 260 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_3775
timestamp 1745462530
transform 1 0 260 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_3776
timestamp 1745462530
transform 1 0 212 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_3777
timestamp 1745462530
transform 1 0 1780 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_3778
timestamp 1745462530
transform 1 0 1732 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_3779
timestamp 1745462530
transform 1 0 1724 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_3780
timestamp 1745462530
transform 1 0 1660 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_3781
timestamp 1745462530
transform 1 0 1660 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_3782
timestamp 1745462530
transform 1 0 1492 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_3783
timestamp 1745462530
transform 1 0 844 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_3784
timestamp 1745462530
transform 1 0 708 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_3785
timestamp 1745462530
transform 1 0 684 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_3786
timestamp 1745462530
transform 1 0 484 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_3787
timestamp 1745462530
transform 1 0 468 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_3788
timestamp 1745462530
transform 1 0 436 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_3789
timestamp 1745462530
transform 1 0 244 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_3790
timestamp 1745462530
transform 1 0 244 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_3791
timestamp 1745462530
transform 1 0 3308 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_3792
timestamp 1745462530
transform 1 0 3076 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_3793
timestamp 1745462530
transform 1 0 3028 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_3794
timestamp 1745462530
transform 1 0 2908 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_3795
timestamp 1745462530
transform 1 0 2908 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_3796
timestamp 1745462530
transform 1 0 2900 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_3797
timestamp 1745462530
transform 1 0 2836 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_3798
timestamp 1745462530
transform 1 0 2812 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_3799
timestamp 1745462530
transform 1 0 2796 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_3800
timestamp 1745462530
transform 1 0 2572 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_3801
timestamp 1745462530
transform 1 0 1836 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_3802
timestamp 1745462530
transform 1 0 1836 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_3803
timestamp 1745462530
transform 1 0 1788 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_3804
timestamp 1745462530
transform 1 0 4308 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_3805
timestamp 1745462530
transform 1 0 4220 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_3806
timestamp 1745462530
transform 1 0 4180 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_3807
timestamp 1745462530
transform 1 0 4156 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_3808
timestamp 1745462530
transform 1 0 4148 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_3809
timestamp 1745462530
transform 1 0 4132 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_3810
timestamp 1745462530
transform 1 0 4124 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_3811
timestamp 1745462530
transform 1 0 4108 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_3812
timestamp 1745462530
transform 1 0 3956 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_3813
timestamp 1745462530
transform 1 0 3884 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_3814
timestamp 1745462530
transform 1 0 3876 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_3815
timestamp 1745462530
transform 1 0 3820 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_3816
timestamp 1745462530
transform 1 0 3820 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_3817
timestamp 1745462530
transform 1 0 3804 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_3818
timestamp 1745462530
transform 1 0 4212 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_3819
timestamp 1745462530
transform 1 0 4212 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_3820
timestamp 1745462530
transform 1 0 4188 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_3821
timestamp 1745462530
transform 1 0 4148 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_3822
timestamp 1745462530
transform 1 0 4084 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_3823
timestamp 1745462530
transform 1 0 4084 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_3824
timestamp 1745462530
transform 1 0 3908 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_3825
timestamp 1745462530
transform 1 0 3852 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_3826
timestamp 1745462530
transform 1 0 3100 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_3827
timestamp 1745462530
transform 1 0 2924 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_3828
timestamp 1745462530
transform 1 0 2876 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_3829
timestamp 1745462530
transform 1 0 2772 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_3830
timestamp 1745462530
transform 1 0 1868 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_3831
timestamp 1745462530
transform 1 0 1852 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_3832
timestamp 1745462530
transform 1 0 1772 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_3833
timestamp 1745462530
transform 1 0 1764 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_3834
timestamp 1745462530
transform 1 0 3804 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_3835
timestamp 1745462530
transform 1 0 3780 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_3836
timestamp 1745462530
transform 1 0 2556 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_3837
timestamp 1745462530
transform 1 0 2468 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_3838
timestamp 1745462530
transform 1 0 3828 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_3839
timestamp 1745462530
transform 1 0 3828 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_3840
timestamp 1745462530
transform 1 0 3732 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_3841
timestamp 1745462530
transform 1 0 3716 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_3842
timestamp 1745462530
transform 1 0 3572 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_3843
timestamp 1745462530
transform 1 0 2428 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_3844
timestamp 1745462530
transform 1 0 2412 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_3845
timestamp 1745462530
transform 1 0 2116 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_3846
timestamp 1745462530
transform 1 0 1940 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_3847
timestamp 1745462530
transform 1 0 1140 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_3848
timestamp 1745462530
transform 1 0 1028 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_3849
timestamp 1745462530
transform 1 0 1004 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_3850
timestamp 1745462530
transform 1 0 956 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_3851
timestamp 1745462530
transform 1 0 3388 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_3852
timestamp 1745462530
transform 1 0 3388 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_3853
timestamp 1745462530
transform 1 0 3324 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_3854
timestamp 1745462530
transform 1 0 3324 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_3855
timestamp 1745462530
transform 1 0 2812 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_3856
timestamp 1745462530
transform 1 0 2452 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_3857
timestamp 1745462530
transform 1 0 2428 0 1 1255
box -2 -2 2 2
use M2_M1  M2_M1_3858
timestamp 1745462530
transform 1 0 2428 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_3859
timestamp 1745462530
transform 1 0 2412 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_3860
timestamp 1745462530
transform 1 0 1476 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_3861
timestamp 1745462530
transform 1 0 1212 0 1 1995
box -2 -2 2 2
use M2_M1  M2_M1_3862
timestamp 1745462530
transform 1 0 1212 0 1 1955
box -2 -2 2 2
use M2_M1  M2_M1_3863
timestamp 1745462530
transform 1 0 1204 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_3864
timestamp 1745462530
transform 1 0 1204 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_3865
timestamp 1745462530
transform 1 0 1180 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_3866
timestamp 1745462530
transform 1 0 1108 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_3867
timestamp 1745462530
transform 1 0 1044 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_3868
timestamp 1745462530
transform 1 0 1036 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_3869
timestamp 1745462530
transform 1 0 972 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_3870
timestamp 1745462530
transform 1 0 4124 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_3871
timestamp 1745462530
transform 1 0 4116 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_3872
timestamp 1745462530
transform 1 0 4068 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_3873
timestamp 1745462530
transform 1 0 4004 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_3874
timestamp 1745462530
transform 1 0 3964 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_3875
timestamp 1745462530
transform 1 0 3060 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_3876
timestamp 1745462530
transform 1 0 2404 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_3877
timestamp 1745462530
transform 1 0 2060 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_3878
timestamp 1745462530
transform 1 0 1868 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_3879
timestamp 1745462530
transform 1 0 1724 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_3880
timestamp 1745462530
transform 1 0 932 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_3881
timestamp 1745462530
transform 1 0 908 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_3882
timestamp 1745462530
transform 1 0 892 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_3883
timestamp 1745462530
transform 1 0 3228 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_3884
timestamp 1745462530
transform 1 0 3220 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_3885
timestamp 1745462530
transform 1 0 3212 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_3886
timestamp 1745462530
transform 1 0 3140 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_3887
timestamp 1745462530
transform 1 0 3124 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_3888
timestamp 1745462530
transform 1 0 2436 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_3889
timestamp 1745462530
transform 1 0 2348 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_3890
timestamp 1745462530
transform 1 0 1660 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_3891
timestamp 1745462530
transform 1 0 1428 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_3892
timestamp 1745462530
transform 1 0 1332 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_3893
timestamp 1745462530
transform 1 0 1068 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_3894
timestamp 1745462530
transform 1 0 1068 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_3895
timestamp 1745462530
transform 1 0 1004 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_3896
timestamp 1745462530
transform 1 0 3812 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_3897
timestamp 1745462530
transform 1 0 3796 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_3898
timestamp 1745462530
transform 1 0 3700 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_3899
timestamp 1745462530
transform 1 0 3692 0 1 1595
box -2 -2 2 2
use M2_M1  M2_M1_3900
timestamp 1745462530
transform 1 0 3684 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_3901
timestamp 1745462530
transform 1 0 3580 0 1 2155
box -2 -2 2 2
use M2_M1  M2_M1_3902
timestamp 1745462530
transform 1 0 3572 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_3903
timestamp 1745462530
transform 1 0 3556 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_3904
timestamp 1745462530
transform 1 0 2380 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_3905
timestamp 1745462530
transform 1 0 2364 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_3906
timestamp 1745462530
transform 1 0 2348 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_3907
timestamp 1745462530
transform 1 0 2092 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_3908
timestamp 1745462530
transform 1 0 1924 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_3909
timestamp 1745462530
transform 1 0 1124 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_3910
timestamp 1745462530
transform 1 0 1012 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_3911
timestamp 1745462530
transform 1 0 980 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_3912
timestamp 1745462530
transform 1 0 940 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_3913
timestamp 1745462530
transform 1 0 3372 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_3914
timestamp 1745462530
transform 1 0 3356 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_3915
timestamp 1745462530
transform 1 0 3300 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_3916
timestamp 1745462530
transform 1 0 3292 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_3917
timestamp 1745462530
transform 1 0 2788 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_3918
timestamp 1745462530
transform 1 0 2436 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_3919
timestamp 1745462530
transform 1 0 2372 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_3920
timestamp 1745462530
transform 1 0 1460 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_3921
timestamp 1745462530
transform 1 0 1164 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_3922
timestamp 1745462530
transform 1 0 1092 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_3923
timestamp 1745462530
transform 1 0 1020 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_3924
timestamp 1745462530
transform 1 0 1012 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_3925
timestamp 1745462530
transform 1 0 924 0 1 905
box -2 -2 2 2
use M2_M1  M2_M1_3926
timestamp 1745462530
transform 1 0 4100 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_3927
timestamp 1745462530
transform 1 0 4100 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_3928
timestamp 1745462530
transform 1 0 4028 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_3929
timestamp 1745462530
transform 1 0 3988 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_3930
timestamp 1745462530
transform 1 0 3948 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_3931
timestamp 1745462530
transform 1 0 3036 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_3932
timestamp 1745462530
transform 1 0 2340 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_3933
timestamp 1745462530
transform 1 0 2028 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_3934
timestamp 1745462530
transform 1 0 1828 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_3935
timestamp 1745462530
transform 1 0 1684 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_3936
timestamp 1745462530
transform 1 0 892 0 1 2185
box -2 -2 2 2
use M2_M1  M2_M1_3937
timestamp 1745462530
transform 1 0 892 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_3938
timestamp 1745462530
transform 1 0 876 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_3939
timestamp 1745462530
transform 1 0 876 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_3940
timestamp 1745462530
transform 1 0 3212 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_3941
timestamp 1745462530
transform 1 0 3172 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_3942
timestamp 1745462530
transform 1 0 3156 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_3943
timestamp 1745462530
transform 1 0 3124 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_3944
timestamp 1745462530
transform 1 0 3108 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_3945
timestamp 1745462530
transform 1 0 2332 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_3946
timestamp 1745462530
transform 1 0 2324 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_3947
timestamp 1745462530
transform 1 0 1644 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_3948
timestamp 1745462530
transform 1 0 1412 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_3949
timestamp 1745462530
transform 1 0 1404 0 1 685
box -2 -2 2 2
use M2_M1  M2_M1_3950
timestamp 1745462530
transform 1 0 1380 0 1 685
box -2 -2 2 2
use M2_M1  M2_M1_3951
timestamp 1745462530
transform 1 0 1316 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_3952
timestamp 1745462530
transform 1 0 1052 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_3953
timestamp 1745462530
transform 1 0 1020 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_3954
timestamp 1745462530
transform 1 0 988 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_3955
timestamp 1745462530
transform 1 0 3660 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_3956
timestamp 1745462530
transform 1 0 3548 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_3957
timestamp 1745462530
transform 1 0 3076 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_3958
timestamp 1745462530
transform 1 0 3052 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_3959
timestamp 1745462530
transform 1 0 3036 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_3960
timestamp 1745462530
transform 1 0 2636 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_3961
timestamp 1745462530
transform 1 0 2524 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_3962
timestamp 1745462530
transform 1 0 2516 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_3963
timestamp 1745462530
transform 1 0 2092 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_3964
timestamp 1745462530
transform 1 0 1932 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_3965
timestamp 1745462530
transform 1 0 1220 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_3966
timestamp 1745462530
transform 1 0 1028 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_3967
timestamp 1745462530
transform 1 0 924 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_3968
timestamp 1745462530
transform 1 0 876 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_3969
timestamp 1745462530
transform 1 0 3308 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_3970
timestamp 1745462530
transform 1 0 2876 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_3971
timestamp 1745462530
transform 1 0 2732 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_3972
timestamp 1745462530
transform 1 0 2716 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_3973
timestamp 1745462530
transform 1 0 2516 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_3974
timestamp 1745462530
transform 1 0 2476 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_3975
timestamp 1745462530
transform 1 0 2460 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_3976
timestamp 1745462530
transform 1 0 1332 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_3977
timestamp 1745462530
transform 1 0 1316 0 1 1595
box -2 -2 2 2
use M2_M1  M2_M1_3978
timestamp 1745462530
transform 1 0 1260 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_3979
timestamp 1745462530
transform 1 0 1164 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_3980
timestamp 1745462530
transform 1 0 1164 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_3981
timestamp 1745462530
transform 1 0 1116 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_3982
timestamp 1745462530
transform 1 0 996 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_3983
timestamp 1745462530
transform 1 0 3892 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_3984
timestamp 1745462530
transform 1 0 3860 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_3985
timestamp 1745462530
transform 1 0 3108 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_3986
timestamp 1745462530
transform 1 0 3084 0 1 1755
box -2 -2 2 2
use M2_M1  M2_M1_3987
timestamp 1745462530
transform 1 0 3084 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_3988
timestamp 1745462530
transform 1 0 3068 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_3989
timestamp 1745462530
transform 1 0 3044 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_3990
timestamp 1745462530
transform 1 0 2980 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_3991
timestamp 1745462530
transform 1 0 2948 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_3992
timestamp 1745462530
transform 1 0 2932 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_3993
timestamp 1745462530
transform 1 0 2484 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_3994
timestamp 1745462530
transform 1 0 2012 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_3995
timestamp 1745462530
transform 1 0 1940 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_3996
timestamp 1745462530
transform 1 0 1916 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_3997
timestamp 1745462530
transform 1 0 1900 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_3998
timestamp 1745462530
transform 1 0 1692 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_3999
timestamp 1745462530
transform 1 0 988 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_4000
timestamp 1745462530
transform 1 0 932 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_4001
timestamp 1745462530
transform 1 0 924 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_4002
timestamp 1745462530
transform 1 0 3092 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_4003
timestamp 1745462530
transform 1 0 2980 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_4004
timestamp 1745462530
transform 1 0 2876 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_4005
timestamp 1745462530
transform 1 0 2732 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_4006
timestamp 1745462530
transform 1 0 2612 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_4007
timestamp 1745462530
transform 1 0 2508 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_4008
timestamp 1745462530
transform 1 0 2332 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_4009
timestamp 1745462530
transform 1 0 1516 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_4010
timestamp 1745462530
transform 1 0 1516 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_4011
timestamp 1745462530
transform 1 0 1492 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_4012
timestamp 1745462530
transform 1 0 1252 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_4013
timestamp 1745462530
transform 1 0 1028 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_4014
timestamp 1745462530
transform 1 0 996 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_4015
timestamp 1745462530
transform 1 0 956 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_4016
timestamp 1745462530
transform 1 0 3796 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_4017
timestamp 1745462530
transform 1 0 3772 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_4018
timestamp 1745462530
transform 1 0 3708 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_4019
timestamp 1745462530
transform 1 0 3652 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_4020
timestamp 1745462530
transform 1 0 3612 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_4021
timestamp 1745462530
transform 1 0 2564 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_4022
timestamp 1745462530
transform 1 0 2556 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_4023
timestamp 1745462530
transform 1 0 2036 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_4024
timestamp 1745462530
transform 1 0 1852 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_4025
timestamp 1745462530
transform 1 0 1092 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_4026
timestamp 1745462530
transform 1 0 820 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_4027
timestamp 1745462530
transform 1 0 804 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_4028
timestamp 1745462530
transform 1 0 780 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_4029
timestamp 1745462530
transform 1 0 3612 0 1 1995
box -2 -2 2 2
use M2_M1  M2_M1_4030
timestamp 1745462530
transform 1 0 3612 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_4031
timestamp 1745462530
transform 1 0 3612 0 1 1555
box -2 -2 2 2
use M2_M1  M2_M1_4032
timestamp 1745462530
transform 1 0 3604 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_4033
timestamp 1745462530
transform 1 0 3580 0 1 1555
box -2 -2 2 2
use M2_M1  M2_M1_4034
timestamp 1745462530
transform 1 0 3548 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_4035
timestamp 1745462530
transform 1 0 3460 0 1 635
box -2 -2 2 2
use M2_M1  M2_M1_4036
timestamp 1745462530
transform 1 0 2732 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_4037
timestamp 1745462530
transform 1 0 2588 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_4038
timestamp 1745462530
transform 1 0 2436 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_4039
timestamp 1745462530
transform 1 0 2404 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_4040
timestamp 1745462530
transform 1 0 1548 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_4041
timestamp 1745462530
transform 1 0 1212 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_4042
timestamp 1745462530
transform 1 0 1172 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_4043
timestamp 1745462530
transform 1 0 876 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_4044
timestamp 1745462530
transform 1 0 644 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_4045
timestamp 1745462530
transform 1 0 580 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_4046
timestamp 1745462530
transform 1 0 4148 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4047
timestamp 1745462530
transform 1 0 4140 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_4048
timestamp 1745462530
transform 1 0 4076 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_4049
timestamp 1745462530
transform 1 0 3940 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_4050
timestamp 1745462530
transform 1 0 3876 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_4051
timestamp 1745462530
transform 1 0 2988 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_4052
timestamp 1745462530
transform 1 0 2652 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_4053
timestamp 1745462530
transform 1 0 1996 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4054
timestamp 1745462530
transform 1 0 1772 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_4055
timestamp 1745462530
transform 1 0 1652 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_4056
timestamp 1745462530
transform 1 0 652 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4057
timestamp 1745462530
transform 1 0 612 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4058
timestamp 1745462530
transform 1 0 604 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_4059
timestamp 1745462530
transform 1 0 3460 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_4060
timestamp 1745462530
transform 1 0 3444 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_4061
timestamp 1745462530
transform 1 0 3444 0 1 1435
box -2 -2 2 2
use M2_M1  M2_M1_4062
timestamp 1745462530
transform 1 0 3364 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_4063
timestamp 1745462530
transform 1 0 3244 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4064
timestamp 1745462530
transform 1 0 3236 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_4065
timestamp 1745462530
transform 1 0 2924 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_4066
timestamp 1745462530
transform 1 0 2628 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_4067
timestamp 1745462530
transform 1 0 2252 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_4068
timestamp 1745462530
transform 1 0 1692 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_4069
timestamp 1745462530
transform 1 0 1396 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_4070
timestamp 1745462530
transform 1 0 1372 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_4071
timestamp 1745462530
transform 1 0 612 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_4072
timestamp 1745462530
transform 1 0 612 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_4073
timestamp 1745462530
transform 1 0 540 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_4074
timestamp 1745462530
transform 1 0 3796 0 1 2635
box -2 -2 2 2
use M2_M1  M2_M1_4075
timestamp 1745462530
transform 1 0 3780 0 1 2595
box -2 -2 2 2
use M2_M1  M2_M1_4076
timestamp 1745462530
transform 1 0 3756 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_4077
timestamp 1745462530
transform 1 0 3756 0 1 1505
box -2 -2 2 2
use M2_M1  M2_M1_4078
timestamp 1745462530
transform 1 0 3740 0 1 1505
box -2 -2 2 2
use M2_M1  M2_M1_4079
timestamp 1745462530
transform 1 0 3740 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_4080
timestamp 1745462530
transform 1 0 3676 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_4081
timestamp 1745462530
transform 1 0 2516 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_4082
timestamp 1745462530
transform 1 0 2500 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_4083
timestamp 1745462530
transform 1 0 1988 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_4084
timestamp 1745462530
transform 1 0 1820 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_4085
timestamp 1745462530
transform 1 0 1060 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_4086
timestamp 1745462530
transform 1 0 788 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_4087
timestamp 1745462530
transform 1 0 772 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_4088
timestamp 1745462530
transform 1 0 3620 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_4089
timestamp 1745462530
transform 1 0 3580 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_4090
timestamp 1745462530
transform 1 0 3580 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_4091
timestamp 1745462530
transform 1 0 3548 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_4092
timestamp 1745462530
transform 1 0 3516 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_4093
timestamp 1745462530
transform 1 0 3420 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_4094
timestamp 1745462530
transform 1 0 2700 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_4095
timestamp 1745462530
transform 1 0 2476 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_4096
timestamp 1745462530
transform 1 0 1500 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_4097
timestamp 1745462530
transform 1 0 1180 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_4098
timestamp 1745462530
transform 1 0 1116 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_4099
timestamp 1745462530
transform 1 0 836 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_4100
timestamp 1745462530
transform 1 0 748 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_4101
timestamp 1745462530
transform 1 0 612 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_4102
timestamp 1745462530
transform 1 0 548 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_4103
timestamp 1745462530
transform 1 0 4108 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_4104
timestamp 1745462530
transform 1 0 4100 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_4105
timestamp 1745462530
transform 1 0 4020 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_4106
timestamp 1745462530
transform 1 0 3908 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_4107
timestamp 1745462530
transform 1 0 3572 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_4108
timestamp 1745462530
transform 1 0 2956 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_4109
timestamp 1745462530
transform 1 0 2532 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_4110
timestamp 1745462530
transform 1 0 2356 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_4111
timestamp 1745462530
transform 1 0 1948 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4112
timestamp 1745462530
transform 1 0 1740 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_4113
timestamp 1745462530
transform 1 0 1620 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_4114
timestamp 1745462530
transform 1 0 1596 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_4115
timestamp 1745462530
transform 1 0 620 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4116
timestamp 1745462530
transform 1 0 580 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4117
timestamp 1745462530
transform 1 0 572 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_4118
timestamp 1745462530
transform 1 0 3844 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_4119
timestamp 1745462530
transform 1 0 3380 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_4120
timestamp 1745462530
transform 1 0 3348 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_4121
timestamp 1745462530
transform 1 0 3332 0 1 1435
box -2 -2 2 2
use M2_M1  M2_M1_4122
timestamp 1745462530
transform 1 0 3300 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_4123
timestamp 1745462530
transform 1 0 3212 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4124
timestamp 1745462530
transform 1 0 3204 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_4125
timestamp 1745462530
transform 1 0 2876 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_4126
timestamp 1745462530
transform 1 0 2452 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_4127
timestamp 1745462530
transform 1 0 2220 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_4128
timestamp 1745462530
transform 1 0 1660 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_4129
timestamp 1745462530
transform 1 0 1364 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_4130
timestamp 1745462530
transform 1 0 1332 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_4131
timestamp 1745462530
transform 1 0 572 0 1 2845
box -2 -2 2 2
use M2_M1  M2_M1_4132
timestamp 1745462530
transform 1 0 572 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_4133
timestamp 1745462530
transform 1 0 508 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_4134
timestamp 1745462530
transform 1 0 3748 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4135
timestamp 1745462530
transform 1 0 3740 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_4136
timestamp 1745462530
transform 1 0 3716 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_4137
timestamp 1745462530
transform 1 0 3620 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4138
timestamp 1745462530
transform 1 0 3620 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_4139
timestamp 1745462530
transform 1 0 2540 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_4140
timestamp 1745462530
transform 1 0 2500 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_4141
timestamp 1745462530
transform 1 0 2036 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_4142
timestamp 1745462530
transform 1 0 1852 0 1 2505
box -2 -2 2 2
use M2_M1  M2_M1_4143
timestamp 1745462530
transform 1 0 1068 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_4144
timestamp 1745462530
transform 1 0 812 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_4145
timestamp 1745462530
transform 1 0 788 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_4146
timestamp 1745462530
transform 1 0 772 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4147
timestamp 1745462530
transform 1 0 3420 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_4148
timestamp 1745462530
transform 1 0 3412 0 1 2625
box -2 -2 2 2
use M2_M1  M2_M1_4149
timestamp 1745462530
transform 1 0 3404 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_4150
timestamp 1745462530
transform 1 0 3380 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_4151
timestamp 1745462530
transform 1 0 2788 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_4152
timestamp 1745462530
transform 1 0 2460 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_4153
timestamp 1745462530
transform 1 0 2452 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_4154
timestamp 1745462530
transform 1 0 1484 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_4155
timestamp 1745462530
transform 1 0 1180 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_4156
timestamp 1745462530
transform 1 0 1084 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_4157
timestamp 1745462530
transform 1 0 860 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_4158
timestamp 1745462530
transform 1 0 844 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_4159
timestamp 1745462530
transform 1 0 796 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_4160
timestamp 1745462530
transform 1 0 4108 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4161
timestamp 1745462530
transform 1 0 4092 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4162
timestamp 1745462530
transform 1 0 4004 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_4163
timestamp 1745462530
transform 1 0 4004 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_4164
timestamp 1745462530
transform 1 0 3988 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_4165
timestamp 1745462530
transform 1 0 3124 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_4166
timestamp 1745462530
transform 1 0 2428 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_4167
timestamp 1745462530
transform 1 0 2036 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4168
timestamp 1745462530
transform 1 0 1780 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_4169
timestamp 1745462530
transform 1 0 1612 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_4170
timestamp 1745462530
transform 1 0 636 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_4171
timestamp 1745462530
transform 1 0 564 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_4172
timestamp 1745462530
transform 1 0 548 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_4173
timestamp 1745462530
transform 1 0 3268 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_4174
timestamp 1745462530
transform 1 0 3252 0 1 1785
box -2 -2 2 2
use M2_M1  M2_M1_4175
timestamp 1745462530
transform 1 0 3236 0 1 1795
box -2 -2 2 2
use M2_M1  M2_M1_4176
timestamp 1745462530
transform 1 0 3236 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_4177
timestamp 1745462530
transform 1 0 3228 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_4178
timestamp 1745462530
transform 1 0 3228 0 1 2305
box -2 -2 2 2
use M2_M1  M2_M1_4179
timestamp 1745462530
transform 1 0 3220 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4180
timestamp 1745462530
transform 1 0 3220 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_4181
timestamp 1745462530
transform 1 0 3172 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_4182
timestamp 1745462530
transform 1 0 3124 0 1 1495
box -2 -2 2 2
use M2_M1  M2_M1_4183
timestamp 1745462530
transform 1 0 3020 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_4184
timestamp 1745462530
transform 1 0 2492 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_4185
timestamp 1745462530
transform 1 0 2252 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_4186
timestamp 1745462530
transform 1 0 1612 0 1 2715
box -2 -2 2 2
use M2_M1  M2_M1_4187
timestamp 1745462530
transform 1 0 1508 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_4188
timestamp 1745462530
transform 1 0 1332 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_4189
timestamp 1745462530
transform 1 0 620 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4190
timestamp 1745462530
transform 1 0 604 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_4191
timestamp 1745462530
transform 1 0 580 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_4192
timestamp 1745462530
transform 1 0 3692 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4193
timestamp 1745462530
transform 1 0 3668 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_4194
timestamp 1745462530
transform 1 0 3604 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_4195
timestamp 1745462530
transform 1 0 3524 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4196
timestamp 1745462530
transform 1 0 3220 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_4197
timestamp 1745462530
transform 1 0 2524 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_4198
timestamp 1745462530
transform 1 0 2508 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_4199
timestamp 1745462530
transform 1 0 2148 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_4200
timestamp 1745462530
transform 1 0 1972 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4201
timestamp 1745462530
transform 1 0 1036 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_4202
timestamp 1745462530
transform 1 0 772 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4203
timestamp 1745462530
transform 1 0 740 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_4204
timestamp 1745462530
transform 1 0 740 0 1 2155
box -2 -2 2 2
use M2_M1  M2_M1_4205
timestamp 1745462530
transform 1 0 740 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_4206
timestamp 1745462530
transform 1 0 740 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_4207
timestamp 1745462530
transform 1 0 3308 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_4208
timestamp 1745462530
transform 1 0 3292 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4209
timestamp 1745462530
transform 1 0 3220 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_4210
timestamp 1745462530
transform 1 0 3052 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_4211
timestamp 1745462530
transform 1 0 2764 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_4212
timestamp 1745462530
transform 1 0 2484 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_4213
timestamp 1745462530
transform 1 0 2388 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_4214
timestamp 1745462530
transform 1 0 1492 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4215
timestamp 1745462530
transform 1 0 1172 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4216
timestamp 1745462530
transform 1 0 1106 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_4217
timestamp 1745462530
transform 1 0 900 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_4218
timestamp 1745462530
transform 1 0 900 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_4219
timestamp 1745462530
transform 1 0 876 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_4220
timestamp 1745462530
transform 1 0 4020 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4221
timestamp 1745462530
transform 1 0 4012 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4222
timestamp 1745462530
transform 1 0 4004 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_4223
timestamp 1745462530
transform 1 0 3956 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_4224
timestamp 1745462530
transform 1 0 3932 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_4225
timestamp 1745462530
transform 1 0 3156 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_4226
timestamp 1745462530
transform 1 0 2540 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_4227
timestamp 1745462530
transform 1 0 2052 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4228
timestamp 1745462530
transform 1 0 1844 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_4229
timestamp 1745462530
transform 1 0 1740 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_4230
timestamp 1745462530
transform 1 0 604 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_4231
timestamp 1745462530
transform 1 0 532 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_4232
timestamp 1745462530
transform 1 0 532 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_4233
timestamp 1745462530
transform 1 0 524 0 1 2155
box -2 -2 2 2
use M2_M1  M2_M1_4234
timestamp 1745462530
transform 1 0 516 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_4235
timestamp 1745462530
transform 1 0 3124 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_4236
timestamp 1745462530
transform 1 0 3108 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_4237
timestamp 1745462530
transform 1 0 3092 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4238
timestamp 1745462530
transform 1 0 3092 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_4239
timestamp 1745462530
transform 1 0 3028 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_4240
timestamp 1745462530
transform 1 0 2564 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_4241
timestamp 1745462530
transform 1 0 2220 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_4242
timestamp 1745462530
transform 1 0 1652 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4243
timestamp 1745462530
transform 1 0 1548 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_4244
timestamp 1745462530
transform 1 0 1364 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4245
timestamp 1745462530
transform 1 0 652 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_4246
timestamp 1745462530
transform 1 0 596 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_4247
timestamp 1745462530
transform 1 0 588 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_4248
timestamp 1745462530
transform 1 0 3652 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_4249
timestamp 1745462530
transform 1 0 3636 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4250
timestamp 1745462530
transform 1 0 3588 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_4251
timestamp 1745462530
transform 1 0 3508 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4252
timestamp 1745462530
transform 1 0 3204 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_4253
timestamp 1745462530
transform 1 0 2556 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4254
timestamp 1745462530
transform 1 0 2508 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_4255
timestamp 1745462530
transform 1 0 2132 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_4256
timestamp 1745462530
transform 1 0 1932 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4257
timestamp 1745462530
transform 1 0 1012 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_4258
timestamp 1745462530
transform 1 0 756 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4259
timestamp 1745462530
transform 1 0 740 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4260
timestamp 1745462530
transform 1 0 724 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_4261
timestamp 1745462530
transform 1 0 724 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_4262
timestamp 1745462530
transform 1 0 3292 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_4263
timestamp 1745462530
transform 1 0 3276 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4264
timestamp 1745462530
transform 1 0 3188 0 1 1945
box -2 -2 2 2
use M2_M1  M2_M1_4265
timestamp 1745462530
transform 1 0 3116 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_4266
timestamp 1745462530
transform 1 0 3100 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_4267
timestamp 1745462530
transform 1 0 3036 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_4268
timestamp 1745462530
transform 1 0 2748 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_4269
timestamp 1745462530
transform 1 0 2588 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4270
timestamp 1745462530
transform 1 0 2372 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_4271
timestamp 1745462530
transform 1 0 1468 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4272
timestamp 1745462530
transform 1 0 1156 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4273
timestamp 1745462530
transform 1 0 1052 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_4274
timestamp 1745462530
transform 1 0 932 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_4275
timestamp 1745462530
transform 1 0 916 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_4276
timestamp 1745462530
transform 1 0 884 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_4277
timestamp 1745462530
transform 1 0 884 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_4278
timestamp 1745462530
transform 1 0 860 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_4279
timestamp 1745462530
transform 1 0 3980 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4280
timestamp 1745462530
transform 1 0 3980 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_4281
timestamp 1745462530
transform 1 0 3972 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4282
timestamp 1745462530
transform 1 0 3940 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_4283
timestamp 1745462530
transform 1 0 3908 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_4284
timestamp 1745462530
transform 1 0 3908 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_4285
timestamp 1745462530
transform 1 0 3900 0 1 2145
box -2 -2 2 2
use M2_M1  M2_M1_4286
timestamp 1745462530
transform 1 0 3900 0 1 1945
box -2 -2 2 2
use M2_M1  M2_M1_4287
timestamp 1745462530
transform 1 0 3140 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_4288
timestamp 1745462530
transform 1 0 2612 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_4289
timestamp 1745462530
transform 1 0 2036 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4290
timestamp 1745462530
transform 1 0 1828 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_4291
timestamp 1745462530
transform 1 0 1724 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_4292
timestamp 1745462530
transform 1 0 588 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_4293
timestamp 1745462530
transform 1 0 516 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_4294
timestamp 1745462530
transform 1 0 476 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_4295
timestamp 1745462530
transform 1 0 3084 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_4296
timestamp 1745462530
transform 1 0 3076 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_4297
timestamp 1745462530
transform 1 0 3060 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4298
timestamp 1745462530
transform 1 0 3060 0 1 1495
box -2 -2 2 2
use M2_M1  M2_M1_4299
timestamp 1745462530
transform 1 0 3012 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_4300
timestamp 1745462530
transform 1 0 2628 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4301
timestamp 1745462530
transform 1 0 2204 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_4302
timestamp 1745462530
transform 1 0 1636 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4303
timestamp 1745462530
transform 1 0 1524 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_4304
timestamp 1745462530
transform 1 0 1348 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4305
timestamp 1745462530
transform 1 0 612 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_4306
timestamp 1745462530
transform 1 0 580 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_4307
timestamp 1745462530
transform 1 0 572 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_4308
timestamp 1745462530
transform 1 0 3124 0 1 3345
box -2 -2 2 2
use M2_M1  M2_M1_4309
timestamp 1745462530
transform 1 0 2804 0 1 3425
box -2 -2 2 2
use M2_M1  M2_M1_4310
timestamp 1745462530
transform 1 0 2228 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_4311
timestamp 1745462530
transform 1 0 2212 0 1 3225
box -2 -2 2 2
use M2_M1  M2_M1_4312
timestamp 1745462530
transform 1 0 2164 0 1 3225
box -2 -2 2 2
use M2_M1  M2_M1_4313
timestamp 1745462530
transform 1 0 2164 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_4314
timestamp 1745462530
transform 1 0 3852 0 1 3225
box -2 -2 2 2
use M2_M1  M2_M1_4315
timestamp 1745462530
transform 1 0 3836 0 1 3315
box -2 -2 2 2
use M2_M1  M2_M1_4316
timestamp 1745462530
transform 1 0 3820 0 1 3225
box -2 -2 2 2
use M2_M1  M2_M1_4317
timestamp 1745462530
transform 1 0 3772 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_4318
timestamp 1745462530
transform 1 0 3772 0 1 3225
box -2 -2 2 2
use M2_M1  M2_M1_4319
timestamp 1745462530
transform 1 0 3724 0 1 3315
box -2 -2 2 2
use M2_M1  M2_M1_4320
timestamp 1745462530
transform 1 0 3684 0 1 3225
box -2 -2 2 2
use M2_M1  M2_M1_4321
timestamp 1745462530
transform 1 0 2092 0 1 3155
box -2 -2 2 2
use M2_M1  M2_M1_4322
timestamp 1745462530
transform 1 0 2004 0 1 3315
box -2 -2 2 2
use M2_M1  M2_M1_4323
timestamp 1745462530
transform 1 0 1940 0 1 3225
box -2 -2 2 2
use M2_M1  M2_M1_4324
timestamp 1745462530
transform 1 0 1884 0 1 3315
box -2 -2 2 2
use M2_M1  M2_M1_4325
timestamp 1745462530
transform 1 0 1844 0 1 3315
box -2 -2 2 2
use M2_M1  M2_M1_4326
timestamp 1745462530
transform 1 0 1844 0 1 3225
box -2 -2 2 2
use M2_M1  M2_M1_4327
timestamp 1745462530
transform 1 0 3868 0 1 3425
box -2 -2 2 2
use M2_M1  M2_M1_4328
timestamp 1745462530
transform 1 0 3836 0 1 3425
box -2 -2 2 2
use M2_M1  M2_M1_4329
timestamp 1745462530
transform 1 0 3812 0 1 3515
box -2 -2 2 2
use M2_M1  M2_M1_4330
timestamp 1745462530
transform 1 0 3796 0 1 3315
box -2 -2 2 2
use M2_M1  M2_M1_4331
timestamp 1745462530
transform 1 0 3764 0 1 3425
box -2 -2 2 2
use M2_M1  M2_M1_4332
timestamp 1745462530
transform 1 0 3020 0 1 3425
box -2 -2 2 2
use M2_M1  M2_M1_4333
timestamp 1745462530
transform 1 0 2652 0 1 3315
box -2 -2 2 2
use M2_M1  M2_M1_4334
timestamp 1745462530
transform 1 0 2068 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_4335
timestamp 1745462530
transform 1 0 2020 0 1 3515
box -2 -2 2 2
use M2_M1  M2_M1_4336
timestamp 1745462530
transform 1 0 2020 0 1 3435
box -2 -2 2 2
use M2_M1  M2_M1_4337
timestamp 1745462530
transform 1 0 2004 0 1 3425
box -2 -2 2 2
use M2_M1  M2_M1_4338
timestamp 1745462530
transform 1 0 1996 0 1 3225
box -2 -2 2 2
use M2_M1  M2_M1_4339
timestamp 1745462530
transform 1 0 1932 0 1 3515
box -2 -2 2 2
use M2_M1  M2_M1_4340
timestamp 1745462530
transform 1 0 1924 0 1 3425
box -2 -2 2 2
use M2_M1  M2_M1_4341
timestamp 1745462530
transform 1 0 3884 0 1 3515
box -2 -2 2 2
use M2_M1  M2_M1_4342
timestamp 1745462530
transform 1 0 3828 0 1 3625
box -2 -2 2 2
use M2_M1  M2_M1_4343
timestamp 1745462530
transform 1 0 3796 0 1 3625
box -2 -2 2 2
use M2_M1  M2_M1_4344
timestamp 1745462530
transform 1 0 3772 0 1 3515
box -2 -2 2 2
use M2_M1  M2_M1_4345
timestamp 1745462530
transform 1 0 3756 0 1 3715
box -2 -2 2 2
use M2_M1  M2_M1_4346
timestamp 1745462530
transform 1 0 3756 0 1 3625
box -2 -2 2 2
use M2_M1  M2_M1_4347
timestamp 1745462530
transform 1 0 3684 0 1 3715
box -2 -2 2 2
use M2_M1  M2_M1_4348
timestamp 1745462530
transform 1 0 2948 0 1 3715
box -2 -2 2 2
use M2_M1  M2_M1_4349
timestamp 1745462530
transform 1 0 2924 0 1 3625
box -2 -2 2 2
use M2_M1  M2_M1_4350
timestamp 1745462530
transform 1 0 2740 0 1 3625
box -2 -2 2 2
use M2_M1  M2_M1_4351
timestamp 1745462530
transform 1 0 2484 0 1 3715
box -2 -2 2 2
use M2_M1  M2_M1_4352
timestamp 1745462530
transform 1 0 2276 0 1 3625
box -2 -2 2 2
use M2_M1  M2_M1_4353
timestamp 1745462530
transform 1 0 2228 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_4354
timestamp 1745462530
transform 1 0 3252 0 1 3715
box -2 -2 2 2
use M2_M1  M2_M1_4355
timestamp 1745462530
transform 1 0 3220 0 1 3715
box -2 -2 2 2
use M2_M1  M2_M1_4356
timestamp 1745462530
transform 1 0 3204 0 1 3625
box -2 -2 2 2
use M2_M1  M2_M1_4357
timestamp 1745462530
transform 1 0 3180 0 1 3715
box -2 -2 2 2
use M2_M1  M2_M1_4358
timestamp 1745462530
transform 1 0 3148 0 1 3715
box -2 -2 2 2
use M2_M1  M2_M1_4359
timestamp 1745462530
transform 1 0 3012 0 1 3715
box -2 -2 2 2
use M2_M1  M2_M1_4360
timestamp 1745462530
transform 1 0 2796 0 1 3625
box -2 -2 2 2
use M2_M1  M2_M1_4361
timestamp 1745462530
transform 1 0 2764 0 1 3715
box -2 -2 2 2
use M2_M1  M2_M1_4362
timestamp 1745462530
transform 1 0 2452 0 1 3715
box -2 -2 2 2
use M2_M1  M2_M1_4363
timestamp 1745462530
transform 1 0 2380 0 1 3715
box -2 -2 2 2
use M2_M1  M2_M1_4364
timestamp 1745462530
transform 1 0 2300 0 1 3715
box -2 -2 2 2
use M2_M1  M2_M1_4365
timestamp 1745462530
transform 1 0 2244 0 1 3715
box -2 -2 2 2
use M2_M1  M2_M1_4366
timestamp 1745462530
transform 1 0 2244 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_4367
timestamp 1745462530
transform 1 0 3620 0 1 3625
box -2 -2 2 2
use M2_M1  M2_M1_4368
timestamp 1745462530
transform 1 0 3548 0 1 3645
box -2 -2 2 2
use M2_M1  M2_M1_4369
timestamp 1745462530
transform 1 0 3452 0 1 3625
box -2 -2 2 2
use M2_M1  M2_M1_4370
timestamp 1745462530
transform 1 0 3444 0 1 3715
box -2 -2 2 2
use M2_M1  M2_M1_4371
timestamp 1745462530
transform 1 0 3372 0 1 3715
box -2 -2 2 2
use M2_M1  M2_M1_4372
timestamp 1745462530
transform 1 0 3372 0 1 3625
box -2 -2 2 2
use M2_M1  M2_M1_4373
timestamp 1745462530
transform 1 0 3148 0 1 3625
box -2 -2 2 2
use M2_M1  M2_M1_4374
timestamp 1745462530
transform 1 0 3084 0 1 3715
box -2 -2 2 2
use M2_M1  M2_M1_4375
timestamp 1745462530
transform 1 0 2996 0 1 3625
box -2 -2 2 2
use M2_M1  M2_M1_4376
timestamp 1745462530
transform 1 0 2852 0 1 3625
box -2 -2 2 2
use M2_M1  M2_M1_4377
timestamp 1745462530
transform 1 0 2364 0 1 3625
box -2 -2 2 2
use M2_M1  M2_M1_4378
timestamp 1745462530
transform 1 0 2204 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_4379
timestamp 1745462530
transform 1 0 2180 0 1 3625
box -2 -2 2 2
use M2_M1  M2_M1_4380
timestamp 1745462530
transform 1 0 2132 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_4381
timestamp 1745462530
transform 1 0 2124 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_4382
timestamp 1745462530
transform 1 0 2068 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_4383
timestamp 1745462530
transform 1 0 2052 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_4384
timestamp 1745462530
transform 1 0 2220 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_4385
timestamp 1745462530
transform 1 0 2212 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_4386
timestamp 1745462530
transform 1 0 2196 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_4387
timestamp 1745462530
transform 1 0 2188 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_4388
timestamp 1745462530
transform 1 0 2692 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4389
timestamp 1745462530
transform 1 0 2668 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4390
timestamp 1745462530
transform 1 0 2308 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_4391
timestamp 1745462530
transform 1 0 2260 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_4392
timestamp 1745462530
transform 1 0 2164 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_4393
timestamp 1745462530
transform 1 0 1580 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_4394
timestamp 1745462530
transform 1 0 1500 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_4395
timestamp 1745462530
transform 1 0 2988 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_4396
timestamp 1745462530
transform 1 0 2948 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4397
timestamp 1745462530
transform 1 0 2684 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_4398
timestamp 1745462530
transform 1 0 1180 0 1 3035
box -2 -2 2 2
use M2_M1  M2_M1_4399
timestamp 1745462530
transform 1 0 900 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_4400
timestamp 1745462530
transform 1 0 1516 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_4401
timestamp 1745462530
transform 1 0 1500 0 1 2305
box -2 -2 2 2
use M2_M1  M2_M1_4402
timestamp 1745462530
transform 1 0 1484 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_4403
timestamp 1745462530
transform 1 0 1476 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_4404
timestamp 1745462530
transform 1 0 1460 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4405
timestamp 1745462530
transform 1 0 716 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_4406
timestamp 1745462530
transform 1 0 644 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_4407
timestamp 1745462530
transform 1 0 524 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_4408
timestamp 1745462530
transform 1 0 484 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_4409
timestamp 1745462530
transform 1 0 1612 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_4410
timestamp 1745462530
transform 1 0 1500 0 1 1315
box -2 -2 2 2
use M2_M1  M2_M1_4411
timestamp 1745462530
transform 1 0 1476 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_4412
timestamp 1745462530
transform 1 0 1460 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_4413
timestamp 1745462530
transform 1 0 1092 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_4414
timestamp 1745462530
transform 1 0 1044 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_4415
timestamp 1745462530
transform 1 0 988 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_4416
timestamp 1745462530
transform 1 0 932 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_4417
timestamp 1745462530
transform 1 0 3252 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_4418
timestamp 1745462530
transform 1 0 3164 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_4419
timestamp 1745462530
transform 1 0 2836 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_4420
timestamp 1745462530
transform 1 0 2796 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_4421
timestamp 1745462530
transform 1 0 2740 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_4422
timestamp 1745462530
transform 1 0 2724 0 1 1035
box -2 -2 2 2
use M2_M1  M2_M1_4423
timestamp 1745462530
transform 1 0 2716 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_4424
timestamp 1745462530
transform 1 0 2708 0 1 1035
box -2 -2 2 2
use M2_M1  M2_M1_4425
timestamp 1745462530
transform 1 0 2404 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_4426
timestamp 1745462530
transform 1 0 2340 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_4427
timestamp 1745462530
transform 1 0 2308 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_4428
timestamp 1745462530
transform 1 0 3452 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_4429
timestamp 1745462530
transform 1 0 3412 0 1 1155
box -2 -2 2 2
use M2_M1  M2_M1_4430
timestamp 1745462530
transform 1 0 3388 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_4431
timestamp 1745462530
transform 1 0 2180 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_4432
timestamp 1745462530
transform 1 0 2036 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_4433
timestamp 1745462530
transform 1 0 3148 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_4434
timestamp 1745462530
transform 1 0 3036 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_4435
timestamp 1745462530
transform 1 0 2996 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_4436
timestamp 1745462530
transform 1 0 2932 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_4437
timestamp 1745462530
transform 1 0 3092 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_4438
timestamp 1745462530
transform 1 0 3060 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_4439
timestamp 1745462530
transform 1 0 3044 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_4440
timestamp 1745462530
transform 1 0 2844 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_4441
timestamp 1745462530
transform 1 0 2724 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_4442
timestamp 1745462530
transform 1 0 3004 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_4443
timestamp 1745462530
transform 1 0 3004 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_4444
timestamp 1745462530
transform 1 0 2956 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_4445
timestamp 1745462530
transform 1 0 4012 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_4446
timestamp 1745462530
transform 1 0 3972 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_4447
timestamp 1745462530
transform 1 0 3844 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_4448
timestamp 1745462530
transform 1 0 3836 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4449
timestamp 1745462530
transform 1 0 3836 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_4450
timestamp 1745462530
transform 1 0 3804 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_4451
timestamp 1745462530
transform 1 0 3772 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_4452
timestamp 1745462530
transform 1 0 2868 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_4453
timestamp 1745462530
transform 1 0 2676 0 1 2995
box -2 -2 2 2
use M2_M1  M2_M1_4454
timestamp 1745462530
transform 1 0 2660 0 1 2995
box -2 -2 2 2
use M2_M1  M2_M1_4455
timestamp 1745462530
transform 1 0 2540 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_4456
timestamp 1745462530
transform 1 0 2468 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_4457
timestamp 1745462530
transform 1 0 2452 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_4458
timestamp 1745462530
transform 1 0 1284 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_4459
timestamp 1745462530
transform 1 0 1276 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_4460
timestamp 1745462530
transform 1 0 2052 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_4461
timestamp 1745462530
transform 1 0 1884 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_4462
timestamp 1745462530
transform 1 0 1452 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_4463
timestamp 1745462530
transform 1 0 1396 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_4464
timestamp 1745462530
transform 1 0 1364 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4465
timestamp 1745462530
transform 1 0 1284 0 1 555
box -2 -2 2 2
use M2_M1  M2_M1_4466
timestamp 1745462530
transform 1 0 1268 0 1 555
box -2 -2 2 2
use M2_M1  M2_M1_4467
timestamp 1745462530
transform 1 0 1244 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_4468
timestamp 1745462530
transform 1 0 1212 0 1 485
box -2 -2 2 2
use M2_M1  M2_M1_4469
timestamp 1745462530
transform 1 0 980 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4470
timestamp 1745462530
transform 1 0 956 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4471
timestamp 1745462530
transform 1 0 724 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4472
timestamp 1745462530
transform 1 0 516 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4473
timestamp 1745462530
transform 1 0 500 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_4474
timestamp 1745462530
transform 1 0 460 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4475
timestamp 1745462530
transform 1 0 452 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_4476
timestamp 1745462530
transform 1 0 452 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_4477
timestamp 1745462530
transform 1 0 444 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_4478
timestamp 1745462530
transform 1 0 428 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_4479
timestamp 1745462530
transform 1 0 420 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_4480
timestamp 1745462530
transform 1 0 2612 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_4481
timestamp 1745462530
transform 1 0 2572 0 1 2105
box -2 -2 2 2
use M2_M1  M2_M1_4482
timestamp 1745462530
transform 1 0 2436 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_4483
timestamp 1745462530
transform 1 0 1740 0 1 2085
box -2 -2 2 2
use M2_M1  M2_M1_4484
timestamp 1745462530
transform 1 0 1380 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_4485
timestamp 1745462530
transform 1 0 1364 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_4486
timestamp 1745462530
transform 1 0 1300 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_4487
timestamp 1745462530
transform 1 0 1468 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_4488
timestamp 1745462530
transform 1 0 1412 0 1 2515
box -2 -2 2 2
use M2_M1  M2_M1_4489
timestamp 1745462530
transform 1 0 1412 0 1 2455
box -2 -2 2 2
use M2_M1  M2_M1_4490
timestamp 1745462530
transform 1 0 1412 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_4491
timestamp 1745462530
transform 1 0 1404 0 1 2305
box -2 -2 2 2
use M2_M1  M2_M1_4492
timestamp 1745462530
transform 1 0 1388 0 1 2455
box -2 -2 2 2
use M2_M1  M2_M1_4493
timestamp 1745462530
transform 1 0 1388 0 1 2345
box -2 -2 2 2
use M2_M1  M2_M1_4494
timestamp 1745462530
transform 1 0 1380 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_4495
timestamp 1745462530
transform 1 0 1100 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_4496
timestamp 1745462530
transform 1 0 1324 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_4497
timestamp 1745462530
transform 1 0 1316 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_4498
timestamp 1745462530
transform 1 0 1260 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_4499
timestamp 1745462530
transform 1 0 1020 0 1 2515
box -2 -2 2 2
use M2_M1  M2_M1_4500
timestamp 1745462530
transform 1 0 980 0 1 2515
box -2 -2 2 2
use M2_M1  M2_M1_4501
timestamp 1745462530
transform 1 0 740 0 1 2515
box -2 -2 2 2
use M2_M1  M2_M1_4502
timestamp 1745462530
transform 1 0 540 0 1 2515
box -2 -2 2 2
use M2_M1  M2_M1_4503
timestamp 1745462530
transform 1 0 540 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_4504
timestamp 1745462530
transform 1 0 476 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_4505
timestamp 1745462530
transform 1 0 460 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_4506
timestamp 1745462530
transform 1 0 460 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_4507
timestamp 1745462530
transform 1 0 436 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_4508
timestamp 1745462530
transform 1 0 3820 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_4509
timestamp 1745462530
transform 1 0 3796 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_4510
timestamp 1745462530
transform 1 0 3604 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_4511
timestamp 1745462530
transform 1 0 3572 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_4512
timestamp 1745462530
transform 1 0 3532 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_4513
timestamp 1745462530
transform 1 0 2676 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_4514
timestamp 1745462530
transform 1 0 2660 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_4515
timestamp 1745462530
transform 1 0 2652 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_4516
timestamp 1745462530
transform 1 0 2636 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_4517
timestamp 1745462530
transform 1 0 2596 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_4518
timestamp 1745462530
transform 1 0 2004 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_4519
timestamp 1745462530
transform 1 0 1932 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_4520
timestamp 1745462530
transform 1 0 4028 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_4521
timestamp 1745462530
transform 1 0 3988 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_4522
timestamp 1745462530
transform 1 0 3884 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_4523
timestamp 1745462530
transform 1 0 3876 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_4524
timestamp 1745462530
transform 1 0 3868 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_4525
timestamp 1745462530
transform 1 0 2604 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_4526
timestamp 1745462530
transform 1 0 1468 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_4527
timestamp 1745462530
transform 1 0 1396 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_4528
timestamp 1745462530
transform 1 0 1268 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_4529
timestamp 1745462530
transform 1 0 1236 0 1 3025
box -2 -2 2 2
use M2_M1  M2_M1_4530
timestamp 1745462530
transform 1 0 1068 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_4531
timestamp 1745462530
transform 1 0 1004 0 1 3225
box -2 -2 2 2
use M2_M1  M2_M1_4532
timestamp 1745462530
transform 1 0 964 0 1 3225
box -2 -2 2 2
use M2_M1  M2_M1_4533
timestamp 1745462530
transform 1 0 1852 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_4534
timestamp 1745462530
transform 1 0 1844 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_4535
timestamp 1745462530
transform 1 0 1772 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_4536
timestamp 1745462530
transform 1 0 1764 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_4537
timestamp 1745462530
transform 1 0 1676 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_4538
timestamp 1745462530
transform 1 0 1596 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_4539
timestamp 1745462530
transform 1 0 3468 0 1 1345
box -2 -2 2 2
use M2_M1  M2_M1_4540
timestamp 1745462530
transform 1 0 3468 0 1 1145
box -2 -2 2 2
use M2_M1  M2_M1_4541
timestamp 1745462530
transform 1 0 3404 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_4542
timestamp 1745462530
transform 1 0 3276 0 1 995
box -2 -2 2 2
use M2_M1  M2_M1_4543
timestamp 1745462530
transform 1 0 3196 0 1 985
box -2 -2 2 2
use M2_M1  M2_M1_4544
timestamp 1745462530
transform 1 0 3132 0 1 2745
box -2 -2 2 2
use M2_M1  M2_M1_4545
timestamp 1745462530
transform 1 0 3084 0 1 2595
box -2 -2 2 2
use M2_M1  M2_M1_4546
timestamp 1745462530
transform 1 0 3084 0 1 2145
box -2 -2 2 2
use M2_M1  M2_M1_4547
timestamp 1745462530
transform 1 0 3044 0 1 2745
box -2 -2 2 2
use M2_M1  M2_M1_4548
timestamp 1745462530
transform 1 0 2868 0 1 995
box -2 -2 2 2
use M2_M1  M2_M1_4549
timestamp 1745462530
transform 1 0 2820 0 1 995
box -2 -2 2 2
use M2_M1  M2_M1_4550
timestamp 1745462530
transform 1 0 2780 0 1 1345
box -2 -2 2 2
use M2_M1  M2_M1_4551
timestamp 1745462530
transform 1 0 2428 0 1 2745
box -2 -2 2 2
use M2_M1  M2_M1_4552
timestamp 1745462530
transform 1 0 2340 0 1 995
box -2 -2 2 2
use M2_M1  M2_M1_4553
timestamp 1745462530
transform 1 0 2172 0 1 3145
box -2 -2 2 2
use M2_M1  M2_M1_4554
timestamp 1745462530
transform 1 0 1564 0 1 1345
box -2 -2 2 2
use M2_M1  M2_M1_4555
timestamp 1745462530
transform 1 0 1540 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_4556
timestamp 1745462530
transform 1 0 1492 0 1 1145
box -2 -2 2 2
use M2_M1  M2_M1_4557
timestamp 1745462530
transform 1 0 1492 0 1 995
box -2 -2 2 2
use M2_M1  M2_M1_4558
timestamp 1745462530
transform 1 0 1156 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_4559
timestamp 1745462530
transform 1 0 1124 0 1 995
box -2 -2 2 2
use M2_M1  M2_M1_4560
timestamp 1745462530
transform 1 0 1108 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_4561
timestamp 1745462530
transform 1 0 1076 0 1 1195
box -2 -2 2 2
use M2_M1  M2_M1_4562
timestamp 1745462530
transform 1 0 1020 0 1 1145
box -2 -2 2 2
use M2_M1  M2_M1_4563
timestamp 1745462530
transform 1 0 3820 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_4564
timestamp 1745462530
transform 1 0 2780 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_4565
timestamp 1745462530
transform 1 0 2156 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_4566
timestamp 1745462530
transform 1 0 1580 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_4567
timestamp 1745462530
transform 1 0 1556 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_4568
timestamp 1745462530
transform 1 0 4220 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_4569
timestamp 1745462530
transform 1 0 4212 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_4570
timestamp 1745462530
transform 1 0 4212 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_4571
timestamp 1745462530
transform 1 0 4196 0 1 3155
box -2 -2 2 2
use M2_M1  M2_M1_4572
timestamp 1745462530
transform 1 0 4028 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_4573
timestamp 1745462530
transform 1 0 4028 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_4574
timestamp 1745462530
transform 1 0 3948 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_4575
timestamp 1745462530
transform 1 0 2172 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_4576
timestamp 1745462530
transform 1 0 1764 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_4577
timestamp 1745462530
transform 1 0 1700 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_4578
timestamp 1745462530
transform 1 0 1652 0 1 4005
box -2 -2 2 2
use M2_M1  M2_M1_4579
timestamp 1745462530
transform 1 0 1644 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_4580
timestamp 1745462530
transform 1 0 1644 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_4581
timestamp 1745462530
transform 1 0 4132 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_4582
timestamp 1745462530
transform 1 0 4044 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_4583
timestamp 1745462530
transform 1 0 4044 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_4584
timestamp 1745462530
transform 1 0 3964 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_4585
timestamp 1745462530
transform 1 0 3956 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_4586
timestamp 1745462530
transform 1 0 2852 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_4587
timestamp 1745462530
transform 1 0 2676 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_4588
timestamp 1745462530
transform 1 0 2148 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_4589
timestamp 1745462530
transform 1 0 2012 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_4590
timestamp 1745462530
transform 1 0 2012 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_4591
timestamp 1745462530
transform 1 0 1980 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_4592
timestamp 1745462530
transform 1 0 1924 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_4593
timestamp 1745462530
transform 1 0 1860 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_4594
timestamp 1745462530
transform 1 0 4300 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_4595
timestamp 1745462530
transform 1 0 4228 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_4596
timestamp 1745462530
transform 1 0 4212 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_4597
timestamp 1745462530
transform 1 0 3852 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_4598
timestamp 1745462530
transform 1 0 3756 0 1 4005
box -2 -2 2 2
use M2_M1  M2_M1_4599
timestamp 1745462530
transform 1 0 3708 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_4600
timestamp 1745462530
transform 1 0 3684 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_4601
timestamp 1745462530
transform 1 0 2980 0 1 4005
box -2 -2 2 2
use M2_M1  M2_M1_4602
timestamp 1745462530
transform 1 0 2916 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_4603
timestamp 1745462530
transform 1 0 2588 0 1 4005
box -2 -2 2 2
use M2_M1  M2_M1_4604
timestamp 1745462530
transform 1 0 2484 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_4605
timestamp 1745462530
transform 1 0 2292 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_4606
timestamp 1745462530
transform 1 0 2284 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_4607
timestamp 1745462530
transform 1 0 3500 0 1 4005
box -2 -2 2 2
use M2_M1  M2_M1_4608
timestamp 1745462530
transform 1 0 3484 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_4609
timestamp 1745462530
transform 1 0 3380 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_4610
timestamp 1745462530
transform 1 0 3228 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_4611
timestamp 1745462530
transform 1 0 3172 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_4612
timestamp 1745462530
transform 1 0 3012 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_4613
timestamp 1745462530
transform 1 0 2740 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_4614
timestamp 1745462530
transform 1 0 2644 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_4615
timestamp 1745462530
transform 1 0 2404 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_4616
timestamp 1745462530
transform 1 0 2372 0 1 4005
box -2 -2 2 2
use M2_M1  M2_M1_4617
timestamp 1745462530
transform 1 0 2212 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_4618
timestamp 1745462530
transform 1 0 2172 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_4619
timestamp 1745462530
transform 1 0 3628 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_4620
timestamp 1745462530
transform 1 0 3596 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_4621
timestamp 1745462530
transform 1 0 3588 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_4622
timestamp 1745462530
transform 1 0 3356 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_4623
timestamp 1745462530
transform 1 0 3348 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_4624
timestamp 1745462530
transform 1 0 3276 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_4625
timestamp 1745462530
transform 1 0 3140 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_4626
timestamp 1745462530
transform 1 0 3116 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_4627
timestamp 1745462530
transform 1 0 3084 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_4628
timestamp 1745462530
transform 1 0 2836 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_4629
timestamp 1745462530
transform 1 0 2380 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_4630
timestamp 1745462530
transform 1 0 2260 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_4631
timestamp 1745462530
transform 1 0 2068 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_4632
timestamp 1745462530
transform 1 0 804 0 1 4115
box -2 -2 2 2
use M2_M1  M2_M1_4633
timestamp 1745462530
transform 1 0 628 0 1 4105
box -2 -2 2 2
use M2_M1  M2_M1_4634
timestamp 1745462530
transform 1 0 4100 0 1 4225
box -2 -2 2 2
use M2_M1  M2_M1_4635
timestamp 1745462530
transform 1 0 4068 0 1 4115
box -2 -2 2 2
use M2_M1  M2_M1_4636
timestamp 1745462530
transform 1 0 3988 0 1 4025
box -2 -2 2 2
use M2_M1  M2_M1_4637
timestamp 1745462530
transform 1 0 3980 0 1 4115
box -2 -2 2 2
use M2_M1  M2_M1_4638
timestamp 1745462530
transform 1 0 2908 0 1 4225
box -2 -2 2 2
use M2_M1  M2_M1_4639
timestamp 1745462530
transform 1 0 2668 0 1 4225
box -2 -2 2 2
use M2_M1  M2_M1_4640
timestamp 1745462530
transform 1 0 1940 0 1 4225
box -2 -2 2 2
use M2_M1  M2_M1_4641
timestamp 1745462530
transform 1 0 1892 0 1 4115
box -2 -2 2 2
use M2_M1  M2_M1_4642
timestamp 1745462530
transform 1 0 1348 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_4643
timestamp 1745462530
transform 1 0 1348 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_4644
timestamp 1745462530
transform 1 0 1324 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_4645
timestamp 1745462530
transform 1 0 1260 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_4646
timestamp 1745462530
transform 1 0 1084 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_4647
timestamp 1745462530
transform 1 0 884 0 1 4005
box -2 -2 2 2
use M2_M1  M2_M1_4648
timestamp 1745462530
transform 1 0 1164 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_4649
timestamp 1745462530
transform 1 0 1132 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_4650
timestamp 1745462530
transform 1 0 1012 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_4651
timestamp 1745462530
transform 1 0 916 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_4652
timestamp 1745462530
transform 1 0 908 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_4653
timestamp 1745462530
transform 1 0 900 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_4654
timestamp 1745462530
transform 1 0 884 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_4655
timestamp 1745462530
transform 1 0 3548 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_4656
timestamp 1745462530
transform 1 0 3548 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_4657
timestamp 1745462530
transform 1 0 3524 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_4658
timestamp 1745462530
transform 1 0 3420 0 1 4105
box -2 -2 2 2
use M2_M1  M2_M1_4659
timestamp 1745462530
transform 1 0 3036 0 1 4035
box -2 -2 2 2
use M2_M1  M2_M1_4660
timestamp 1745462530
transform 1 0 2668 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_4661
timestamp 1745462530
transform 1 0 2540 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_4662
timestamp 1745462530
transform 1 0 2340 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_4663
timestamp 1745462530
transform 1 0 2228 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_4664
timestamp 1745462530
transform 1 0 2180 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_4665
timestamp 1745462530
transform 1 0 3556 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_4666
timestamp 1745462530
transform 1 0 3508 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_4667
timestamp 1745462530
transform 1 0 3492 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_4668
timestamp 1745462530
transform 1 0 3276 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_4669
timestamp 1745462530
transform 1 0 3068 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_4670
timestamp 1745462530
transform 1 0 2796 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_4671
timestamp 1745462530
transform 1 0 2548 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_4672
timestamp 1745462530
transform 1 0 2364 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_4673
timestamp 1745462530
transform 1 0 2188 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_4674
timestamp 1745462530
transform 1 0 2140 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_4675
timestamp 1745462530
transform 1 0 3076 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_4676
timestamp 1745462530
transform 1 0 3068 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_4677
timestamp 1745462530
transform 1 0 3028 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_4678
timestamp 1745462530
transform 1 0 2996 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_4679
timestamp 1745462530
transform 1 0 2956 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_4680
timestamp 1745462530
transform 1 0 2924 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_4681
timestamp 1745462530
transform 1 0 2924 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_4682
timestamp 1745462530
transform 1 0 2900 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_4683
timestamp 1745462530
transform 1 0 2900 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_4684
timestamp 1745462530
transform 1 0 2764 0 1 3825
box -2 -2 2 2
use M2_M1  M2_M1_4685
timestamp 1745462530
transform 1 0 2036 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_4686
timestamp 1745462530
transform 1 0 3588 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_4687
timestamp 1745462530
transform 1 0 3572 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_4688
timestamp 1745462530
transform 1 0 3540 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_4689
timestamp 1745462530
transform 1 0 3508 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_4690
timestamp 1745462530
transform 1 0 3508 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_4691
timestamp 1745462530
transform 1 0 3476 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_4692
timestamp 1745462530
transform 1 0 3356 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_4693
timestamp 1745462530
transform 1 0 3292 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_4694
timestamp 1745462530
transform 1 0 3284 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_4695
timestamp 1745462530
transform 1 0 3204 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_4696
timestamp 1745462530
transform 1 0 2428 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_4697
timestamp 1745462530
transform 1 0 2668 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_4698
timestamp 1745462530
transform 1 0 2628 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_4699
timestamp 1745462530
transform 1 0 2564 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_4700
timestamp 1745462530
transform 1 0 2524 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_4701
timestamp 1745462530
transform 1 0 2524 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_4702
timestamp 1745462530
transform 1 0 2516 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_4703
timestamp 1745462530
transform 1 0 2484 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_4704
timestamp 1745462530
transform 1 0 2444 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_4705
timestamp 1745462530
transform 1 0 2300 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_4706
timestamp 1745462530
transform 1 0 2284 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_4707
timestamp 1745462530
transform 1 0 3500 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_4708
timestamp 1745462530
transform 1 0 3492 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_4709
timestamp 1745462530
transform 1 0 3452 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_4710
timestamp 1745462530
transform 1 0 3396 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_4711
timestamp 1745462530
transform 1 0 3372 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_4712
timestamp 1745462530
transform 1 0 3236 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_4713
timestamp 1745462530
transform 1 0 3204 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_4714
timestamp 1745462530
transform 1 0 3148 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_4715
timestamp 1745462530
transform 1 0 3132 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_4716
timestamp 1745462530
transform 1 0 2060 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_4717
timestamp 1745462530
transform 1 0 3948 0 1 1315
box -2 -2 2 2
use M2_M1  M2_M1_4718
timestamp 1745462530
transform 1 0 3900 0 1 1315
box -2 -2 2 2
use M2_M1  M2_M1_4719
timestamp 1745462530
transform 1 0 3692 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_4720
timestamp 1745462530
transform 1 0 3564 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_4721
timestamp 1745462530
transform 1 0 3364 0 1 1315
box -2 -2 2 2
use M2_M1  M2_M1_4722
timestamp 1745462530
transform 1 0 3140 0 1 1315
box -2 -2 2 2
use M2_M1  M2_M1_4723
timestamp 1745462530
transform 1 0 3140 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_4724
timestamp 1745462530
transform 1 0 3028 0 1 1315
box -2 -2 2 2
use M2_M1  M2_M1_4725
timestamp 1745462530
transform 1 0 2756 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_4726
timestamp 1745462530
transform 1 0 2556 0 1 1315
box -2 -2 2 2
use M2_M1  M2_M1_4727
timestamp 1745462530
transform 1 0 2476 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_4728
timestamp 1745462530
transform 1 0 2348 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_4729
timestamp 1745462530
transform 1 0 2244 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_4730
timestamp 1745462530
transform 1 0 3100 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_4731
timestamp 1745462530
transform 1 0 3084 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_4732
timestamp 1745462530
transform 1 0 3052 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_4733
timestamp 1745462530
transform 1 0 2996 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_4734
timestamp 1745462530
transform 1 0 2956 0 1 2305
box -2 -2 2 2
use M2_M1  M2_M1_4735
timestamp 1745462530
transform 1 0 2924 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_4736
timestamp 1745462530
transform 1 0 2916 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_4737
timestamp 1745462530
transform 1 0 2764 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_4738
timestamp 1745462530
transform 1 0 2748 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_4739
timestamp 1745462530
transform 1 0 2684 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_4740
timestamp 1745462530
transform 1 0 2652 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_4741
timestamp 1745462530
transform 1 0 2564 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_4742
timestamp 1745462530
transform 1 0 2244 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_4743
timestamp 1745462530
transform 1 0 2084 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_4744
timestamp 1745462530
transform 1 0 2036 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_4745
timestamp 1745462530
transform 1 0 1948 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_4746
timestamp 1745462530
transform 1 0 1540 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_4747
timestamp 1745462530
transform 1 0 1380 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_4748
timestamp 1745462530
transform 1 0 1284 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_4749
timestamp 1745462530
transform 1 0 1180 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_4750
timestamp 1745462530
transform 1 0 1044 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_4751
timestamp 1745462530
transform 1 0 1020 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_4752
timestamp 1745462530
transform 1 0 1012 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_4753
timestamp 1745462530
transform 1 0 940 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_4754
timestamp 1745462530
transform 1 0 940 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_4755
timestamp 1745462530
transform 1 0 932 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_4756
timestamp 1745462530
transform 1 0 2132 0 1 1315
box -2 -2 2 2
use M2_M1  M2_M1_4757
timestamp 1745462530
transform 1 0 2108 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_4758
timestamp 1745462530
transform 1 0 1916 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_4759
timestamp 1745462530
transform 1 0 1740 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_4760
timestamp 1745462530
transform 1 0 1532 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_4761
timestamp 1745462530
transform 1 0 1276 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_4762
timestamp 1745462530
transform 1 0 1244 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_4763
timestamp 1745462530
transform 1 0 1180 0 1 1315
box -2 -2 2 2
use M2_M1  M2_M1_4764
timestamp 1745462530
transform 1 0 1132 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_4765
timestamp 1745462530
transform 1 0 1076 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_4766
timestamp 1745462530
transform 1 0 1044 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_4767
timestamp 1745462530
transform 1 0 972 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_4768
timestamp 1745462530
transform 1 0 964 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_4769
timestamp 1745462530
transform 1 0 508 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_4770
timestamp 1745462530
transform 1 0 348 0 1 3595
box -2 -2 2 2
use M2_M1  M2_M1_4771
timestamp 1745462530
transform 1 0 284 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_4772
timestamp 1745462530
transform 1 0 276 0 1 3595
box -2 -2 2 2
use M2_M1  M2_M1_4773
timestamp 1745462530
transform 1 0 252 0 1 3545
box -2 -2 2 2
use M2_M1  M2_M1_4774
timestamp 1745462530
transform 1 0 220 0 1 3545
box -2 -2 2 2
use M2_M1  M2_M1_4775
timestamp 1745462530
transform 1 0 460 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_4776
timestamp 1745462530
transform 1 0 420 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_4777
timestamp 1745462530
transform 1 0 356 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_4778
timestamp 1745462530
transform 1 0 332 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_4779
timestamp 1745462530
transform 1 0 324 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_4780
timestamp 1745462530
transform 1 0 348 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_4781
timestamp 1745462530
transform 1 0 332 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_4782
timestamp 1745462530
transform 1 0 308 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_4783
timestamp 1745462530
transform 1 0 284 0 1 3515
box -2 -2 2 2
use M2_M1  M2_M1_4784
timestamp 1745462530
transform 1 0 164 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_4785
timestamp 1745462530
transform 1 0 412 0 1 3515
box -2 -2 2 2
use M2_M1  M2_M1_4786
timestamp 1745462530
transform 1 0 356 0 1 3515
box -2 -2 2 2
use M2_M1  M2_M1_4787
timestamp 1745462530
transform 1 0 276 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_4788
timestamp 1745462530
transform 1 0 276 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_4789
timestamp 1745462530
transform 1 0 236 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_4790
timestamp 1745462530
transform 1 0 188 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_4791
timestamp 1745462530
transform 1 0 180 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_4792
timestamp 1745462530
transform 1 0 116 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_4793
timestamp 1745462530
transform 1 0 348 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_4794
timestamp 1745462530
transform 1 0 316 0 1 3625
box -2 -2 2 2
use M2_M1  M2_M1_4795
timestamp 1745462530
transform 1 0 276 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_4796
timestamp 1745462530
transform 1 0 212 0 1 3625
box -2 -2 2 2
use M2_M1  M2_M1_4797
timestamp 1745462530
transform 1 0 212 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_4798
timestamp 1745462530
transform 1 0 212 0 1 3425
box -2 -2 2 2
use M2_M1  M2_M1_4799
timestamp 1745462530
transform 1 0 268 0 1 3515
box -2 -2 2 2
use M2_M1  M2_M1_4800
timestamp 1745462530
transform 1 0 268 0 1 3425
box -2 -2 2 2
use M2_M1  M2_M1_4801
timestamp 1745462530
transform 1 0 428 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_4802
timestamp 1745462530
transform 1 0 348 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_4803
timestamp 1745462530
transform 1 0 316 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_4804
timestamp 1745462530
transform 1 0 308 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_4805
timestamp 1745462530
transform 1 0 212 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_4806
timestamp 1745462530
transform 1 0 180 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_4807
timestamp 1745462530
transform 1 0 212 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_4808
timestamp 1745462530
transform 1 0 140 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_4809
timestamp 1745462530
transform 1 0 124 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_4810
timestamp 1745462530
transform 1 0 116 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_4811
timestamp 1745462530
transform 1 0 268 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_4812
timestamp 1745462530
transform 1 0 196 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_4813
timestamp 1745462530
transform 1 0 2972 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_4814
timestamp 1745462530
transform 1 0 2956 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_4815
timestamp 1745462530
transform 1 0 2924 0 1 2645
box -2 -2 2 2
use M2_M1  M2_M1_4816
timestamp 1745462530
transform 1 0 2924 0 1 2625
box -2 -2 2 2
use M2_M1  M2_M1_4817
timestamp 1745462530
transform 1 0 2924 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_4818
timestamp 1745462530
transform 1 0 2764 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_4819
timestamp 1745462530
transform 1 0 2724 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_4820
timestamp 1745462530
transform 1 0 2700 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_4821
timestamp 1745462530
transform 1 0 2908 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_4822
timestamp 1745462530
transform 1 0 2884 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_4823
timestamp 1745462530
transform 1 0 2884 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_4824
timestamp 1745462530
transform 1 0 3140 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4825
timestamp 1745462530
transform 1 0 3076 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_4826
timestamp 1745462530
transform 1 0 3028 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_4827
timestamp 1745462530
transform 1 0 2868 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_4828
timestamp 1745462530
transform 1 0 2820 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4829
timestamp 1745462530
transform 1 0 2820 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4830
timestamp 1745462530
transform 1 0 3044 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4831
timestamp 1745462530
transform 1 0 3020 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_4832
timestamp 1745462530
transform 1 0 2916 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4833
timestamp 1745462530
transform 1 0 4164 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_4834
timestamp 1745462530
transform 1 0 4132 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_4835
timestamp 1745462530
transform 1 0 4076 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4836
timestamp 1745462530
transform 1 0 4044 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4837
timestamp 1745462530
transform 1 0 3156 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4838
timestamp 1745462530
transform 1 0 3140 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_4839
timestamp 1745462530
transform 1 0 3124 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4840
timestamp 1745462530
transform 1 0 4204 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_4841
timestamp 1745462530
transform 1 0 4092 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_4842
timestamp 1745462530
transform 1 0 4052 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4843
timestamp 1745462530
transform 1 0 4052 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_4844
timestamp 1745462530
transform 1 0 3900 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_4845
timestamp 1745462530
transform 1 0 3820 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_4846
timestamp 1745462530
transform 1 0 3820 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4847
timestamp 1745462530
transform 1 0 3700 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4848
timestamp 1745462530
transform 1 0 3316 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4849
timestamp 1745462530
transform 1 0 3284 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_4850
timestamp 1745462530
transform 1 0 2948 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_4851
timestamp 1745462530
transform 1 0 3548 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_4852
timestamp 1745462530
transform 1 0 3532 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4853
timestamp 1745462530
transform 1 0 3500 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_4854
timestamp 1745462530
transform 1 0 3468 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4855
timestamp 1745462530
transform 1 0 4372 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_4856
timestamp 1745462530
transform 1 0 4260 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_4857
timestamp 1745462530
transform 1 0 4100 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_4858
timestamp 1745462530
transform 1 0 3212 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_4859
timestamp 1745462530
transform 1 0 3172 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_4860
timestamp 1745462530
transform 1 0 3172 0 1 2045
box -2 -2 2 2
use M2_M1  M2_M1_4861
timestamp 1745462530
transform 1 0 4244 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_4862
timestamp 1745462530
transform 1 0 4132 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_4863
timestamp 1745462530
transform 1 0 4092 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_4864
timestamp 1745462530
transform 1 0 4060 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_4865
timestamp 1745462530
transform 1 0 3892 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_4866
timestamp 1745462530
transform 1 0 3804 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_4867
timestamp 1745462530
transform 1 0 3500 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_4868
timestamp 1745462530
transform 1 0 3316 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_4869
timestamp 1745462530
transform 1 0 3284 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_4870
timestamp 1745462530
transform 1 0 3748 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_4871
timestamp 1745462530
transform 1 0 3572 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_4872
timestamp 1745462530
transform 1 0 3540 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_4873
timestamp 1745462530
transform 1 0 4372 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4874
timestamp 1745462530
transform 1 0 4244 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4875
timestamp 1745462530
transform 1 0 4116 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4876
timestamp 1745462530
transform 1 0 3356 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4877
timestamp 1745462530
transform 1 0 3252 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_4878
timestamp 1745462530
transform 1 0 3212 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4879
timestamp 1745462530
transform 1 0 4356 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4880
timestamp 1745462530
transform 1 0 4188 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_4881
timestamp 1745462530
transform 1 0 4076 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_4882
timestamp 1745462530
transform 1 0 3972 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4883
timestamp 1745462530
transform 1 0 3796 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4884
timestamp 1745462530
transform 1 0 3764 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4885
timestamp 1745462530
transform 1 0 3468 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4886
timestamp 1745462530
transform 1 0 3436 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_4887
timestamp 1745462530
transform 1 0 3412 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_4888
timestamp 1745462530
transform 1 0 3796 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4889
timestamp 1745462530
transform 1 0 3612 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_4890
timestamp 1745462530
transform 1 0 3604 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4891
timestamp 1745462530
transform 1 0 4332 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_4892
timestamp 1745462530
transform 1 0 4204 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_4893
timestamp 1745462530
transform 1 0 4148 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_4894
timestamp 1745462530
transform 1 0 4076 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_4895
timestamp 1745462530
transform 1 0 3244 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_4896
timestamp 1745462530
transform 1 0 3164 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_4897
timestamp 1745462530
transform 1 0 3036 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_4898
timestamp 1745462530
transform 1 0 4372 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_4899
timestamp 1745462530
transform 1 0 4260 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_4900
timestamp 1745462530
transform 1 0 4124 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_4901
timestamp 1745462530
transform 1 0 4076 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_4902
timestamp 1745462530
transform 1 0 3876 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_4903
timestamp 1745462530
transform 1 0 3844 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_4904
timestamp 1745462530
transform 1 0 3820 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_4905
timestamp 1745462530
transform 1 0 3764 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_4906
timestamp 1745462530
transform 1 0 3444 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_4907
timestamp 1745462530
transform 1 0 3348 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_4908
timestamp 1745462530
transform 1 0 3348 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_4909
timestamp 1745462530
transform 1 0 3324 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_4910
timestamp 1745462530
transform 1 0 3684 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_4911
timestamp 1745462530
transform 1 0 3588 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_4912
timestamp 1745462530
transform 1 0 3588 0 1 2385
box -2 -2 2 2
use M2_M1  M2_M1_4913
timestamp 1745462530
transform 1 0 3588 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_4914
timestamp 1745462530
transform 1 0 3564 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_4915
timestamp 1745462530
transform 1 0 3564 0 1 2385
box -2 -2 2 2
use M2_M1  M2_M1_4916
timestamp 1745462530
transform 1 0 4268 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_4917
timestamp 1745462530
transform 1 0 4084 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_4918
timestamp 1745462530
transform 1 0 4044 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_4919
timestamp 1745462530
transform 1 0 3148 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_4920
timestamp 1745462530
transform 1 0 3004 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_4921
timestamp 1745462530
transform 1 0 4372 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_4922
timestamp 1745462530
transform 1 0 4116 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_4923
timestamp 1745462530
transform 1 0 4028 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_4924
timestamp 1745462530
transform 1 0 3988 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_4925
timestamp 1745462530
transform 1 0 3820 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_4926
timestamp 1745462530
transform 1 0 3788 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_4927
timestamp 1745462530
transform 1 0 3452 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_4928
timestamp 1745462530
transform 1 0 3356 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_4929
timestamp 1745462530
transform 1 0 3316 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_4930
timestamp 1745462530
transform 1 0 3772 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_4931
timestamp 1745462530
transform 1 0 3580 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_4932
timestamp 1745462530
transform 1 0 3548 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_4933
timestamp 1745462530
transform 1 0 4076 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_4934
timestamp 1745462530
transform 1 0 3980 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_4935
timestamp 1745462530
transform 1 0 3980 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4936
timestamp 1745462530
transform 1 0 3956 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_4937
timestamp 1745462530
transform 1 0 3124 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4938
timestamp 1745462530
transform 1 0 3068 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4939
timestamp 1745462530
transform 1 0 2972 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_4940
timestamp 1745462530
transform 1 0 4044 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_4941
timestamp 1745462530
transform 1 0 4012 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4942
timestamp 1745462530
transform 1 0 3988 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_4943
timestamp 1745462530
transform 1 0 3932 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_4944
timestamp 1745462530
transform 1 0 3772 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4945
timestamp 1745462530
transform 1 0 3732 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_4946
timestamp 1745462530
transform 1 0 3732 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_4947
timestamp 1745462530
transform 1 0 3652 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4948
timestamp 1745462530
transform 1 0 3404 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_4949
timestamp 1745462530
transform 1 0 3332 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_4950
timestamp 1745462530
transform 1 0 3268 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_4951
timestamp 1745462530
transform 1 0 3260 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_4952
timestamp 1745462530
transform 1 0 3652 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_4953
timestamp 1745462530
transform 1 0 3604 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4954
timestamp 1745462530
transform 1 0 3500 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4955
timestamp 1745462530
transform 1 0 4340 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_4956
timestamp 1745462530
transform 1 0 4156 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_4957
timestamp 1745462530
transform 1 0 3932 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_4958
timestamp 1745462530
transform 1 0 3252 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_4959
timestamp 1745462530
transform 1 0 3172 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_4960
timestamp 1745462530
transform 1 0 3092 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4961
timestamp 1745462530
transform 1 0 4340 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4962
timestamp 1745462530
transform 1 0 4172 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_4963
timestamp 1745462530
transform 1 0 3980 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4964
timestamp 1745462530
transform 1 0 3956 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4965
timestamp 1745462530
transform 1 0 3812 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_4966
timestamp 1745462530
transform 1 0 3740 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4967
timestamp 1745462530
transform 1 0 3540 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_4968
timestamp 1745462530
transform 1 0 3484 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_4969
timestamp 1745462530
transform 1 0 3372 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_4970
timestamp 1745462530
transform 1 0 3716 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4971
timestamp 1745462530
transform 1 0 3628 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_4972
timestamp 1745462530
transform 1 0 3572 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4973
timestamp 1745462530
transform 1 0 3092 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_4974
timestamp 1745462530
transform 1 0 3036 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_4975
timestamp 1745462530
transform 1 0 3020 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_4976
timestamp 1745462530
transform 1 0 2980 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_4977
timestamp 1745462530
transform 1 0 2948 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_4978
timestamp 1745462530
transform 1 0 2900 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_4979
timestamp 1745462530
transform 1 0 2828 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_4980
timestamp 1745462530
transform 1 0 2820 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_4981
timestamp 1745462530
transform 1 0 2884 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_4982
timestamp 1745462530
transform 1 0 2716 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_4983
timestamp 1745462530
transform 1 0 2636 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_4984
timestamp 1745462530
transform 1 0 2604 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_4985
timestamp 1745462530
transform 1 0 3012 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_4986
timestamp 1745462530
transform 1 0 2636 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_4987
timestamp 1745462530
transform 1 0 2636 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_4988
timestamp 1745462530
transform 1 0 2988 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_4989
timestamp 1745462530
transform 1 0 2572 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_4990
timestamp 1745462530
transform 1 0 2540 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_4991
timestamp 1745462530
transform 1 0 3028 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_4992
timestamp 1745462530
transform 1 0 2716 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_4993
timestamp 1745462530
transform 1 0 2716 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_4994
timestamp 1745462530
transform 1 0 2684 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_4995
timestamp 1745462530
transform 1 0 3940 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_4996
timestamp 1745462530
transform 1 0 3276 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_4997
timestamp 1745462530
transform 1 0 3172 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_4998
timestamp 1745462530
transform 1 0 2988 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_4999
timestamp 1745462530
transform 1 0 3148 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_5000
timestamp 1745462530
transform 1 0 2908 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_5001
timestamp 1745462530
transform 1 0 2868 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_5002
timestamp 1745462530
transform 1 0 2820 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_5003
timestamp 1745462530
transform 1 0 3052 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_5004
timestamp 1745462530
transform 1 0 2932 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5005
timestamp 1745462530
transform 1 0 2924 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_5006
timestamp 1745462530
transform 1 0 2852 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_5007
timestamp 1745462530
transform 1 0 3236 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_5008
timestamp 1745462530
transform 1 0 3148 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_5009
timestamp 1745462530
transform 1 0 3028 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_5010
timestamp 1745462530
transform 1 0 2980 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_5011
timestamp 1745462530
transform 1 0 3060 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5012
timestamp 1745462530
transform 1 0 2908 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5013
timestamp 1745462530
transform 1 0 2772 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5014
timestamp 1745462530
transform 1 0 2756 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5015
timestamp 1745462530
transform 1 0 3244 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5016
timestamp 1745462530
transform 1 0 2988 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5017
timestamp 1745462530
transform 1 0 2900 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5018
timestamp 1745462530
transform 1 0 2900 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5019
timestamp 1745462530
transform 1 0 4036 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5020
timestamp 1745462530
transform 1 0 3924 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5021
timestamp 1745462530
transform 1 0 3892 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_5022
timestamp 1745462530
transform 1 0 3852 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_5023
timestamp 1745462530
transform 1 0 3340 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_5024
timestamp 1745462530
transform 1 0 3236 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_5025
timestamp 1745462530
transform 1 0 3116 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_5026
timestamp 1745462530
transform 1 0 3388 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5027
timestamp 1745462530
transform 1 0 3388 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_5028
timestamp 1745462530
transform 1 0 3372 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_5029
timestamp 1745462530
transform 1 0 3332 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_5030
timestamp 1745462530
transform 1 0 3196 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_5031
timestamp 1745462530
transform 1 0 4044 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_5032
timestamp 1745462530
transform 1 0 3916 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_5033
timestamp 1745462530
transform 1 0 3828 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_5034
timestamp 1745462530
transform 1 0 3708 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_5035
timestamp 1745462530
transform 1 0 3532 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5036
timestamp 1745462530
transform 1 0 3468 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_5037
timestamp 1745462530
transform 1 0 3324 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_5038
timestamp 1745462530
transform 1 0 3300 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5039
timestamp 1745462530
transform 1 0 3724 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5040
timestamp 1745462530
transform 1 0 3588 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_5041
timestamp 1745462530
transform 1 0 3532 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_5042
timestamp 1745462530
transform 1 0 3356 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5043
timestamp 1745462530
transform 1 0 4276 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_5044
timestamp 1745462530
transform 1 0 4180 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5045
timestamp 1745462530
transform 1 0 3996 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5046
timestamp 1745462530
transform 1 0 3820 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_5047
timestamp 1745462530
transform 1 0 4292 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_5048
timestamp 1745462530
transform 1 0 4132 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_5049
timestamp 1745462530
transform 1 0 3188 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_5050
timestamp 1745462530
transform 1 0 3156 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_5051
timestamp 1745462530
transform 1 0 4372 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_5052
timestamp 1745462530
transform 1 0 4356 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_5053
timestamp 1745462530
transform 1 0 3316 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_5054
timestamp 1745462530
transform 1 0 3220 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_5055
timestamp 1745462530
transform 1 0 4068 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_5056
timestamp 1745462530
transform 1 0 3916 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_5057
timestamp 1745462530
transform 1 0 3796 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_5058
timestamp 1745462530
transform 1 0 3708 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_5059
timestamp 1745462530
transform 1 0 4180 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_5060
timestamp 1745462530
transform 1 0 4100 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5061
timestamp 1745462530
transform 1 0 3444 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5062
timestamp 1745462530
transform 1 0 3436 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_5063
timestamp 1745462530
transform 1 0 4372 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_5064
timestamp 1745462530
transform 1 0 4324 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5065
timestamp 1745462530
transform 1 0 3540 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_5066
timestamp 1745462530
transform 1 0 3396 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5067
timestamp 1745462530
transform 1 0 4092 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5068
timestamp 1745462530
transform 1 0 3996 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5069
timestamp 1745462530
transform 1 0 3900 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5070
timestamp 1745462530
transform 1 0 3540 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_5071
timestamp 1745462530
transform 1 0 3412 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_5072
timestamp 1745462530
transform 1 0 3156 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_5073
timestamp 1745462530
transform 1 0 3684 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_5074
timestamp 1745462530
transform 1 0 3604 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_5075
timestamp 1745462530
transform 1 0 3604 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_5076
timestamp 1745462530
transform 1 0 3244 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_5077
timestamp 1745462530
transform 1 0 3956 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_5078
timestamp 1745462530
transform 1 0 3844 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_5079
timestamp 1745462530
transform 1 0 3748 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_5080
timestamp 1745462530
transform 1 0 3700 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_5081
timestamp 1745462530
transform 1 0 3636 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5082
timestamp 1745462530
transform 1 0 3348 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5083
timestamp 1745462530
transform 1 0 3796 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_5084
timestamp 1745462530
transform 1 0 3732 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5085
timestamp 1745462530
transform 1 0 3428 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5086
timestamp 1745462530
transform 1 0 4372 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5087
timestamp 1745462530
transform 1 0 4260 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_5088
timestamp 1745462530
transform 1 0 4196 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_5089
timestamp 1745462530
transform 1 0 4028 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_5090
timestamp 1745462530
transform 1 0 4372 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_5091
timestamp 1745462530
transform 1 0 4268 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_5092
timestamp 1745462530
transform 1 0 4364 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_5093
timestamp 1745462530
transform 1 0 4252 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_5094
timestamp 1745462530
transform 1 0 4156 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_5095
timestamp 1745462530
transform 1 0 4092 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5096
timestamp 1745462530
transform 1 0 4380 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_5097
timestamp 1745462530
transform 1 0 4268 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5098
timestamp 1745462530
transform 1 0 4052 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_5099
timestamp 1745462530
transform 1 0 3924 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_5100
timestamp 1745462530
transform 1 0 3908 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5101
timestamp 1745462530
transform 1 0 3588 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_5102
timestamp 1745462530
transform 1 0 3460 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_5103
timestamp 1745462530
transform 1 0 3084 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_5104
timestamp 1745462530
transform 1 0 3716 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_5105
timestamp 1745462530
transform 1 0 3636 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_5106
timestamp 1745462530
transform 1 0 3620 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_5107
timestamp 1745462530
transform 1 0 2988 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_5108
timestamp 1745462530
transform 1 0 3844 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_5109
timestamp 1745462530
transform 1 0 3836 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_5110
timestamp 1745462530
transform 1 0 3172 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_5111
timestamp 1745462530
transform 1 0 3444 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_5112
timestamp 1745462530
transform 1 0 3428 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5113
timestamp 1745462530
transform 1 0 3028 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5114
timestamp 1745462530
transform 1 0 3636 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_5115
timestamp 1745462530
transform 1 0 3196 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5116
timestamp 1745462530
transform 1 0 4156 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_5117
timestamp 1745462530
transform 1 0 4044 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_5118
timestamp 1745462530
transform 1 0 4364 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_5119
timestamp 1745462530
transform 1 0 4252 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_5120
timestamp 1745462530
transform 1 0 4268 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_5121
timestamp 1745462530
transform 1 0 4172 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_5122
timestamp 1745462530
transform 1 0 4028 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_5123
timestamp 1745462530
transform 1 0 3940 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_5124
timestamp 1745462530
transform 1 0 4364 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_5125
timestamp 1745462530
transform 1 0 4260 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_5126
timestamp 1745462530
transform 1 0 4172 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_5127
timestamp 1745462530
transform 1 0 3844 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_5128
timestamp 1745462530
transform 1 0 3844 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_5129
timestamp 1745462530
transform 1 0 3844 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_5130
timestamp 1745462530
transform 1 0 3348 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_5131
timestamp 1745462530
transform 1 0 3316 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_5132
timestamp 1745462530
transform 1 0 3100 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_5133
timestamp 1745462530
transform 1 0 4076 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_5134
timestamp 1745462530
transform 1 0 3964 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_5135
timestamp 1745462530
transform 1 0 3924 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_5136
timestamp 1745462530
transform 1 0 3924 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_5137
timestamp 1745462530
transform 1 0 3788 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_5138
timestamp 1745462530
transform 1 0 3740 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_5139
timestamp 1745462530
transform 1 0 3700 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_5140
timestamp 1745462530
transform 1 0 3668 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_5141
timestamp 1745462530
transform 1 0 3564 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_5142
timestamp 1745462530
transform 1 0 3564 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_5143
timestamp 1745462530
transform 1 0 3412 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_5144
timestamp 1745462530
transform 1 0 3412 0 1 1185
box -2 -2 2 2
use M2_M1  M2_M1_5145
timestamp 1745462530
transform 1 0 3340 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_5146
timestamp 1745462530
transform 1 0 3676 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_5147
timestamp 1745462530
transform 1 0 3660 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_5148
timestamp 1745462530
transform 1 0 3572 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_5149
timestamp 1745462530
transform 1 0 3540 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_5150
timestamp 1745462530
transform 1 0 4268 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_5151
timestamp 1745462530
transform 1 0 4092 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_5152
timestamp 1745462530
transform 1 0 3964 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_5153
timestamp 1745462530
transform 1 0 3812 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_5154
timestamp 1745462530
transform 1 0 3340 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_5155
timestamp 1745462530
transform 1 0 3316 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_5156
timestamp 1745462530
transform 1 0 3276 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_5157
timestamp 1745462530
transform 1 0 3172 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_5158
timestamp 1745462530
transform 1 0 3140 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_5159
timestamp 1745462530
transform 1 0 3140 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_5160
timestamp 1745462530
transform 1 0 4372 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_5161
timestamp 1745462530
transform 1 0 4260 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_5162
timestamp 1745462530
transform 1 0 4012 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_5163
timestamp 1745462530
transform 1 0 3868 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_5164
timestamp 1745462530
transform 1 0 3836 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_5165
timestamp 1745462530
transform 1 0 3748 0 1 995
box -2 -2 2 2
use M2_M1  M2_M1_5166
timestamp 1745462530
transform 1 0 3676 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_5167
timestamp 1745462530
transform 1 0 3668 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_5168
timestamp 1745462530
transform 1 0 3516 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_5169
timestamp 1745462530
transform 1 0 3516 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_5170
timestamp 1745462530
transform 1 0 3500 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_5171
timestamp 1745462530
transform 1 0 3340 0 1 1115
box -2 -2 2 2
use M2_M1  M2_M1_5172
timestamp 1745462530
transform 1 0 4180 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_5173
timestamp 1745462530
transform 1 0 4124 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_5174
timestamp 1745462530
transform 1 0 3612 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_5175
timestamp 1745462530
transform 1 0 3604 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_5176
timestamp 1745462530
transform 1 0 4364 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_5177
timestamp 1745462530
transform 1 0 4364 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_5178
timestamp 1745462530
transform 1 0 3980 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_5179
timestamp 1745462530
transform 1 0 4068 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_5180
timestamp 1745462530
transform 1 0 3988 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_5181
timestamp 1745462530
transform 1 0 3356 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_5182
timestamp 1745462530
transform 1 0 3188 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_5183
timestamp 1745462530
transform 1 0 4372 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_5184
timestamp 1745462530
transform 1 0 4180 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_5185
timestamp 1745462530
transform 1 0 4036 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_5186
timestamp 1745462530
transform 1 0 3980 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_5187
timestamp 1745462530
transform 1 0 4212 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_5188
timestamp 1745462530
transform 1 0 4092 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_5189
timestamp 1745462530
transform 1 0 3900 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_5190
timestamp 1745462530
transform 1 0 3804 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_5191
timestamp 1745462530
transform 1 0 3940 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_5192
timestamp 1745462530
transform 1 0 3916 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_5193
timestamp 1745462530
transform 1 0 3516 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_5194
timestamp 1745462530
transform 1 0 3364 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_5195
timestamp 1745462530
transform 1 0 4372 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_5196
timestamp 1745462530
transform 1 0 4188 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_5197
timestamp 1745462530
transform 1 0 3692 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_5198
timestamp 1745462530
transform 1 0 4244 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_5199
timestamp 1745462530
transform 1 0 4116 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_5200
timestamp 1745462530
transform 1 0 3948 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_5201
timestamp 1745462530
transform 1 0 3916 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_5202
timestamp 1745462530
transform 1 0 4284 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_5203
timestamp 1745462530
transform 1 0 4076 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_5204
timestamp 1745462530
transform 1 0 3324 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_5205
timestamp 1745462530
transform 1 0 3276 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_5206
timestamp 1745462530
transform 1 0 4364 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_5207
timestamp 1745462530
transform 1 0 4364 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_5208
timestamp 1745462530
transform 1 0 4036 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_5209
timestamp 1745462530
transform 1 0 3916 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_5210
timestamp 1745462530
transform 1 0 4372 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_5211
timestamp 1745462530
transform 1 0 4260 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_5212
timestamp 1745462530
transform 1 0 3844 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_5213
timestamp 1745462530
transform 1 0 3748 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_5214
timestamp 1745462530
transform 1 0 4036 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_5215
timestamp 1745462530
transform 1 0 3476 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_5216
timestamp 1745462530
transform 1 0 3380 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_5217
timestamp 1745462530
transform 1 0 4372 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_5218
timestamp 1745462530
transform 1 0 4228 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_5219
timestamp 1745462530
transform 1 0 3612 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_5220
timestamp 1745462530
transform 1 0 3612 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_5221
timestamp 1745462530
transform 1 0 4116 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_5222
timestamp 1745462530
transform 1 0 4036 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_5223
timestamp 1745462530
transform 1 0 4028 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_5224
timestamp 1745462530
transform 1 0 3428 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_5225
timestamp 1745462530
transform 1 0 3324 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_5226
timestamp 1745462530
transform 1 0 3228 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_5227
timestamp 1745462530
transform 1 0 4132 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_5228
timestamp 1745462530
transform 1 0 4076 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_5229
timestamp 1745462530
transform 1 0 3972 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_5230
timestamp 1745462530
transform 1 0 3924 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_5231
timestamp 1745462530
transform 1 0 3836 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_5232
timestamp 1745462530
transform 1 0 3804 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_5233
timestamp 1745462530
transform 1 0 3548 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_5234
timestamp 1745462530
transform 1 0 3396 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_5235
timestamp 1745462530
transform 1 0 3724 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_5236
timestamp 1745462530
transform 1 0 3684 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_5237
timestamp 1745462530
transform 1 0 3684 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_5238
timestamp 1745462530
transform 1 0 4220 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_5239
timestamp 1745462530
transform 1 0 4108 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_5240
timestamp 1745462530
transform 1 0 4196 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_5241
timestamp 1745462530
transform 1 0 4092 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_5242
timestamp 1745462530
transform 1 0 4356 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_5243
timestamp 1745462530
transform 1 0 4244 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_5244
timestamp 1745462530
transform 1 0 4372 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_5245
timestamp 1745462530
transform 1 0 4260 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_5246
timestamp 1745462530
transform 1 0 4084 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_5247
timestamp 1745462530
transform 1 0 3964 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_5248
timestamp 1745462530
transform 1 0 3764 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_5249
timestamp 1745462530
transform 1 0 3708 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_5250
timestamp 1745462530
transform 1 0 3996 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_5251
timestamp 1745462530
transform 1 0 3940 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_5252
timestamp 1745462530
transform 1 0 3932 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_5253
timestamp 1745462530
transform 1 0 3196 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_5254
timestamp 1745462530
transform 1 0 3180 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_5255
timestamp 1745462530
transform 1 0 3084 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_5256
timestamp 1745462530
transform 1 0 3972 0 1 1095
box -2 -2 2 2
use M2_M1  M2_M1_5257
timestamp 1745462530
transform 1 0 3884 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_5258
timestamp 1745462530
transform 1 0 3828 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_5259
timestamp 1745462530
transform 1 0 3772 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_5260
timestamp 1745462530
transform 1 0 3652 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_5261
timestamp 1745462530
transform 1 0 3644 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_5262
timestamp 1745462530
transform 1 0 3492 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_5263
timestamp 1745462530
transform 1 0 3412 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_5264
timestamp 1745462530
transform 1 0 3276 0 1 1105
box -2 -2 2 2
use M2_M1  M2_M1_5265
timestamp 1745462530
transform 1 0 3652 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_5266
timestamp 1745462530
transform 1 0 3604 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_5267
timestamp 1745462530
transform 1 0 3564 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_5268
timestamp 1745462530
transform 1 0 3428 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_5269
timestamp 1745462530
transform 1 0 3380 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_5270
timestamp 1745462530
transform 1 0 3540 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_5271
timestamp 1745462530
transform 1 0 3492 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_5272
timestamp 1745462530
transform 1 0 3316 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_5273
timestamp 1745462530
transform 1 0 3268 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_5274
timestamp 1745462530
transform 1 0 3084 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_5275
timestamp 1745462530
transform 1 0 2972 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_5276
timestamp 1745462530
transform 1 0 2972 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_5277
timestamp 1745462530
transform 1 0 2860 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_5278
timestamp 1745462530
transform 1 0 3028 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_5279
timestamp 1745462530
transform 1 0 3004 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_5280
timestamp 1745462530
transform 1 0 3004 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_5281
timestamp 1745462530
transform 1 0 2892 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_5282
timestamp 1745462530
transform 1 0 2468 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_5283
timestamp 1745462530
transform 1 0 2324 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_5284
timestamp 1745462530
transform 1 0 2324 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_5285
timestamp 1745462530
transform 1 0 2652 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_5286
timestamp 1745462530
transform 1 0 2556 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_5287
timestamp 1745462530
transform 1 0 2548 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_5288
timestamp 1745462530
transform 1 0 2516 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_5289
timestamp 1745462530
transform 1 0 2532 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_5290
timestamp 1745462530
transform 1 0 2452 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_5291
timestamp 1745462530
transform 1 0 2444 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_5292
timestamp 1745462530
transform 1 0 2812 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_5293
timestamp 1745462530
transform 1 0 2756 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_5294
timestamp 1745462530
transform 1 0 2708 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_5295
timestamp 1745462530
transform 1 0 2692 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_5296
timestamp 1745462530
transform 1 0 3164 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_5297
timestamp 1745462530
transform 1 0 3084 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_5298
timestamp 1745462530
transform 1 0 2908 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_5299
timestamp 1745462530
transform 1 0 2892 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_5300
timestamp 1745462530
transform 1 0 3100 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_5301
timestamp 1745462530
transform 1 0 2972 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_5302
timestamp 1745462530
transform 1 0 2868 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_5303
timestamp 1745462530
transform 1 0 2428 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_5304
timestamp 1745462530
transform 1 0 2268 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_5305
timestamp 1745462530
transform 1 0 2244 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_5306
timestamp 1745462530
transform 1 0 2244 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_5307
timestamp 1745462530
transform 1 0 2676 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_5308
timestamp 1745462530
transform 1 0 2564 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_5309
timestamp 1745462530
transform 1 0 2532 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_5310
timestamp 1745462530
transform 1 0 2524 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_5311
timestamp 1745462530
transform 1 0 2484 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_5312
timestamp 1745462530
transform 1 0 2412 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_5313
timestamp 1745462530
transform 1 0 2412 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_5314
timestamp 1745462530
transform 1 0 2412 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_5315
timestamp 1745462530
transform 1 0 2788 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_5316
timestamp 1745462530
transform 1 0 2780 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_5317
timestamp 1745462530
transform 1 0 2716 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_5318
timestamp 1745462530
transform 1 0 3100 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_5319
timestamp 1745462530
transform 1 0 3036 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_5320
timestamp 1745462530
transform 1 0 3036 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_5321
timestamp 1745462530
transform 1 0 3012 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_5322
timestamp 1745462530
transform 1 0 2956 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_5323
timestamp 1745462530
transform 1 0 3076 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_5324
timestamp 1745462530
transform 1 0 2988 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_5325
timestamp 1745462530
transform 1 0 2884 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_5326
timestamp 1745462530
transform 1 0 2500 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_5327
timestamp 1745462530
transform 1 0 2404 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_5328
timestamp 1745462530
transform 1 0 2316 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_5329
timestamp 1745462530
transform 1 0 2276 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_5330
timestamp 1745462530
transform 1 0 2532 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_5331
timestamp 1745462530
transform 1 0 2388 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_5332
timestamp 1745462530
transform 1 0 2300 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_5333
timestamp 1745462530
transform 1 0 2244 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_5334
timestamp 1745462530
transform 1 0 2692 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_5335
timestamp 1745462530
transform 1 0 2668 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_5336
timestamp 1745462530
transform 1 0 2516 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_5337
timestamp 1745462530
transform 1 0 2428 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_5338
timestamp 1745462530
transform 1 0 2868 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_5339
timestamp 1745462530
transform 1 0 2772 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_5340
timestamp 1745462530
transform 1 0 2764 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_5341
timestamp 1745462530
transform 1 0 2756 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_5342
timestamp 1745462530
transform 1 0 3204 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_5343
timestamp 1745462530
transform 1 0 3156 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_5344
timestamp 1745462530
transform 1 0 3116 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_5345
timestamp 1745462530
transform 1 0 3060 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_5346
timestamp 1745462530
transform 1 0 3116 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_5347
timestamp 1745462530
transform 1 0 3044 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_5348
timestamp 1745462530
transform 1 0 3012 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_5349
timestamp 1745462530
transform 1 0 2996 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_5350
timestamp 1745462530
transform 1 0 2468 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_5351
timestamp 1745462530
transform 1 0 2444 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_5352
timestamp 1745462530
transform 1 0 2244 0 1 795
box -2 -2 2 2
use M2_M1  M2_M1_5353
timestamp 1745462530
transform 1 0 2556 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_5354
timestamp 1745462530
transform 1 0 2540 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_5355
timestamp 1745462530
transform 1 0 2508 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_5356
timestamp 1745462530
transform 1 0 2500 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_5357
timestamp 1745462530
transform 1 0 2676 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_5358
timestamp 1745462530
transform 1 0 2628 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_5359
timestamp 1745462530
transform 1 0 2580 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_5360
timestamp 1745462530
transform 1 0 2452 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_5361
timestamp 1745462530
transform 1 0 3092 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_5362
timestamp 1745462530
transform 1 0 2980 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_5363
timestamp 1745462530
transform 1 0 2828 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_5364
timestamp 1745462530
transform 1 0 2780 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_5365
timestamp 1745462530
transform 1 0 3084 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_5366
timestamp 1745462530
transform 1 0 3068 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_5367
timestamp 1745462530
transform 1 0 2972 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_5368
timestamp 1745462530
transform 1 0 3156 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_5369
timestamp 1745462530
transform 1 0 3148 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_5370
timestamp 1745462530
transform 1 0 3044 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_5371
timestamp 1745462530
transform 1 0 2380 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_5372
timestamp 1745462530
transform 1 0 2196 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_5373
timestamp 1745462530
transform 1 0 2436 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_5374
timestamp 1745462530
transform 1 0 2420 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_5375
timestamp 1745462530
transform 1 0 2356 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_5376
timestamp 1745462530
transform 1 0 2460 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_5377
timestamp 1745462530
transform 1 0 2340 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_5378
timestamp 1745462530
transform 1 0 2212 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_5379
timestamp 1745462530
transform 1 0 2836 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_5380
timestamp 1745462530
transform 1 0 2804 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_5381
timestamp 1745462530
transform 1 0 2748 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_5382
timestamp 1745462530
transform 1 0 2876 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_5383
timestamp 1745462530
transform 1 0 2860 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_5384
timestamp 1745462530
transform 1 0 3196 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_5385
timestamp 1745462530
transform 1 0 3108 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_5386
timestamp 1745462530
transform 1 0 3068 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_5387
timestamp 1745462530
transform 1 0 3228 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_5388
timestamp 1745462530
transform 1 0 3116 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_5389
timestamp 1745462530
transform 1 0 3068 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_5390
timestamp 1745462530
transform 1 0 2196 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_5391
timestamp 1745462530
transform 1 0 2164 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_5392
timestamp 1745462530
transform 1 0 2492 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_5393
timestamp 1745462530
transform 1 0 2428 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_5394
timestamp 1745462530
transform 1 0 2356 0 1 985
box -2 -2 2 2
use M2_M1  M2_M1_5395
timestamp 1745462530
transform 1 0 2244 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_5396
timestamp 1745462530
transform 1 0 2180 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_5397
timestamp 1745462530
transform 1 0 2900 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_5398
timestamp 1745462530
transform 1 0 2788 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_5399
timestamp 1745462530
transform 1 0 2740 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_5400
timestamp 1745462530
transform 1 0 2988 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_5401
timestamp 1745462530
transform 1 0 2964 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_5402
timestamp 1745462530
transform 1 0 2932 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_5403
timestamp 1745462530
transform 1 0 2884 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_5404
timestamp 1745462530
transform 1 0 2436 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_5405
timestamp 1745462530
transform 1 0 2412 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_5406
timestamp 1745462530
transform 1 0 2772 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_5407
timestamp 1745462530
transform 1 0 2692 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_5408
timestamp 1745462530
transform 1 0 1796 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_5409
timestamp 1745462530
transform 1 0 1756 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_5410
timestamp 1745462530
transform 1 0 1716 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_5411
timestamp 1745462530
transform 1 0 1700 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_5412
timestamp 1745462530
transform 1 0 1692 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_5413
timestamp 1745462530
transform 1 0 1660 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_5414
timestamp 1745462530
transform 1 0 1644 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_5415
timestamp 1745462530
transform 1 0 1540 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_5416
timestamp 1745462530
transform 1 0 1508 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_5417
timestamp 1745462530
transform 1 0 1948 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_5418
timestamp 1745462530
transform 1 0 1948 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_5419
timestamp 1745462530
transform 1 0 1884 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_5420
timestamp 1745462530
transform 1 0 1884 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_5421
timestamp 1745462530
transform 1 0 2164 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_5422
timestamp 1745462530
transform 1 0 2108 0 1 1155
box -2 -2 2 2
use M2_M1  M2_M1_5423
timestamp 1745462530
transform 1 0 2068 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_5424
timestamp 1745462530
transform 1 0 2052 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_5425
timestamp 1745462530
transform 1 0 1460 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_5426
timestamp 1745462530
transform 1 0 1284 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_5427
timestamp 1745462530
transform 1 0 1252 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_5428
timestamp 1745462530
transform 1 0 2100 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_5429
timestamp 1745462530
transform 1 0 1972 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_5430
timestamp 1745462530
transform 1 0 1340 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_5431
timestamp 1745462530
transform 1 0 1220 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_5432
timestamp 1745462530
transform 1 0 1796 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_5433
timestamp 1745462530
transform 1 0 1748 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_5434
timestamp 1745462530
transform 1 0 1636 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_5435
timestamp 1745462530
transform 1 0 1636 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_5436
timestamp 1745462530
transform 1 0 1580 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_5437
timestamp 1745462530
transform 1 0 1532 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_5438
timestamp 1745462530
transform 1 0 1484 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_5439
timestamp 1745462530
transform 1 0 1972 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_5440
timestamp 1745462530
transform 1 0 1924 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_5441
timestamp 1745462530
transform 1 0 1884 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_5442
timestamp 1745462530
transform 1 0 1876 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_5443
timestamp 1745462530
transform 1 0 2236 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_5444
timestamp 1745462530
transform 1 0 2188 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_5445
timestamp 1745462530
transform 1 0 2116 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_5446
timestamp 1745462530
transform 1 0 2036 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_5447
timestamp 1745462530
transform 1 0 1396 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_5448
timestamp 1745462530
transform 1 0 1244 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_5449
timestamp 1745462530
transform 1 0 1148 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_5450
timestamp 1745462530
transform 1 0 1372 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_5451
timestamp 1745462530
transform 1 0 1324 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_5452
timestamp 1745462530
transform 1 0 1252 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_5453
timestamp 1745462530
transform 1 0 1052 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_5454
timestamp 1745462530
transform 1 0 1828 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_5455
timestamp 1745462530
transform 1 0 1764 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_5456
timestamp 1745462530
transform 1 0 1700 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_5457
timestamp 1745462530
transform 1 0 1700 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_5458
timestamp 1745462530
transform 1 0 1604 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_5459
timestamp 1745462530
transform 1 0 1556 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_5460
timestamp 1745462530
transform 1 0 1500 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_5461
timestamp 1745462530
transform 1 0 1396 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_5462
timestamp 1745462530
transform 1 0 1980 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_5463
timestamp 1745462530
transform 1 0 1924 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_5464
timestamp 1745462530
transform 1 0 1836 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_5465
timestamp 1745462530
transform 1 0 2140 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_5466
timestamp 1745462530
transform 1 0 2092 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_5467
timestamp 1745462530
transform 1 0 1980 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_5468
timestamp 1745462530
transform 1 0 1964 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_5469
timestamp 1745462530
transform 1 0 1372 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_5470
timestamp 1745462530
transform 1 0 1252 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_5471
timestamp 1745462530
transform 1 0 1124 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_5472
timestamp 1745462530
transform 1 0 1372 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_5473
timestamp 1745462530
transform 1 0 1252 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_5474
timestamp 1745462530
transform 1 0 1116 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_5475
timestamp 1745462530
transform 1 0 1796 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_5476
timestamp 1745462530
transform 1 0 1684 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_5477
timestamp 1745462530
transform 1 0 1628 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_5478
timestamp 1745462530
transform 1 0 1628 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_5479
timestamp 1745462530
transform 1 0 1652 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_5480
timestamp 1745462530
transform 1 0 1540 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_5481
timestamp 1745462530
transform 1 0 1484 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_5482
timestamp 1745462530
transform 1 0 1468 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_5483
timestamp 1745462530
transform 1 0 2060 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_5484
timestamp 1745462530
transform 1 0 1948 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_5485
timestamp 1745462530
transform 1 0 1884 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_5486
timestamp 1745462530
transform 1 0 1772 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_5487
timestamp 1745462530
transform 1 0 2068 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_5488
timestamp 1745462530
transform 1 0 2028 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_5489
timestamp 1745462530
transform 1 0 1948 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_5490
timestamp 1745462530
transform 1 0 1948 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_5491
timestamp 1745462530
transform 1 0 1356 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_5492
timestamp 1745462530
transform 1 0 1340 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_5493
timestamp 1745462530
transform 1 0 1196 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_5494
timestamp 1745462530
transform 1 0 1076 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_5495
timestamp 1745462530
transform 1 0 1260 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_5496
timestamp 1745462530
transform 1 0 1196 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_5497
timestamp 1745462530
transform 1 0 1044 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_5498
timestamp 1745462530
transform 1 0 1756 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_5499
timestamp 1745462530
transform 1 0 1732 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_5500
timestamp 1745462530
transform 1 0 1676 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_5501
timestamp 1745462530
transform 1 0 1468 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_5502
timestamp 1745462530
transform 1 0 1436 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_5503
timestamp 1745462530
transform 1 0 1404 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_5504
timestamp 1745462530
transform 1 0 1900 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_5505
timestamp 1745462530
transform 1 0 1884 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_5506
timestamp 1745462530
transform 1 0 1788 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_5507
timestamp 1745462530
transform 1 0 2124 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_5508
timestamp 1745462530
transform 1 0 2060 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_5509
timestamp 1745462530
transform 1 0 1940 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_5510
timestamp 1745462530
transform 1 0 1292 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_5511
timestamp 1745462530
transform 1 0 1268 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_5512
timestamp 1745462530
transform 1 0 1220 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_5513
timestamp 1745462530
transform 1 0 1204 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_5514
timestamp 1745462530
transform 1 0 1172 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_5515
timestamp 1745462530
transform 1 0 1460 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_5516
timestamp 1745462530
transform 1 0 1412 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_5517
timestamp 1745462530
transform 1 0 1868 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_5518
timestamp 1745462530
transform 1 0 1844 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_5519
timestamp 1745462530
transform 1 0 2060 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_5520
timestamp 1745462530
transform 1 0 1948 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_5521
timestamp 1745462530
transform 1 0 1276 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_5522
timestamp 1745462530
transform 1 0 1212 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_5523
timestamp 1745462530
transform 1 0 1332 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_5524
timestamp 1745462530
transform 1 0 1220 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_5525
timestamp 1745462530
transform 1 0 1828 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_5526
timestamp 1745462530
transform 1 0 1724 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_5527
timestamp 1745462530
transform 1 0 1692 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_5528
timestamp 1745462530
transform 1 0 1580 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_5529
timestamp 1745462530
transform 1 0 1524 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_5530
timestamp 1745462530
transform 1 0 1468 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_5531
timestamp 1745462530
transform 1 0 1876 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_5532
timestamp 1745462530
transform 1 0 1868 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_5533
timestamp 1745462530
transform 1 0 1820 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_5534
timestamp 1745462530
transform 1 0 2124 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_5535
timestamp 1745462530
transform 1 0 2068 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_5536
timestamp 1745462530
transform 1 0 2052 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_5537
timestamp 1745462530
transform 1 0 1092 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_5538
timestamp 1745462530
transform 1 0 1076 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_5539
timestamp 1745462530
transform 1 0 1044 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_5540
timestamp 1745462530
transform 1 0 996 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_5541
timestamp 1745462530
transform 1 0 980 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_5542
timestamp 1745462530
transform 1 0 1476 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_5543
timestamp 1745462530
transform 1 0 1460 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_5544
timestamp 1745462530
transform 1 0 1756 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_5545
timestamp 1745462530
transform 1 0 1748 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_5546
timestamp 1745462530
transform 1 0 1652 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_5547
timestamp 1745462530
transform 1 0 1572 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_5548
timestamp 1745462530
transform 1 0 924 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_5549
timestamp 1745462530
transform 1 0 772 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_5550
timestamp 1745462530
transform 1 0 668 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_5551
timestamp 1745462530
transform 1 0 644 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_5552
timestamp 1745462530
transform 1 0 996 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_5553
timestamp 1745462530
transform 1 0 724 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_5554
timestamp 1745462530
transform 1 0 660 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_5555
timestamp 1745462530
transform 1 0 932 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_5556
timestamp 1745462530
transform 1 0 780 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_5557
timestamp 1745462530
transform 1 0 764 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_5558
timestamp 1745462530
transform 1 0 1020 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_5559
timestamp 1745462530
transform 1 0 900 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_5560
timestamp 1745462530
transform 1 0 900 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_5561
timestamp 1745462530
transform 1 0 852 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_5562
timestamp 1745462530
transform 1 0 1148 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_5563
timestamp 1745462530
transform 1 0 1100 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_5564
timestamp 1745462530
transform 1 0 1012 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_5565
timestamp 1745462530
transform 1 0 988 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_5566
timestamp 1745462530
transform 1 0 1084 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_5567
timestamp 1745462530
transform 1 0 900 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_5568
timestamp 1745462530
transform 1 0 836 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_5569
timestamp 1745462530
transform 1 0 836 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_5570
timestamp 1745462530
transform 1 0 628 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_5571
timestamp 1745462530
transform 1 0 620 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_5572
timestamp 1745462530
transform 1 0 540 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_5573
timestamp 1745462530
transform 1 0 516 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_5574
timestamp 1745462530
transform 1 0 668 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_5575
timestamp 1745462530
transform 1 0 612 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_5576
timestamp 1745462530
transform 1 0 540 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_5577
timestamp 1745462530
transform 1 0 412 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_5578
timestamp 1745462530
transform 1 0 708 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_5579
timestamp 1745462530
transform 1 0 596 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_5580
timestamp 1745462530
transform 1 0 364 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_5581
timestamp 1745462530
transform 1 0 364 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_5582
timestamp 1745462530
transform 1 0 788 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_5583
timestamp 1745462530
transform 1 0 748 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_5584
timestamp 1745462530
transform 1 0 196 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_5585
timestamp 1745462530
transform 1 0 148 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_5586
timestamp 1745462530
transform 1 0 956 0 1 1195
box -2 -2 2 2
use M2_M1  M2_M1_5587
timestamp 1745462530
transform 1 0 908 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_5588
timestamp 1745462530
transform 1 0 180 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_5589
timestamp 1745462530
transform 1 0 908 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_5590
timestamp 1745462530
transform 1 0 780 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_5591
timestamp 1745462530
transform 1 0 460 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_5592
timestamp 1745462530
transform 1 0 460 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_5593
timestamp 1745462530
transform 1 0 876 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_5594
timestamp 1745462530
transform 1 0 844 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_5595
timestamp 1745462530
transform 1 0 828 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_5596
timestamp 1745462530
transform 1 0 724 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_5597
timestamp 1745462530
transform 1 0 1020 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_5598
timestamp 1745462530
transform 1 0 1004 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_5599
timestamp 1745462530
transform 1 0 932 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_5600
timestamp 1745462530
transform 1 0 716 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_5601
timestamp 1745462530
transform 1 0 964 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_5602
timestamp 1745462530
transform 1 0 892 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_5603
timestamp 1745462530
transform 1 0 868 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_5604
timestamp 1745462530
transform 1 0 804 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_5605
timestamp 1745462530
transform 1 0 980 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_5606
timestamp 1745462530
transform 1 0 972 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_5607
timestamp 1745462530
transform 1 0 956 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_5608
timestamp 1745462530
transform 1 0 940 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_5609
timestamp 1745462530
transform 1 0 964 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_5610
timestamp 1745462530
transform 1 0 948 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_5611
timestamp 1745462530
transform 1 0 916 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_5612
timestamp 1745462530
transform 1 0 1004 0 1 905
box -2 -2 2 2
use M2_M1  M2_M1_5613
timestamp 1745462530
transform 1 0 820 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_5614
timestamp 1745462530
transform 1 0 804 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_5615
timestamp 1745462530
transform 1 0 772 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_5616
timestamp 1745462530
transform 1 0 652 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_5617
timestamp 1745462530
transform 1 0 652 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_5618
timestamp 1745462530
transform 1 0 628 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_5619
timestamp 1745462530
transform 1 0 772 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_5620
timestamp 1745462530
transform 1 0 676 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_5621
timestamp 1745462530
transform 1 0 644 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_5622
timestamp 1745462530
transform 1 0 620 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_5623
timestamp 1745462530
transform 1 0 612 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_5624
timestamp 1745462530
transform 1 0 716 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_5625
timestamp 1745462530
transform 1 0 572 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_5626
timestamp 1745462530
transform 1 0 572 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_5627
timestamp 1745462530
transform 1 0 532 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_5628
timestamp 1745462530
transform 1 0 916 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_5629
timestamp 1745462530
transform 1 0 876 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_5630
timestamp 1745462530
transform 1 0 852 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_5631
timestamp 1745462530
transform 1 0 804 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_5632
timestamp 1745462530
transform 1 0 756 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_5633
timestamp 1745462530
transform 1 0 868 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_5634
timestamp 1745462530
transform 1 0 836 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_5635
timestamp 1745462530
transform 1 0 740 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_5636
timestamp 1745462530
transform 1 0 788 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_5637
timestamp 1745462530
transform 1 0 788 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_5638
timestamp 1745462530
transform 1 0 676 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_5639
timestamp 1745462530
transform 1 0 668 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_5640
timestamp 1745462530
transform 1 0 900 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_5641
timestamp 1745462530
transform 1 0 652 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_5642
timestamp 1745462530
transform 1 0 612 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_5643
timestamp 1745462530
transform 1 0 1076 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_5644
timestamp 1745462530
transform 1 0 468 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_5645
timestamp 1745462530
transform 1 0 444 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_5646
timestamp 1745462530
transform 1 0 1012 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_5647
timestamp 1745462530
transform 1 0 364 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_5648
timestamp 1745462530
transform 1 0 356 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_5649
timestamp 1745462530
transform 1 0 1036 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_5650
timestamp 1745462530
transform 1 0 276 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_5651
timestamp 1745462530
transform 1 0 180 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_5652
timestamp 1745462530
transform 1 0 980 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_5653
timestamp 1745462530
transform 1 0 300 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_5654
timestamp 1745462530
transform 1 0 180 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_5655
timestamp 1745462530
transform 1 0 1044 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_5656
timestamp 1745462530
transform 1 0 588 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_5657
timestamp 1745462530
transform 1 0 532 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_5658
timestamp 1745462530
transform 1 0 388 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_5659
timestamp 1745462530
transform 1 0 356 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_5660
timestamp 1745462530
transform 1 0 180 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_5661
timestamp 1745462530
transform 1 0 156 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_5662
timestamp 1745462530
transform 1 0 500 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_5663
timestamp 1745462530
transform 1 0 292 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_5664
timestamp 1745462530
transform 1 0 180 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_5665
timestamp 1745462530
transform 1 0 548 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_5666
timestamp 1745462530
transform 1 0 428 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_5667
timestamp 1745462530
transform 1 0 564 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_5668
timestamp 1745462530
transform 1 0 420 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_5669
timestamp 1745462530
transform 1 0 356 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_5670
timestamp 1745462530
transform 1 0 708 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_5671
timestamp 1745462530
transform 1 0 236 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_5672
timestamp 1745462530
transform 1 0 188 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_5673
timestamp 1745462530
transform 1 0 844 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_5674
timestamp 1745462530
transform 1 0 236 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_5675
timestamp 1745462530
transform 1 0 180 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_5676
timestamp 1745462530
transform 1 0 844 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_5677
timestamp 1745462530
transform 1 0 412 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_5678
timestamp 1745462530
transform 1 0 348 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_5679
timestamp 1745462530
transform 1 0 940 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5680
timestamp 1745462530
transform 1 0 756 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5681
timestamp 1745462530
transform 1 0 668 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_5682
timestamp 1745462530
transform 1 0 620 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5683
timestamp 1745462530
transform 1 0 988 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_5684
timestamp 1745462530
transform 1 0 916 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_5685
timestamp 1745462530
transform 1 0 812 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5686
timestamp 1745462530
transform 1 0 772 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_5687
timestamp 1745462530
transform 1 0 900 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_5688
timestamp 1745462530
transform 1 0 676 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5689
timestamp 1745462530
transform 1 0 628 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_5690
timestamp 1745462530
transform 1 0 628 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_5691
timestamp 1745462530
transform 1 0 900 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5692
timestamp 1745462530
transform 1 0 900 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_5693
timestamp 1745462530
transform 1 0 844 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_5694
timestamp 1745462530
transform 1 0 724 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_5695
timestamp 1745462530
transform 1 0 980 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_5696
timestamp 1745462530
transform 1 0 964 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5697
timestamp 1745462530
transform 1 0 876 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_5698
timestamp 1745462530
transform 1 0 748 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_5699
timestamp 1745462530
transform 1 0 852 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_5700
timestamp 1745462530
transform 1 0 828 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5701
timestamp 1745462530
transform 1 0 580 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_5702
timestamp 1745462530
transform 1 0 580 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_5703
timestamp 1745462530
transform 1 0 692 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5704
timestamp 1745462530
transform 1 0 540 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_5705
timestamp 1745462530
transform 1 0 316 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5706
timestamp 1745462530
transform 1 0 300 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5707
timestamp 1745462530
transform 1 0 764 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5708
timestamp 1745462530
transform 1 0 668 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_5709
timestamp 1745462530
transform 1 0 452 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5710
timestamp 1745462530
transform 1 0 644 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5711
timestamp 1745462530
transform 1 0 628 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5712
timestamp 1745462530
transform 1 0 628 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5713
timestamp 1745462530
transform 1 0 524 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_5714
timestamp 1745462530
transform 1 0 460 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_5715
timestamp 1745462530
transform 1 0 836 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5716
timestamp 1745462530
transform 1 0 748 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_5717
timestamp 1745462530
transform 1 0 388 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_5718
timestamp 1745462530
transform 1 0 380 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_5719
timestamp 1745462530
transform 1 0 908 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5720
timestamp 1745462530
transform 1 0 884 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5721
timestamp 1745462530
transform 1 0 268 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_5722
timestamp 1745462530
transform 1 0 204 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_5723
timestamp 1745462530
transform 1 0 780 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_5724
timestamp 1745462530
transform 1 0 772 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5725
timestamp 1745462530
transform 1 0 180 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5726
timestamp 1745462530
transform 1 0 900 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_5727
timestamp 1745462530
transform 1 0 652 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5728
timestamp 1745462530
transform 1 0 316 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5729
timestamp 1745462530
transform 1 0 308 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5730
timestamp 1745462530
transform 1 0 1036 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5731
timestamp 1745462530
transform 1 0 668 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_5732
timestamp 1745462530
transform 1 0 556 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5733
timestamp 1745462530
transform 1 0 452 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5734
timestamp 1745462530
transform 1 0 868 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5735
timestamp 1745462530
transform 1 0 628 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5736
timestamp 1745462530
transform 1 0 500 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_5737
timestamp 1745462530
transform 1 0 500 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5738
timestamp 1745462530
transform 1 0 932 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5739
timestamp 1745462530
transform 1 0 828 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_5740
timestamp 1745462530
transform 1 0 388 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5741
timestamp 1745462530
transform 1 0 348 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5742
timestamp 1745462530
transform 1 0 1020 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_5743
timestamp 1745462530
transform 1 0 844 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_5744
timestamp 1745462530
transform 1 0 172 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_5745
timestamp 1745462530
transform 1 0 972 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5746
timestamp 1745462530
transform 1 0 740 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5747
timestamp 1745462530
transform 1 0 180 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5748
timestamp 1745462530
transform 1 0 604 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5749
timestamp 1745462530
transform 1 0 540 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_5750
timestamp 1745462530
transform 1 0 516 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_5751
timestamp 1745462530
transform 1 0 364 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_5752
timestamp 1745462530
transform 1 0 308 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_5753
timestamp 1745462530
transform 1 0 620 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_5754
timestamp 1745462530
transform 1 0 612 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_5755
timestamp 1745462530
transform 1 0 500 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_5756
timestamp 1745462530
transform 1 0 436 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_5757
timestamp 1745462530
transform 1 0 580 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_5758
timestamp 1745462530
transform 1 0 580 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_5759
timestamp 1745462530
transform 1 0 508 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_5760
timestamp 1745462530
transform 1 0 388 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_5761
timestamp 1745462530
transform 1 0 772 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5762
timestamp 1745462530
transform 1 0 756 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_5763
timestamp 1745462530
transform 1 0 436 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_5764
timestamp 1745462530
transform 1 0 364 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_5765
timestamp 1745462530
transform 1 0 852 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_5766
timestamp 1745462530
transform 1 0 804 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5767
timestamp 1745462530
transform 1 0 180 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_5768
timestamp 1745462530
transform 1 0 180 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5769
timestamp 1745462530
transform 1 0 764 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_5770
timestamp 1745462530
transform 1 0 692 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5771
timestamp 1745462530
transform 1 0 252 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_5772
timestamp 1745462530
transform 1 0 172 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_5773
timestamp 1745462530
transform 1 0 988 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_5774
timestamp 1745462530
transform 1 0 940 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_5775
timestamp 1745462530
transform 1 0 900 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_5776
timestamp 1745462530
transform 1 0 1204 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_5777
timestamp 1745462530
transform 1 0 1076 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5778
timestamp 1745462530
transform 1 0 1004 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_5779
timestamp 1745462530
transform 1 0 1092 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_5780
timestamp 1745462530
transform 1 0 916 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_5781
timestamp 1745462530
transform 1 0 916 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5782
timestamp 1745462530
transform 1 0 1092 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_5783
timestamp 1745462530
transform 1 0 964 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5784
timestamp 1745462530
transform 1 0 908 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_5785
timestamp 1745462530
transform 1 0 1076 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_5786
timestamp 1745462530
transform 1 0 1060 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_5787
timestamp 1745462530
transform 1 0 1020 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_5788
timestamp 1745462530
transform 1 0 1060 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_5789
timestamp 1745462530
transform 1 0 1036 0 1 2045
box -2 -2 2 2
use M2_M1  M2_M1_5790
timestamp 1745462530
transform 1 0 972 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_5791
timestamp 1745462530
transform 1 0 972 0 1 2195
box -2 -2 2 2
use M2_M1  M2_M1_5792
timestamp 1745462530
transform 1 0 956 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_5793
timestamp 1745462530
transform 1 0 524 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_5794
timestamp 1745462530
transform 1 0 476 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_5795
timestamp 1745462530
transform 1 0 172 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_5796
timestamp 1745462530
transform 1 0 172 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_5797
timestamp 1745462530
transform 1 0 596 0 1 2395
box -2 -2 2 2
use M2_M1  M2_M1_5798
timestamp 1745462530
transform 1 0 548 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_5799
timestamp 1745462530
transform 1 0 508 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_5800
timestamp 1745462530
transform 1 0 644 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_5801
timestamp 1745462530
transform 1 0 628 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_5802
timestamp 1745462530
transform 1 0 620 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_5803
timestamp 1745462530
transform 1 0 612 0 1 2555
box -2 -2 2 2
use M2_M1  M2_M1_5804
timestamp 1745462530
transform 1 0 612 0 1 2495
box -2 -2 2 2
use M2_M1  M2_M1_5805
timestamp 1745462530
transform 1 0 564 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5806
timestamp 1745462530
transform 1 0 548 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_5807
timestamp 1745462530
transform 1 0 484 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_5808
timestamp 1745462530
transform 1 0 732 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_5809
timestamp 1745462530
transform 1 0 716 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_5810
timestamp 1745462530
transform 1 0 716 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_5811
timestamp 1745462530
transform 1 0 892 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_5812
timestamp 1745462530
transform 1 0 852 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5813
timestamp 1745462530
transform 1 0 812 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_5814
timestamp 1745462530
transform 1 0 732 0 1 2395
box -2 -2 2 2
use M2_M1  M2_M1_5815
timestamp 1745462530
transform 1 0 612 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_5816
timestamp 1745462530
transform 1 0 572 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_5817
timestamp 1745462530
transform 1 0 572 0 1 2645
box -2 -2 2 2
use M2_M1  M2_M1_5818
timestamp 1745462530
transform 1 0 572 0 1 2625
box -2 -2 2 2
use M2_M1  M2_M1_5819
timestamp 1745462530
transform 1 0 412 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_5820
timestamp 1745462530
transform 1 0 364 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_5821
timestamp 1745462530
transform 1 0 836 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_5822
timestamp 1745462530
transform 1 0 796 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_5823
timestamp 1745462530
transform 1 0 948 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_5824
timestamp 1745462530
transform 1 0 868 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_5825
timestamp 1745462530
transform 1 0 196 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_5826
timestamp 1745462530
transform 1 0 180 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_5827
timestamp 1745462530
transform 1 0 2004 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_5828
timestamp 1745462530
transform 1 0 1844 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_5829
timestamp 1745462530
transform 1 0 1316 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_5830
timestamp 1745462530
transform 1 0 1220 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_5831
timestamp 1745462530
transform 1 0 1204 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_5832
timestamp 1745462530
transform 1 0 1196 0 1 1785
box -2 -2 2 2
use M2_M1  M2_M1_5833
timestamp 1745462530
transform 1 0 1636 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_5834
timestamp 1745462530
transform 1 0 1516 0 1 1795
box -2 -2 2 2
use M2_M1  M2_M1_5835
timestamp 1745462530
transform 1 0 1516 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_5836
timestamp 1745462530
transform 1 0 1972 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5837
timestamp 1745462530
transform 1 0 1908 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_5838
timestamp 1745462530
transform 1 0 1852 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5839
timestamp 1745462530
transform 1 0 1204 0 1 1985
box -2 -2 2 2
use M2_M1  M2_M1_5840
timestamp 1745462530
transform 1 0 1148 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_5841
timestamp 1745462530
transform 1 0 1124 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5842
timestamp 1745462530
transform 1 0 1420 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_5843
timestamp 1745462530
transform 1 0 1412 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_5844
timestamp 1745462530
transform 1 0 1340 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_5845
timestamp 1745462530
transform 1 0 2060 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_5846
timestamp 1745462530
transform 1 0 1820 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_5847
timestamp 1745462530
transform 1 0 1372 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_5848
timestamp 1745462530
transform 1 0 1292 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_5849
timestamp 1745462530
transform 1 0 1276 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_5850
timestamp 1745462530
transform 1 0 1684 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_5851
timestamp 1745462530
transform 1 0 1660 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_5852
timestamp 1745462530
transform 1 0 1572 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_5853
timestamp 1745462530
transform 1 0 1996 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_5854
timestamp 1745462530
transform 1 0 1820 0 1 2545
box -2 -2 2 2
use M2_M1  M2_M1_5855
timestamp 1745462530
transform 1 0 1812 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_5856
timestamp 1745462530
transform 1 0 1180 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_5857
timestamp 1745462530
transform 1 0 1156 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_5858
timestamp 1745462530
transform 1 0 1500 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_5859
timestamp 1745462530
transform 1 0 1468 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_5860
timestamp 1745462530
transform 1 0 1396 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_5861
timestamp 1745462530
transform 1 0 2172 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5862
timestamp 1745462530
transform 1 0 2036 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5863
timestamp 1745462530
transform 1 0 2004 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5864
timestamp 1745462530
transform 1 0 1388 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5865
timestamp 1745462530
transform 1 0 1308 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5866
timestamp 1745462530
transform 1 0 1276 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5867
timestamp 1745462530
transform 1 0 1276 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5868
timestamp 1745462530
transform 1 0 1764 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5869
timestamp 1745462530
transform 1 0 1636 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5870
timestamp 1745462530
transform 1 0 1636 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5871
timestamp 1745462530
transform 1 0 2060 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5872
timestamp 1745462530
transform 1 0 1900 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5873
timestamp 1745462530
transform 1 0 1884 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5874
timestamp 1745462530
transform 1 0 1132 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5875
timestamp 1745462530
transform 1 0 1084 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5876
timestamp 1745462530
transform 1 0 1460 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5877
timestamp 1745462530
transform 1 0 1460 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5878
timestamp 1745462530
transform 1 0 1452 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_5879
timestamp 1745462530
transform 1 0 2092 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_5880
timestamp 1745462530
transform 1 0 2020 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_5881
timestamp 1745462530
transform 1 0 2004 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_5882
timestamp 1745462530
transform 1 0 1324 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_5883
timestamp 1745462530
transform 1 0 1316 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_5884
timestamp 1745462530
transform 1 0 1308 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_5885
timestamp 1745462530
transform 1 0 1812 0 1 2705
box -2 -2 2 2
use M2_M1  M2_M1_5886
timestamp 1745462530
transform 1 0 1652 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_5887
timestamp 1745462530
transform 1 0 1620 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_5888
timestamp 1745462530
transform 1 0 1956 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_5889
timestamp 1745462530
transform 1 0 1868 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_5890
timestamp 1745462530
transform 1 0 1860 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_5891
timestamp 1745462530
transform 1 0 1204 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_5892
timestamp 1745462530
transform 1 0 1164 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_5893
timestamp 1745462530
transform 1 0 1604 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_5894
timestamp 1745462530
transform 1 0 1516 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_5895
timestamp 1745462530
transform 1 0 1468 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_5896
timestamp 1745462530
transform 1 0 2132 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5897
timestamp 1745462530
transform 1 0 2068 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5898
timestamp 1745462530
transform 1 0 2028 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_5899
timestamp 1745462530
transform 1 0 2020 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_5900
timestamp 1745462530
transform 1 0 1396 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_5901
timestamp 1745462530
transform 1 0 1364 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_5902
timestamp 1745462530
transform 1 0 1356 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5903
timestamp 1745462530
transform 1 0 1340 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_5904
timestamp 1745462530
transform 1 0 1748 0 1 2185
box -2 -2 2 2
use M2_M1  M2_M1_5905
timestamp 1745462530
transform 1 0 1732 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5906
timestamp 1745462530
transform 1 0 1732 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_5907
timestamp 1745462530
transform 1 0 1708 0 1 1955
box -2 -2 2 2
use M2_M1  M2_M1_5908
timestamp 1745462530
transform 1 0 1692 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_5909
timestamp 1745462530
transform 1 0 1660 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_5910
timestamp 1745462530
transform 1 0 1996 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_5911
timestamp 1745462530
transform 1 0 1964 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_5912
timestamp 1745462530
transform 1 0 1948 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5913
timestamp 1745462530
transform 1 0 1932 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_5914
timestamp 1745462530
transform 1 0 1236 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_5915
timestamp 1745462530
transform 1 0 1188 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_5916
timestamp 1745462530
transform 1 0 1124 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_5917
timestamp 1745462530
transform 1 0 1116 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5918
timestamp 1745462530
transform 1 0 1628 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_5919
timestamp 1745462530
transform 1 0 1564 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_5920
timestamp 1745462530
transform 1 0 1524 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_5921
timestamp 1745462530
transform 1 0 1516 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_5922
timestamp 1745462530
transform 1 0 2020 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_5923
timestamp 1745462530
transform 1 0 1964 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_5924
timestamp 1745462530
transform 1 0 1964 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_5925
timestamp 1745462530
transform 1 0 1420 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_5926
timestamp 1745462530
transform 1 0 1380 0 1 2625
box -2 -2 2 2
use M2_M1  M2_M1_5927
timestamp 1745462530
transform 1 0 1380 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_5928
timestamp 1745462530
transform 1 0 1372 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_5929
timestamp 1745462530
transform 1 0 1340 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_5930
timestamp 1745462530
transform 1 0 1788 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_5931
timestamp 1745462530
transform 1 0 1716 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_5932
timestamp 1745462530
transform 1 0 1652 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_5933
timestamp 1745462530
transform 1 0 1900 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_5934
timestamp 1745462530
transform 1 0 1900 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_5935
timestamp 1745462530
transform 1 0 1844 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_5936
timestamp 1745462530
transform 1 0 1180 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_5937
timestamp 1745462530
transform 1 0 1148 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_5938
timestamp 1745462530
transform 1 0 1636 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_5939
timestamp 1745462530
transform 1 0 1564 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_5940
timestamp 1745462530
transform 1 0 1532 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_5941
timestamp 1745462530
transform 1 0 2852 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_5942
timestamp 1745462530
transform 1 0 2748 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_5943
timestamp 1745462530
transform 1 0 2020 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_5944
timestamp 1745462530
transform 1 0 2012 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_5945
timestamp 1745462530
transform 1 0 2764 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_5946
timestamp 1745462530
transform 1 0 1452 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_5947
timestamp 1745462530
transform 1 0 1340 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_5948
timestamp 1745462530
transform 1 0 2588 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_5949
timestamp 1745462530
transform 1 0 2572 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_5950
timestamp 1745462530
transform 1 0 1684 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_5951
timestamp 1745462530
transform 1 0 1628 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_5952
timestamp 1745462530
transform 1 0 2476 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_5953
timestamp 1745462530
transform 1 0 2468 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_5954
timestamp 1745462530
transform 1 0 1964 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_5955
timestamp 1745462530
transform 1 0 1948 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_5956
timestamp 1745462530
transform 1 0 2740 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_5957
timestamp 1745462530
transform 1 0 2660 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_5958
timestamp 1745462530
transform 1 0 1468 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_5959
timestamp 1745462530
transform 1 0 1148 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_5960
timestamp 1745462530
transform 1 0 2604 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_5961
timestamp 1745462530
transform 1 0 2556 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_5962
timestamp 1745462530
transform 1 0 1524 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_5963
timestamp 1745462530
transform 1 0 1444 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_5964
timestamp 1745462530
transform 1 0 3196 0 1 2145
box -2 -2 2 2
use M2_M1  M2_M1_5965
timestamp 1745462530
transform 1 0 3092 0 1 2745
box -2 -2 2 2
use M2_M1  M2_M1_5966
timestamp 1745462530
transform 1 0 3028 0 1 2595
box -2 -2 2 2
use M2_M1  M2_M1_5967
timestamp 1745462530
transform 1 0 2996 0 1 2795
box -2 -2 2 2
use M2_M1  M2_M1_5968
timestamp 1745462530
transform 1 0 2956 0 1 2145
box -2 -2 2 2
use M2_M1  M2_M1_5969
timestamp 1745462530
transform 1 0 2436 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5970
timestamp 1745462530
transform 1 0 1540 0 1 2345
box -2 -2 2 2
use M2_M1  M2_M1_5971
timestamp 1745462530
transform 1 0 1508 0 1 2545
box -2 -2 2 2
use M2_M1  M2_M1_5972
timestamp 1745462530
transform 1 0 1492 0 1 2795
box -2 -2 2 2
use M2_M1  M2_M1_5973
timestamp 1745462530
transform 1 0 1492 0 1 2545
box -2 -2 2 2
use M2_M1  M2_M1_5974
timestamp 1745462530
transform 1 0 1404 0 1 3145
box -2 -2 2 2
use M2_M1  M2_M1_5975
timestamp 1745462530
transform 1 0 1340 0 1 3195
box -2 -2 2 2
use M2_M1  M2_M1_5976
timestamp 1745462530
transform 1 0 1316 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_5977
timestamp 1745462530
transform 1 0 1292 0 1 3345
box -2 -2 2 2
use M2_M1  M2_M1_5978
timestamp 1745462530
transform 1 0 956 0 1 3545
box -2 -2 2 2
use M2_M1  M2_M1_5979
timestamp 1745462530
transform 1 0 956 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_5980
timestamp 1745462530
transform 1 0 948 0 1 3395
box -2 -2 2 2
use M2_M1  M2_M1_5981
timestamp 1745462530
transform 1 0 924 0 1 3545
box -2 -2 2 2
use M2_M1  M2_M1_5982
timestamp 1745462530
transform 1 0 908 0 1 3395
box -2 -2 2 2
use M2_M1  M2_M1_5983
timestamp 1745462530
transform 1 0 748 0 1 1945
box -2 -2 2 2
use M2_M1  M2_M1_5984
timestamp 1745462530
transform 1 0 660 0 1 1995
box -2 -2 2 2
use M2_M1  M2_M1_5985
timestamp 1745462530
transform 1 0 644 0 1 3235
box -2 -2 2 2
use M2_M1  M2_M1_5986
timestamp 1745462530
transform 1 0 620 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_5987
timestamp 1745462530
transform 1 0 572 0 1 2105
box -2 -2 2 2
use M2_M1  M2_M1_5988
timestamp 1745462530
transform 1 0 556 0 1 2145
box -2 -2 2 2
use M2_M1  M2_M1_5989
timestamp 1745462530
transform 1 0 540 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_5990
timestamp 1745462530
transform 1 0 500 0 1 1945
box -2 -2 2 2
use M2_M1  M2_M1_5991
timestamp 1745462530
transform 1 0 1332 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_5992
timestamp 1745462530
transform 1 0 1220 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_5993
timestamp 1745462530
transform 1 0 1412 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_5994
timestamp 1745462530
transform 1 0 1340 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_5995
timestamp 1745462530
transform 1 0 1468 0 1 3425
box -2 -2 2 2
use M2_M1  M2_M1_5996
timestamp 1745462530
transform 1 0 1228 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_5997
timestamp 1745462530
transform 1 0 1428 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_5998
timestamp 1745462530
transform 1 0 1324 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_5999
timestamp 1745462530
transform 1 0 1284 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_6000
timestamp 1745462530
transform 1 0 1212 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_6001
timestamp 1745462530
transform 1 0 1420 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_6002
timestamp 1745462530
transform 1 0 1220 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_6003
timestamp 1745462530
transform 1 0 2284 0 1 2715
box -2 -2 2 2
use M2_M1  M2_M1_6004
timestamp 1745462530
transform 1 0 1604 0 1 3035
box -2 -2 2 2
use M2_M1  M2_M1_6005
timestamp 1745462530
transform 1 0 1524 0 1 2995
box -2 -2 2 2
use M2_M1  M2_M1_6006
timestamp 1745462530
transform 1 0 1124 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_6007
timestamp 1745462530
transform 1 0 1068 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_6008
timestamp 1745462530
transform 1 0 980 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_6009
timestamp 1745462530
transform 1 0 892 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_6010
timestamp 1745462530
transform 1 0 860 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_6011
timestamp 1745462530
transform 1 0 548 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_6012
timestamp 1745462530
transform 1 0 548 0 1 3115
box -2 -2 2 2
use M2_M1  M2_M1_6013
timestamp 1745462530
transform 1 0 460 0 1 3115
box -2 -2 2 2
use M2_M1  M2_M1_6014
timestamp 1745462530
transform 1 0 436 0 1 3185
box -2 -2 2 2
use M2_M1  M2_M1_6015
timestamp 1745462530
transform 1 0 356 0 1 3115
box -2 -2 2 2
use M2_M1  M2_M1_6016
timestamp 1745462530
transform 1 0 340 0 1 3185
box -2 -2 2 2
use M2_M1  M2_M1_6017
timestamp 1745462530
transform 1 0 236 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_6018
timestamp 1745462530
transform 1 0 236 0 1 3025
box -2 -2 2 2
use M2_M1  M2_M1_6019
timestamp 1745462530
transform 1 0 228 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_6020
timestamp 1745462530
transform 1 0 140 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_6021
timestamp 1745462530
transform 1 0 2092 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_6022
timestamp 1745462530
transform 1 0 860 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_6023
timestamp 1745462530
transform 1 0 2196 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_6024
timestamp 1745462530
transform 1 0 676 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_6025
timestamp 1745462530
transform 1 0 2196 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_6026
timestamp 1745462530
transform 1 0 636 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_6027
timestamp 1745462530
transform 1 0 2156 0 1 3035
box -2 -2 2 2
use M2_M1  M2_M1_6028
timestamp 1745462530
transform 1 0 532 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_6029
timestamp 1745462530
transform 1 0 2068 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_6030
timestamp 1745462530
transform 1 0 412 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_6031
timestamp 1745462530
transform 1 0 2140 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_6032
timestamp 1745462530
transform 1 0 292 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_6033
timestamp 1745462530
transform 1 0 2404 0 1 2595
box -2 -2 2 2
use M2_M1  M2_M1_6034
timestamp 1745462530
transform 1 0 2388 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_6035
timestamp 1745462530
transform 1 0 2268 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_6036
timestamp 1745462530
transform 1 0 2132 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_6037
timestamp 1745462530
transform 1 0 2532 0 1 1595
box -2 -2 2 2
use M2_M1  M2_M1_6038
timestamp 1745462530
transform 1 0 2460 0 1 1595
box -2 -2 2 2
use M2_M1  M2_M1_6039
timestamp 1745462530
transform 1 0 2420 0 1 1945
box -2 -2 2 2
use M2_M1  M2_M1_6040
timestamp 1745462530
transform 1 0 2388 0 1 1595
box -2 -2 2 2
use M2_M1  M2_M1_6041
timestamp 1745462530
transform 1 0 2324 0 1 1945
box -2 -2 2 2
use M2_M1  M2_M1_6042
timestamp 1745462530
transform 1 0 2316 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_6043
timestamp 1745462530
transform 1 0 2308 0 1 1595
box -2 -2 2 2
use M2_M1  M2_M1_6044
timestamp 1745462530
transform 1 0 2236 0 1 2635
box -2 -2 2 2
use M2_M1  M2_M1_6045
timestamp 1745462530
transform 1 0 2092 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_6046
timestamp 1745462530
transform 1 0 2212 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_6047
timestamp 1745462530
transform 1 0 2148 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_6048
timestamp 1745462530
transform 1 0 2132 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_6049
timestamp 1745462530
transform 1 0 2132 0 1 1795
box -2 -2 2 2
use M2_M1  M2_M1_6050
timestamp 1745462530
transform 1 0 2116 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_6051
timestamp 1745462530
transform 1 0 2044 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_6052
timestamp 1745462530
transform 1 0 2180 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_6053
timestamp 1745462530
transform 1 0 2172 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_6054
timestamp 1745462530
transform 1 0 2156 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_6055
timestamp 1745462530
transform 1 0 2148 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_6056
timestamp 1745462530
transform 1 0 2148 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_6057
timestamp 1745462530
transform 1 0 2108 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_6058
timestamp 1745462530
transform 1 0 3556 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_6059
timestamp 1745462530
transform 1 0 3548 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_6060
timestamp 1745462530
transform 1 0 3516 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_6061
timestamp 1745462530
transform 1 0 2788 0 1 2995
box -2 -2 2 2
use M2_M1  M2_M1_6062
timestamp 1745462530
transform 1 0 2660 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_6063
timestamp 1745462530
transform 1 0 2620 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_6064
timestamp 1745462530
transform 1 0 2596 0 1 895
box -2 -2 2 2
use M2_M1  M2_M1_6065
timestamp 1745462530
transform 1 0 2596 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_6066
timestamp 1745462530
transform 1 0 2588 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_6067
timestamp 1745462530
transform 1 0 2580 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_6068
timestamp 1745462530
transform 1 0 2564 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_6069
timestamp 1745462530
transform 1 0 2252 0 1 3115
box -2 -2 2 2
use M2_M1  M2_M1_6070
timestamp 1745462530
transform 1 0 2252 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_6071
timestamp 1745462530
transform 1 0 2204 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_6072
timestamp 1745462530
transform 1 0 1972 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_6073
timestamp 1745462530
transform 1 0 1628 0 1 3025
box -2 -2 2 2
use M2_M1  M2_M1_6074
timestamp 1745462530
transform 1 0 1140 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_6075
timestamp 1745462530
transform 1 0 1156 0 1 3825
box -2 -2 2 2
use M2_M1  M2_M1_6076
timestamp 1745462530
transform 1 0 1132 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_6077
timestamp 1745462530
transform 1 0 1236 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_6078
timestamp 1745462530
transform 1 0 1132 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_6079
timestamp 1745462530
transform 1 0 1724 0 1 3025
box -2 -2 2 2
use M2_M1  M2_M1_6080
timestamp 1745462530
transform 1 0 1212 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_6081
timestamp 1745462530
transform 1 0 1212 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_6082
timestamp 1745462530
transform 1 0 1204 0 1 3025
box -2 -2 2 2
use M2_M1  M2_M1_6083
timestamp 1745462530
transform 1 0 1356 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_6084
timestamp 1745462530
transform 1 0 1188 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_6085
timestamp 1745462530
transform 1 0 1524 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_6086
timestamp 1745462530
transform 1 0 1452 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_6087
timestamp 1745462530
transform 1 0 1436 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_6088
timestamp 1745462530
transform 1 0 1396 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_6089
timestamp 1745462530
transform 1 0 1236 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_6090
timestamp 1745462530
transform 1 0 1188 0 1 2625
box -2 -2 2 2
use M2_M1  M2_M1_6091
timestamp 1745462530
transform 1 0 1188 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_6092
timestamp 1745462530
transform 1 0 1172 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_6093
timestamp 1745462530
transform 1 0 1156 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_6094
timestamp 1745462530
transform 1 0 1780 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_6095
timestamp 1745462530
transform 1 0 1708 0 1 3025
box -2 -2 2 2
use M2_M1  M2_M1_6096
timestamp 1745462530
transform 1 0 1820 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_6097
timestamp 1745462530
transform 1 0 1716 0 1 3035
box -2 -2 2 2
use M2_M1  M2_M1_6098
timestamp 1745462530
transform 1 0 1884 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_6099
timestamp 1745462530
transform 1 0 1796 0 1 2995
box -2 -2 2 2
use M2_M1  M2_M1_6100
timestamp 1745462530
transform 1 0 1812 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_6101
timestamp 1745462530
transform 1 0 1796 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_6102
timestamp 1745462530
transform 1 0 1756 0 1 1945
box -2 -2 2 2
use M2_M1  M2_M1_6103
timestamp 1745462530
transform 1 0 1756 0 1 1905
box -2 -2 2 2
use M2_M1  M2_M1_6104
timestamp 1745462530
transform 1 0 1756 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_6105
timestamp 1745462530
transform 1 0 1740 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_6106
timestamp 1745462530
transform 1 0 1740 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_6107
timestamp 1745462530
transform 1 0 1740 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_6108
timestamp 1745462530
transform 1 0 1828 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_6109
timestamp 1745462530
transform 1 0 1820 0 1 2235
box -2 -2 2 2
use M2_M1  M2_M1_6110
timestamp 1745462530
transform 1 0 1684 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_6111
timestamp 1745462530
transform 1 0 1660 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_6112
timestamp 1745462530
transform 1 0 1548 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_6113
timestamp 1745462530
transform 1 0 1924 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_6114
timestamp 1745462530
transform 1 0 1836 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_6115
timestamp 1745462530
transform 1 0 1804 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_6116
timestamp 1745462530
transform 1 0 876 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_6117
timestamp 1745462530
transform 1 0 796 0 1 3225
box -2 -2 2 2
use M2_M1  M2_M1_6118
timestamp 1745462530
transform 1 0 796 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_6119
timestamp 1745462530
transform 1 0 996 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_6120
timestamp 1745462530
transform 1 0 948 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_6121
timestamp 1745462530
transform 1 0 924 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_6122
timestamp 1745462530
transform 1 0 812 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_6123
timestamp 1745462530
transform 1 0 828 0 1 3225
box -2 -2 2 2
use M2_M1  M2_M1_6124
timestamp 1745462530
transform 1 0 804 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_6125
timestamp 1745462530
transform 1 0 940 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_6126
timestamp 1745462530
transform 1 0 876 0 1 3195
box -2 -2 2 2
use M2_M1  M2_M1_6127
timestamp 1745462530
transform 1 0 700 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_6128
timestamp 1745462530
transform 1 0 676 0 1 3225
box -2 -2 2 2
use M2_M1  M2_M1_6129
timestamp 1745462530
transform 1 0 620 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_6130
timestamp 1745462530
transform 1 0 3156 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_6131
timestamp 1745462530
transform 1 0 3124 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_6132
timestamp 1745462530
transform 1 0 3116 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_6133
timestamp 1745462530
transform 1 0 3100 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_6134
timestamp 1745462530
transform 1 0 3092 0 1 3485
box -2 -2 2 2
use M2_M1  M2_M1_6135
timestamp 1745462530
transform 1 0 3084 0 1 3595
box -2 -2 2 2
use M2_M1  M2_M1_6136
timestamp 1745462530
transform 1 0 3084 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_6137
timestamp 1745462530
transform 1 0 3100 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_6138
timestamp 1745462530
transform 1 0 2996 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_6139
timestamp 1745462530
transform 1 0 3412 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_6140
timestamp 1745462530
transform 1 0 3348 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_6141
timestamp 1745462530
transform 1 0 3348 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_6142
timestamp 1745462530
transform 1 0 3124 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_6143
timestamp 1745462530
transform 1 0 2972 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_6144
timestamp 1745462530
transform 1 0 2780 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_6145
timestamp 1745462530
transform 1 0 2308 0 1 3595
box -2 -2 2 2
use M2_M1  M2_M1_6146
timestamp 1745462530
transform 1 0 2140 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_6147
timestamp 1745462530
transform 1 0 1732 0 1 3515
box -2 -2 2 2
use M2_M1  M2_M1_6148
timestamp 1745462530
transform 1 0 3060 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_6149
timestamp 1745462530
transform 1 0 2988 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_6150
timestamp 1745462530
transform 1 0 2988 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_6151
timestamp 1745462530
transform 1 0 2972 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_6152
timestamp 1745462530
transform 1 0 2916 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_6153
timestamp 1745462530
transform 1 0 2900 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_6154
timestamp 1745462530
transform 1 0 1948 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_6155
timestamp 1745462530
transform 1 0 1844 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_6156
timestamp 1745462530
transform 1 0 1692 0 1 3315
box -2 -2 2 2
use M2_M1  M2_M1_6157
timestamp 1745462530
transform 1 0 2204 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_6158
timestamp 1745462530
transform 1 0 2108 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_6159
timestamp 1745462530
transform 1 0 3308 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_6160
timestamp 1745462530
transform 1 0 3260 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_6161
timestamp 1745462530
transform 1 0 3228 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_6162
timestamp 1745462530
transform 1 0 3156 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_6163
timestamp 1745462530
transform 1 0 3068 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_6164
timestamp 1745462530
transform 1 0 2836 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_6165
timestamp 1745462530
transform 1 0 2396 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_6166
timestamp 1745462530
transform 1 0 2380 0 1 3315
box -2 -2 2 2
use M2_M1  M2_M1_6167
timestamp 1745462530
transform 1 0 2356 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_6168
timestamp 1745462530
transform 1 0 3076 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_6169
timestamp 1745462530
transform 1 0 3052 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_6170
timestamp 1745462530
transform 1 0 3044 0 1 3315
box -2 -2 2 2
use M2_M1  M2_M1_6171
timestamp 1745462530
transform 1 0 3004 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_6172
timestamp 1745462530
transform 1 0 2972 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_6173
timestamp 1745462530
transform 1 0 2932 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_6174
timestamp 1745462530
transform 1 0 2932 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_6175
timestamp 1745462530
transform 1 0 2820 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_6176
timestamp 1745462530
transform 1 0 2820 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_6177
timestamp 1745462530
transform 1 0 3100 0 1 3425
box -2 -2 2 2
use M2_M1  M2_M1_6178
timestamp 1745462530
transform 1 0 3052 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_6179
timestamp 1745462530
transform 1 0 2004 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_6180
timestamp 1745462530
transform 1 0 1948 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_6181
timestamp 1745462530
transform 1 0 3244 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_6182
timestamp 1745462530
transform 1 0 3220 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_6183
timestamp 1745462530
transform 1 0 3196 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_6184
timestamp 1745462530
transform 1 0 3140 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_6185
timestamp 1745462530
transform 1 0 3060 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_6186
timestamp 1745462530
transform 1 0 2892 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_6187
timestamp 1745462530
transform 1 0 2692 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_6188
timestamp 1745462530
transform 1 0 2660 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_6189
timestamp 1745462530
transform 1 0 2612 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_6190
timestamp 1745462530
transform 1 0 3404 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_6191
timestamp 1745462530
transform 1 0 3404 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_6192
timestamp 1745462530
transform 1 0 3372 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_6193
timestamp 1745462530
transform 1 0 3380 0 1 3745
box -2 -2 2 2
use M2_M1  M2_M1_6194
timestamp 1745462530
transform 1 0 3348 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_6195
timestamp 1745462530
transform 1 0 3436 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_6196
timestamp 1745462530
transform 1 0 3412 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_6197
timestamp 1745462530
transform 1 0 3804 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_6198
timestamp 1745462530
transform 1 0 3788 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_6199
timestamp 1745462530
transform 1 0 3764 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_6200
timestamp 1745462530
transform 1 0 3748 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_6201
timestamp 1745462530
transform 1 0 3724 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_6202
timestamp 1745462530
transform 1 0 3596 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_6203
timestamp 1745462530
transform 1 0 3420 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_6204
timestamp 1745462530
transform 1 0 3228 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_6205
timestamp 1745462530
transform 1 0 1796 0 1 3225
box -2 -2 2 2
use M2_M1  M2_M1_6206
timestamp 1745462530
transform 1 0 3676 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_6207
timestamp 1745462530
transform 1 0 3668 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_6208
timestamp 1745462530
transform 1 0 3604 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_6209
timestamp 1745462530
transform 1 0 3588 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_6210
timestamp 1745462530
transform 1 0 3412 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_6211
timestamp 1745462530
transform 1 0 3300 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_6212
timestamp 1745462530
transform 1 0 3300 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_6213
timestamp 1745462530
transform 1 0 3300 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_6214
timestamp 1745462530
transform 1 0 3180 0 1 3225
box -2 -2 2 2
use M2_M1  M2_M1_6215
timestamp 1745462530
transform 1 0 3332 0 1 3315
box -2 -2 2 2
use M2_M1  M2_M1_6216
timestamp 1745462530
transform 1 0 3188 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_6217
timestamp 1745462530
transform 1 0 2372 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_6218
timestamp 1745462530
transform 1 0 2012 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_6219
timestamp 1745462530
transform 1 0 3332 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_6220
timestamp 1745462530
transform 1 0 3284 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_6221
timestamp 1745462530
transform 1 0 3276 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_6222
timestamp 1745462530
transform 1 0 3276 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_6223
timestamp 1745462530
transform 1 0 3268 0 1 3745
box -2 -2 2 2
use M2_M1  M2_M1_6224
timestamp 1745462530
transform 1 0 3372 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_6225
timestamp 1745462530
transform 1 0 3284 0 1 3745
box -2 -2 2 2
use M2_M1  M2_M1_6226
timestamp 1745462530
transform 1 0 3812 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_6227
timestamp 1745462530
transform 1 0 3812 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_6228
timestamp 1745462530
transform 1 0 3764 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_6229
timestamp 1745462530
transform 1 0 3748 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_6230
timestamp 1745462530
transform 1 0 3732 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_6231
timestamp 1745462530
transform 1 0 3732 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_6232
timestamp 1745462530
transform 1 0 3708 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_6233
timestamp 1745462530
transform 1 0 3428 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_6234
timestamp 1745462530
transform 1 0 3356 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_6235
timestamp 1745462530
transform 1 0 3196 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_6236
timestamp 1745462530
transform 1 0 1748 0 1 3315
box -2 -2 2 2
use M2_M1  M2_M1_6237
timestamp 1745462530
transform 1 0 3700 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_6238
timestamp 1745462530
transform 1 0 3660 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_6239
timestamp 1745462530
transform 1 0 3652 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_6240
timestamp 1745462530
transform 1 0 3572 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_6241
timestamp 1745462530
transform 1 0 3436 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_6242
timestamp 1745462530
transform 1 0 3388 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_6243
timestamp 1745462530
transform 1 0 3292 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_6244
timestamp 1745462530
transform 1 0 3236 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_6245
timestamp 1745462530
transform 1 0 3156 0 1 3315
box -2 -2 2 2
use M2_M1  M2_M1_6246
timestamp 1745462530
transform 1 0 3260 0 1 3425
box -2 -2 2 2
use M2_M1  M2_M1_6247
timestamp 1745462530
transform 1 0 3212 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_6248
timestamp 1745462530
transform 1 0 3388 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_6249
timestamp 1745462530
transform 1 0 3340 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_6250
timestamp 1745462530
transform 1 0 3340 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_6251
timestamp 1745462530
transform 1 0 3324 0 1 3595
box -2 -2 2 2
use M2_M1  M2_M1_6252
timestamp 1745462530
transform 1 0 3300 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_6253
timestamp 1745462530
transform 1 0 3372 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_6254
timestamp 1745462530
transform 1 0 3348 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_6255
timestamp 1745462530
transform 1 0 3860 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_6256
timestamp 1745462530
transform 1 0 3844 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_6257
timestamp 1745462530
transform 1 0 3828 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_6258
timestamp 1745462530
transform 1 0 3740 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_6259
timestamp 1745462530
transform 1 0 3644 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_6260
timestamp 1745462530
transform 1 0 3516 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_6261
timestamp 1745462530
transform 1 0 3356 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_6262
timestamp 1745462530
transform 1 0 3172 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_6263
timestamp 1745462530
transform 1 0 1724 0 1 3225
box -2 -2 2 2
use M2_M1  M2_M1_6264
timestamp 1745462530
transform 1 0 3596 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_6265
timestamp 1745462530
transform 1 0 3596 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_6266
timestamp 1745462530
transform 1 0 3540 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_6267
timestamp 1745462530
transform 1 0 3532 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_6268
timestamp 1745462530
transform 1 0 3524 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_6269
timestamp 1745462530
transform 1 0 3396 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_6270
timestamp 1745462530
transform 1 0 3396 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_6271
timestamp 1745462530
transform 1 0 3316 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_6272
timestamp 1745462530
transform 1 0 3276 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_6273
timestamp 1745462530
transform 1 0 3124 0 1 3225
box -2 -2 2 2
use M2_M1  M2_M1_6274
timestamp 1745462530
transform 1 0 3292 0 1 3315
box -2 -2 2 2
use M2_M1  M2_M1_6275
timestamp 1745462530
transform 1 0 3236 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_6276
timestamp 1745462530
transform 1 0 3196 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_6277
timestamp 1745462530
transform 1 0 3164 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_6278
timestamp 1745462530
transform 1 0 3156 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_6279
timestamp 1745462530
transform 1 0 3188 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_6280
timestamp 1745462530
transform 1 0 3156 0 1 3595
box -2 -2 2 2
use M2_M1  M2_M1_6281
timestamp 1745462530
transform 1 0 3172 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_6282
timestamp 1745462530
transform 1 0 3156 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_6283
timestamp 1745462530
transform 1 0 3788 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_6284
timestamp 1745462530
transform 1 0 3772 0 1 3555
box -2 -2 2 2
use M2_M1  M2_M1_6285
timestamp 1745462530
transform 1 0 3740 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_6286
timestamp 1745462530
transform 1 0 3700 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_6287
timestamp 1745462530
transform 1 0 3660 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_6288
timestamp 1745462530
transform 1 0 3156 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_6289
timestamp 1745462530
transform 1 0 3108 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_6290
timestamp 1745462530
transform 1 0 3108 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_6291
timestamp 1745462530
transform 1 0 3084 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_6292
timestamp 1745462530
transform 1 0 1652 0 1 3315
box -2 -2 2 2
use M2_M1  M2_M1_6293
timestamp 1745462530
transform 1 0 3636 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_6294
timestamp 1745462530
transform 1 0 3628 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_6295
timestamp 1745462530
transform 1 0 3580 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_6296
timestamp 1745462530
transform 1 0 3524 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_6297
timestamp 1745462530
transform 1 0 3220 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_6298
timestamp 1745462530
transform 1 0 3212 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_6299
timestamp 1745462530
transform 1 0 3164 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_6300
timestamp 1745462530
transform 1 0 3140 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_6301
timestamp 1745462530
transform 1 0 3092 0 1 3225
box -2 -2 2 2
use M2_M1  M2_M1_6302
timestamp 1745462530
transform 1 0 3180 0 1 3425
box -2 -2 2 2
use M2_M1  M2_M1_6303
timestamp 1745462530
transform 1 0 3132 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_6304
timestamp 1745462530
transform 1 0 2044 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_6305
timestamp 1745462530
transform 1 0 1916 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_6306
timestamp 1745462530
transform 1 0 2420 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_6307
timestamp 1745462530
transform 1 0 2388 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_6308
timestamp 1745462530
transform 1 0 2388 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_6309
timestamp 1745462530
transform 1 0 2420 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_6310
timestamp 1745462530
transform 1 0 2364 0 1 3595
box -2 -2 2 2
use M2_M1  M2_M1_6311
timestamp 1745462530
transform 1 0 2396 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_6312
timestamp 1745462530
transform 1 0 2372 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_6313
timestamp 1745462530
transform 1 0 2460 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_6314
timestamp 1745462530
transform 1 0 2412 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_6315
timestamp 1745462530
transform 1 0 2356 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_6316
timestamp 1745462530
transform 1 0 2340 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_6317
timestamp 1745462530
transform 1 0 2108 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_6318
timestamp 1745462530
transform 1 0 1980 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_6319
timestamp 1745462530
transform 1 0 1908 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_6320
timestamp 1745462530
transform 1 0 1884 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_6321
timestamp 1745462530
transform 1 0 1684 0 1 3225
box -2 -2 2 2
use M2_M1  M2_M1_6322
timestamp 1745462530
transform 1 0 2956 0 1 3225
box -2 -2 2 2
use M2_M1  M2_M1_6323
timestamp 1745462530
transform 1 0 2588 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_6324
timestamp 1745462530
transform 1 0 2500 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_6325
timestamp 1745462530
transform 1 0 2460 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_6326
timestamp 1745462530
transform 1 0 2436 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_6327
timestamp 1745462530
transform 1 0 2436 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_6328
timestamp 1745462530
transform 1 0 2412 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_6329
timestamp 1745462530
transform 1 0 2404 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_6330
timestamp 1745462530
transform 1 0 2364 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_6331
timestamp 1745462530
transform 1 0 2652 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_6332
timestamp 1745462530
transform 1 0 2428 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_6333
timestamp 1745462530
transform 1 0 2260 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_6334
timestamp 1745462530
transform 1 0 1980 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_6335
timestamp 1745462530
transform 1 0 2132 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_6336
timestamp 1745462530
transform 1 0 2108 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_6337
timestamp 1745462530
transform 1 0 2076 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_6338
timestamp 1745462530
transform 1 0 2388 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_6339
timestamp 1745462530
transform 1 0 2100 0 1 3595
box -2 -2 2 2
use M2_M1  M2_M1_6340
timestamp 1745462530
transform 1 0 2164 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_6341
timestamp 1745462530
transform 1 0 2140 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_6342
timestamp 1745462530
transform 1 0 2260 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_6343
timestamp 1745462530
transform 1 0 2236 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_6344
timestamp 1745462530
transform 1 0 2220 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_6345
timestamp 1745462530
transform 1 0 2188 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_6346
timestamp 1745462530
transform 1 0 2148 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_6347
timestamp 1745462530
transform 1 0 1996 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_6348
timestamp 1745462530
transform 1 0 1884 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_6349
timestamp 1745462530
transform 1 0 1804 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_6350
timestamp 1745462530
transform 1 0 1692 0 1 3425
box -2 -2 2 2
use M2_M1  M2_M1_6351
timestamp 1745462530
transform 1 0 2364 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_6352
timestamp 1745462530
transform 1 0 2364 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_6353
timestamp 1745462530
transform 1 0 2348 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_6354
timestamp 1745462530
transform 1 0 2340 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_6355
timestamp 1745462530
transform 1 0 2332 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_6356
timestamp 1745462530
transform 1 0 2316 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_6357
timestamp 1745462530
transform 1 0 2316 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_6358
timestamp 1745462530
transform 1 0 2276 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_6359
timestamp 1745462530
transform 1 0 2276 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_6360
timestamp 1745462530
transform 1 0 2236 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_6361
timestamp 1745462530
transform 1 0 2604 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_6362
timestamp 1745462530
transform 1 0 2380 0 1 3425
box -2 -2 2 2
use M2_M1  M2_M1_6363
timestamp 1745462530
transform 1 0 2892 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_6364
timestamp 1745462530
transform 1 0 2876 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_6365
timestamp 1745462530
transform 1 0 2844 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_6366
timestamp 1745462530
transform 1 0 2860 0 1 3595
box -2 -2 2 2
use M2_M1  M2_M1_6367
timestamp 1745462530
transform 1 0 2860 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_6368
timestamp 1745462530
transform 1 0 2876 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_6369
timestamp 1745462530
transform 1 0 2860 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_6370
timestamp 1745462530
transform 1 0 3604 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_6371
timestamp 1745462530
transform 1 0 3524 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_6372
timestamp 1745462530
transform 1 0 3428 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_6373
timestamp 1745462530
transform 1 0 3124 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_6374
timestamp 1745462530
transform 1 0 3052 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_6375
timestamp 1745462530
transform 1 0 2820 0 1 3635
box -2 -2 2 2
use M2_M1  M2_M1_6376
timestamp 1745462530
transform 1 0 2404 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_6377
timestamp 1745462530
transform 1 0 2276 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_6378
timestamp 1745462530
transform 1 0 1900 0 1 3515
box -2 -2 2 2
use M2_M1  M2_M1_6379
timestamp 1745462530
transform 1 0 2836 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_6380
timestamp 1745462530
transform 1 0 2764 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_6381
timestamp 1745462530
transform 1 0 2764 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_6382
timestamp 1745462530
transform 1 0 2724 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_6383
timestamp 1745462530
transform 1 0 2708 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_6384
timestamp 1745462530
transform 1 0 2604 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_6385
timestamp 1745462530
transform 1 0 1956 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_6386
timestamp 1745462530
transform 1 0 1772 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_6387
timestamp 1745462530
transform 1 0 1756 0 1 3225
box -2 -2 2 2
use M2_M1  M2_M1_6388
timestamp 1745462530
transform 1 0 3428 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_6389
timestamp 1745462530
transform 1 0 3396 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_6390
timestamp 1745462530
transform 1 0 3388 0 1 3595
box -2 -2 2 2
use M2_M1  M2_M1_6391
timestamp 1745462530
transform 1 0 3148 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_6392
timestamp 1745462530
transform 1 0 3060 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_6393
timestamp 1745462530
transform 1 0 2836 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_6394
timestamp 1745462530
transform 1 0 2508 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_6395
timestamp 1745462530
transform 1 0 2316 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_6396
timestamp 1745462530
transform 1 0 2308 0 1 3425
box -2 -2 2 2
use M2_M1  M2_M1_6397
timestamp 1745462530
transform 1 0 3020 0 1 3225
box -2 -2 2 2
use M2_M1  M2_M1_6398
timestamp 1745462530
transform 1 0 2844 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_6399
timestamp 1745462530
transform 1 0 2836 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_6400
timestamp 1745462530
transform 1 0 2740 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_6401
timestamp 1745462530
transform 1 0 2708 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_6402
timestamp 1745462530
transform 1 0 2684 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_6403
timestamp 1745462530
transform 1 0 2684 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_6404
timestamp 1745462530
transform 1 0 2652 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_6405
timestamp 1745462530
transform 1 0 2636 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_6406
timestamp 1745462530
transform 1 0 2604 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_6407
timestamp 1745462530
transform 1 0 2892 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_6408
timestamp 1745462530
transform 1 0 2868 0 1 3495
box -2 -2 2 2
use M2_M1  M2_M1_6409
timestamp 1745462530
transform 1 0 3412 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_6410
timestamp 1745462530
transform 1 0 3388 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_6411
timestamp 1745462530
transform 1 0 3364 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_6412
timestamp 1745462530
transform 1 0 3132 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_6413
timestamp 1745462530
transform 1 0 3084 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_6414
timestamp 1745462530
transform 1 0 2908 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_6415
timestamp 1745462530
transform 1 0 2572 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_6416
timestamp 1745462530
transform 1 0 2540 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_6417
timestamp 1745462530
transform 1 0 2532 0 1 3505
box -2 -2 2 2
use M2_M1  M2_M1_6418
timestamp 1745462530
transform 1 0 2484 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_6419
timestamp 1745462530
transform 1 0 3124 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_6420
timestamp 1745462530
transform 1 0 3100 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_6421
timestamp 1745462530
transform 1 0 3092 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_6422
timestamp 1745462530
transform 1 0 3092 0 1 3745
box -2 -2 2 2
use M2_M1  M2_M1_6423
timestamp 1745462530
transform 1 0 3084 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_6424
timestamp 1745462530
transform 1 0 3108 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_6425
timestamp 1745462530
transform 1 0 3092 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_6426
timestamp 1745462530
transform 1 0 3076 0 1 3625
box -2 -2 2 2
use M2_M1  M2_M1_6427
timestamp 1745462530
transform 1 0 3068 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_6428
timestamp 1745462530
transform 1 0 3652 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_6429
timestamp 1745462530
transform 1 0 3636 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_6430
timestamp 1745462530
transform 1 0 3612 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_6431
timestamp 1745462530
transform 1 0 3628 0 1 3595
box -2 -2 2 2
use M2_M1  M2_M1_6432
timestamp 1745462530
transform 1 0 3460 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_6433
timestamp 1745462530
transform 1 0 3644 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_6434
timestamp 1745462530
transform 1 0 3628 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_6435
timestamp 1745462530
transform 1 0 3444 0 1 3515
box -2 -2 2 2
use M2_M1  M2_M1_6436
timestamp 1745462530
transform 1 0 3348 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_6437
timestamp 1745462530
transform 1 0 3636 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_6438
timestamp 1745462530
transform 1 0 3588 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_6439
timestamp 1745462530
transform 1 0 3492 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_6440
timestamp 1745462530
transform 1 0 3460 0 1 3595
box -2 -2 2 2
use M2_M1  M2_M1_6441
timestamp 1745462530
transform 1 0 3420 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_6442
timestamp 1745462530
transform 1 0 3476 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_6443
timestamp 1745462530
transform 1 0 3460 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_6444
timestamp 1745462530
transform 1 0 3420 0 1 3625
box -2 -2 2 2
use M2_M1  M2_M1_6445
timestamp 1745462530
transform 1 0 3396 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_6446
timestamp 1745462530
transform 1 0 3628 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_6447
timestamp 1745462530
transform 1 0 3596 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_6448
timestamp 1745462530
transform 1 0 3508 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_6449
timestamp 1745462530
transform 1 0 3476 0 1 3595
box -2 -2 2 2
use M2_M1  M2_M1_6450
timestamp 1745462530
transform 1 0 3420 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_6451
timestamp 1745462530
transform 1 0 3540 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_6452
timestamp 1745462530
transform 1 0 3516 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_6453
timestamp 1745462530
transform 1 0 3420 0 1 3425
box -2 -2 2 2
use M2_M1  M2_M1_6454
timestamp 1745462530
transform 1 0 3372 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_6455
timestamp 1745462530
transform 1 0 3268 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_6456
timestamp 1745462530
transform 1 0 3228 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_6457
timestamp 1745462530
transform 1 0 3196 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_6458
timestamp 1745462530
transform 1 0 3180 0 1 3795
box -2 -2 2 2
use M2_M1  M2_M1_6459
timestamp 1745462530
transform 1 0 3164 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_6460
timestamp 1745462530
transform 1 0 3204 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_6461
timestamp 1745462530
transform 1 0 3148 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_6462
timestamp 1745462530
transform 1 0 3172 0 1 3515
box -2 -2 2 2
use M2_M1  M2_M1_6463
timestamp 1745462530
transform 1 0 3116 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_6464
timestamp 1745462530
transform 1 0 2436 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_6465
timestamp 1745462530
transform 1 0 2412 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_6466
timestamp 1745462530
transform 1 0 2380 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_6467
timestamp 1745462530
transform 1 0 2540 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_6468
timestamp 1745462530
transform 1 0 2436 0 1 3795
box -2 -2 2 2
use M2_M1  M2_M1_6469
timestamp 1745462530
transform 1 0 2452 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_6470
timestamp 1745462530
transform 1 0 2452 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_6471
timestamp 1745462530
transform 1 0 2532 0 1 3625
box -2 -2 2 2
use M2_M1  M2_M1_6472
timestamp 1745462530
transform 1 0 2508 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_6473
timestamp 1745462530
transform 1 0 2348 0 1 3755
box -2 -2 2 2
use M2_M1  M2_M1_6474
timestamp 1745462530
transform 1 0 2252 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_6475
timestamp 1745462530
transform 1 0 2212 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_6476
timestamp 1745462530
transform 1 0 2356 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_6477
timestamp 1745462530
transform 1 0 2324 0 1 3745
box -2 -2 2 2
use M2_M1  M2_M1_6478
timestamp 1745462530
transform 1 0 2340 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_6479
timestamp 1745462530
transform 1 0 2324 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_6480
timestamp 1745462530
transform 1 0 1852 0 1 3505
box -2 -2 2 2
use M2_M1  M2_M1_6481
timestamp 1745462530
transform 1 0 1852 0 1 3435
box -2 -2 2 2
use M2_M1  M2_M1_6482
timestamp 1745462530
transform 1 0 2452 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_6483
timestamp 1745462530
transform 1 0 2372 0 1 3515
box -2 -2 2 2
use M2_M1  M2_M1_6484
timestamp 1745462530
transform 1 0 2116 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_6485
timestamp 1745462530
transform 1 0 1900 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_6486
timestamp 1745462530
transform 1 0 2652 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_6487
timestamp 1745462530
transform 1 0 2644 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_6488
timestamp 1745462530
transform 1 0 2628 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_6489
timestamp 1745462530
transform 1 0 2588 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_6490
timestamp 1745462530
transform 1 0 2556 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_6491
timestamp 1745462530
transform 1 0 2548 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_6492
timestamp 1745462530
transform 1 0 2396 0 1 3825
box -2 -2 2 2
use M2_M1  M2_M1_6493
timestamp 1745462530
transform 1 0 1876 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_6494
timestamp 1745462530
transform 1 0 1780 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_6495
timestamp 1745462530
transform 1 0 1628 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_6496
timestamp 1745462530
transform 1 0 2500 0 1 3025
box -2 -2 2 2
use M2_M1  M2_M1_6497
timestamp 1745462530
transform 1 0 2476 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_6498
timestamp 1745462530
transform 1 0 2604 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_6499
timestamp 1745462530
transform 1 0 2596 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_6500
timestamp 1745462530
transform 1 0 2580 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_6501
timestamp 1745462530
transform 1 0 2476 0 1 3025
box -2 -2 2 2
use M2_M1  M2_M1_6502
timestamp 1745462530
transform 1 0 2412 0 1 2995
box -2 -2 2 2
use M2_M1  M2_M1_6503
timestamp 1745462530
transform 1 0 2412 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_6504
timestamp 1745462530
transform 1 0 2548 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_6505
timestamp 1745462530
transform 1 0 2508 0 1 2995
box -2 -2 2 2
use M2_M1  M2_M1_6506
timestamp 1745462530
transform 1 0 2484 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_6507
timestamp 1745462530
transform 1 0 2396 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_6508
timestamp 1745462530
transform 1 0 2372 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_6509
timestamp 1745462530
transform 1 0 2476 0 1 3035
box -2 -2 2 2
use M2_M1  M2_M1_6510
timestamp 1745462530
transform 1 0 2460 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_6511
timestamp 1745462530
transform 1 0 2620 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_6512
timestamp 1745462530
transform 1 0 2612 0 1 3025
box -2 -2 2 2
use M2_M1  M2_M1_6513
timestamp 1745462530
transform 1 0 2572 0 1 3025
box -2 -2 2 2
use M2_M1  M2_M1_6514
timestamp 1745462530
transform 1 0 2428 0 1 2995
box -2 -2 2 2
use M2_M1  M2_M1_6515
timestamp 1745462530
transform 1 0 2364 0 1 3025
box -2 -2 2 2
use M2_M1  M2_M1_6516
timestamp 1745462530
transform 1 0 2284 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_6517
timestamp 1745462530
transform 1 0 2260 0 1 3435
box -2 -2 2 2
use M2_M1  M2_M1_6518
timestamp 1745462530
transform 1 0 2260 0 1 3305
box -2 -2 2 2
use M2_M1  M2_M1_6519
timestamp 1745462530
transform 1 0 2140 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_6520
timestamp 1745462530
transform 1 0 2756 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_6521
timestamp 1745462530
transform 1 0 2748 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_6522
timestamp 1745462530
transform 1 0 2724 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_6523
timestamp 1745462530
transform 1 0 2772 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_6524
timestamp 1745462530
transform 1 0 2748 0 1 3595
box -2 -2 2 2
use M2_M1  M2_M1_6525
timestamp 1745462530
transform 1 0 2796 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_6526
timestamp 1745462530
transform 1 0 2772 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_6527
timestamp 1745462530
transform 1 0 3236 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_6528
timestamp 1745462530
transform 1 0 3188 0 1 3715
box -2 -2 2 2
use M2_M1  M2_M1_6529
timestamp 1745462530
transform 1 0 3180 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_6530
timestamp 1745462530
transform 1 0 3156 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_6531
timestamp 1745462530
transform 1 0 2996 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_6532
timestamp 1745462530
transform 1 0 2780 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_6533
timestamp 1745462530
transform 1 0 2364 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_6534
timestamp 1745462530
transform 1 0 2228 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_6535
timestamp 1745462530
transform 1 0 1852 0 1 3625
box -2 -2 2 2
use M2_M1  M2_M1_6536
timestamp 1745462530
transform 1 0 3316 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_6537
timestamp 1745462530
transform 1 0 3308 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_6538
timestamp 1745462530
transform 1 0 3300 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_6539
timestamp 1745462530
transform 1 0 3220 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_6540
timestamp 1745462530
transform 1 0 3004 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_6541
timestamp 1745462530
transform 1 0 2756 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_6542
timestamp 1745462530
transform 1 0 2404 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_6543
timestamp 1745462530
transform 1 0 2244 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_6544
timestamp 1745462530
transform 1 0 2244 0 1 3425
box -2 -2 2 2
use M2_M1  M2_M1_6545
timestamp 1745462530
transform 1 0 2804 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_6546
timestamp 1745462530
transform 1 0 2780 0 1 3515
box -2 -2 2 2
use M2_M1  M2_M1_6547
timestamp 1745462530
transform 1 0 3308 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_6548
timestamp 1745462530
transform 1 0 3292 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_6549
timestamp 1745462530
transform 1 0 3284 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_6550
timestamp 1745462530
transform 1 0 3212 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_6551
timestamp 1745462530
transform 1 0 3036 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_6552
timestamp 1745462530
transform 1 0 2828 0 1 3545
box -2 -2 2 2
use M2_M1  M2_M1_6553
timestamp 1745462530
transform 1 0 2564 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_6554
timestamp 1745462530
transform 1 0 2492 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_6555
timestamp 1745462530
transform 1 0 2428 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_6556
timestamp 1745462530
transform 1 0 3052 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_6557
timestamp 1745462530
transform 1 0 3052 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_6558
timestamp 1745462530
transform 1 0 3020 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_6559
timestamp 1745462530
transform 1 0 3044 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_6560
timestamp 1745462530
transform 1 0 3020 0 1 3745
box -2 -2 2 2
use M2_M1  M2_M1_6561
timestamp 1745462530
transform 1 0 3036 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_6562
timestamp 1745462530
transform 1 0 3020 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_6563
timestamp 1745462530
transform 1 0 3028 0 1 3625
box -2 -2 2 2
use M2_M1  M2_M1_6564
timestamp 1745462530
transform 1 0 3020 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_6565
timestamp 1745462530
transform 1 0 3492 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_6566
timestamp 1745462530
transform 1 0 3468 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_6567
timestamp 1745462530
transform 1 0 3340 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_6568
timestamp 1745462530
transform 1 0 3324 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_6569
timestamp 1745462530
transform 1 0 3316 0 1 3745
box -2 -2 2 2
use M2_M1  M2_M1_6570
timestamp 1745462530
transform 1 0 3340 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_6571
timestamp 1745462530
transform 1 0 3260 0 1 3715
box -2 -2 2 2
use M2_M1  M2_M1_6572
timestamp 1745462530
transform 1 0 3324 0 1 3515
box -2 -2 2 2
use M2_M1  M2_M1_6573
timestamp 1745462530
transform 1 0 3276 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_6574
timestamp 1745462530
transform 1 0 3388 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_6575
timestamp 1745462530
transform 1 0 3364 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_6576
timestamp 1745462530
transform 1 0 3324 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_6577
timestamp 1745462530
transform 1 0 3324 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_6578
timestamp 1745462530
transform 1 0 3292 0 1 3745
box -2 -2 2 2
use M2_M1  M2_M1_6579
timestamp 1745462530
transform 1 0 3308 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_6580
timestamp 1745462530
transform 1 0 3228 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_6581
timestamp 1745462530
transform 1 0 3316 0 1 3625
box -2 -2 2 2
use M2_M1  M2_M1_6582
timestamp 1745462530
transform 1 0 3268 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_6583
timestamp 1745462530
transform 1 0 3508 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_6584
timestamp 1745462530
transform 1 0 3476 0 1 4005
box -2 -2 2 2
use M2_M1  M2_M1_6585
timestamp 1745462530
transform 1 0 3212 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_6586
timestamp 1745462530
transform 1 0 3340 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_6587
timestamp 1745462530
transform 1 0 3212 0 1 3595
box -2 -2 2 2
use M2_M1  M2_M1_6588
timestamp 1745462530
transform 1 0 3228 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_6589
timestamp 1745462530
transform 1 0 3204 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_6590
timestamp 1745462530
transform 1 0 3340 0 1 3425
box -2 -2 2 2
use M2_M1  M2_M1_6591
timestamp 1745462530
transform 1 0 3292 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_6592
timestamp 1745462530
transform 1 0 3212 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_6593
timestamp 1745462530
transform 1 0 3212 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_6594
timestamp 1745462530
transform 1 0 3180 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_6595
timestamp 1745462530
transform 1 0 3244 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_6596
timestamp 1745462530
transform 1 0 3212 0 1 3795
box -2 -2 2 2
use M2_M1  M2_M1_6597
timestamp 1745462530
transform 1 0 3228 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_6598
timestamp 1745462530
transform 1 0 3188 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_6599
timestamp 1745462530
transform 1 0 3244 0 1 3515
box -2 -2 2 2
use M2_M1  M2_M1_6600
timestamp 1745462530
transform 1 0 3196 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_6601
timestamp 1745462530
transform 1 0 2444 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_6602
timestamp 1745462530
transform 1 0 2412 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_6603
timestamp 1745462530
transform 1 0 2412 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_6604
timestamp 1745462530
transform 1 0 2436 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_6605
timestamp 1745462530
transform 1 0 2404 0 1 3795
box -2 -2 2 2
use M2_M1  M2_M1_6606
timestamp 1745462530
transform 1 0 2420 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_6607
timestamp 1745462530
transform 1 0 2404 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_6608
timestamp 1745462530
transform 1 0 2476 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_6609
timestamp 1745462530
transform 1 0 2452 0 1 3625
box -2 -2 2 2
use M2_M1  M2_M1_6610
timestamp 1745462530
transform 1 0 2212 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_6611
timestamp 1745462530
transform 1 0 2204 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_6612
timestamp 1745462530
transform 1 0 2180 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_6613
timestamp 1745462530
transform 1 0 2268 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_6614
timestamp 1745462530
transform 1 0 2188 0 1 3745
box -2 -2 2 2
use M2_M1  M2_M1_6615
timestamp 1745462530
transform 1 0 2244 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_6616
timestamp 1745462530
transform 1 0 2220 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_6617
timestamp 1745462530
transform 1 0 1812 0 1 3435
box -2 -2 2 2
use M2_M1  M2_M1_6618
timestamp 1745462530
transform 1 0 1804 0 1 3635
box -2 -2 2 2
use M2_M1  M2_M1_6619
timestamp 1745462530
transform 1 0 1748 0 1 3635
box -2 -2 2 2
use M2_M1  M2_M1_6620
timestamp 1745462530
transform 1 0 1740 0 1 3435
box -2 -2 2 2
use M2_M1  M2_M1_6621
timestamp 1745462530
transform 1 0 2404 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_6622
timestamp 1745462530
transform 1 0 2276 0 1 3515
box -2 -2 2 2
use M2_M1  M2_M1_6623
timestamp 1745462530
transform 1 0 2148 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_6624
timestamp 1745462530
transform 1 0 1812 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_6625
timestamp 1745462530
transform 1 0 2396 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_6626
timestamp 1745462530
transform 1 0 2388 0 1 3025
box -2 -2 2 2
use M2_M1  M2_M1_6627
timestamp 1745462530
transform 1 0 2412 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_6628
timestamp 1745462530
transform 1 0 2380 0 1 3035
box -2 -2 2 2
use M2_M1  M2_M1_6629
timestamp 1745462530
transform 1 0 2188 0 1 3825
box -2 -2 2 2
use M2_M1  M2_M1_6630
timestamp 1745462530
transform 1 0 2180 0 1 3395
box -2 -2 2 2
use M2_M1  M2_M1_6631
timestamp 1745462530
transform 1 0 2148 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_6632
timestamp 1745462530
transform 1 0 2140 0 1 3345
box -2 -2 2 2
use M2_M1  M2_M1_6633
timestamp 1745462530
transform 1 0 2100 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_6634
timestamp 1745462530
transform 1 0 2100 0 1 3395
box -2 -2 2 2
use M2_M1  M2_M1_6635
timestamp 1745462530
transform 1 0 2044 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_6636
timestamp 1745462530
transform 1 0 1836 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_6637
timestamp 1745462530
transform 1 0 1764 0 1 3545
box -2 -2 2 2
use M2_M1  M2_M1_6638
timestamp 1745462530
transform 1 0 1716 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_6639
timestamp 1745462530
transform 1 0 1692 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_6640
timestamp 1745462530
transform 1 0 1116 0 1 3315
box -2 -2 2 2
use M2_M1  M2_M1_6641
timestamp 1745462530
transform 1 0 1116 0 1 3225
box -2 -2 2 2
use M2_M1  M2_M1_6642
timestamp 1745462530
transform 1 0 2708 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_6643
timestamp 1745462530
transform 1 0 2692 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_6644
timestamp 1745462530
transform 1 0 2652 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_6645
timestamp 1745462530
transform 1 0 2700 0 1 3745
box -2 -2 2 2
use M2_M1  M2_M1_6646
timestamp 1745462530
transform 1 0 2684 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_6647
timestamp 1745462530
transform 1 0 2764 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_6648
timestamp 1745462530
transform 1 0 2740 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_6649
timestamp 1745462530
transform 1 0 3748 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_6650
timestamp 1745462530
transform 1 0 3724 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_6651
timestamp 1745462530
transform 1 0 3724 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_6652
timestamp 1745462530
transform 1 0 3668 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_6653
timestamp 1745462530
transform 1 0 2932 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_6654
timestamp 1745462530
transform 1 0 2748 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_6655
timestamp 1745462530
transform 1 0 2468 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_6656
timestamp 1745462530
transform 1 0 2260 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_6657
timestamp 1745462530
transform 1 0 1756 0 1 3625
box -2 -2 2 2
use M2_M1  M2_M1_6658
timestamp 1745462530
transform 1 0 3668 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_6659
timestamp 1745462530
transform 1 0 3660 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_6660
timestamp 1745462530
transform 1 0 3644 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_6661
timestamp 1745462530
transform 1 0 3620 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_6662
timestamp 1745462530
transform 1 0 3604 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_6663
timestamp 1745462530
transform 1 0 2940 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_6664
timestamp 1745462530
transform 1 0 2636 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_6665
timestamp 1745462530
transform 1 0 2596 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_6666
timestamp 1745462530
transform 1 0 2580 0 1 3625
box -2 -2 2 2
use M2_M1  M2_M1_6667
timestamp 1745462530
transform 1 0 2292 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_6668
timestamp 1745462530
transform 1 0 2172 0 1 3515
box -2 -2 2 2
use M2_M1  M2_M1_6669
timestamp 1745462530
transform 1 0 2708 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_6670
timestamp 1745462530
transform 1 0 2684 0 1 3515
box -2 -2 2 2
use M2_M1  M2_M1_6671
timestamp 1745462530
transform 1 0 3588 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_6672
timestamp 1745462530
transform 1 0 3580 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_6673
timestamp 1745462530
transform 1 0 3532 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_6674
timestamp 1745462530
transform 1 0 3492 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_6675
timestamp 1745462530
transform 1 0 2996 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_6676
timestamp 1745462530
transform 1 0 2724 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_6677
timestamp 1745462530
transform 1 0 2660 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_6678
timestamp 1745462530
transform 1 0 2636 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_6679
timestamp 1745462530
transform 1 0 2580 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_6680
timestamp 1745462530
transform 1 0 2988 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_6681
timestamp 1745462530
transform 1 0 2972 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_6682
timestamp 1745462530
transform 1 0 2964 0 1 4005
box -2 -2 2 2
use M2_M1  M2_M1_6683
timestamp 1745462530
transform 1 0 2964 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_6684
timestamp 1745462530
transform 1 0 2956 0 1 3745
box -2 -2 2 2
use M2_M1  M2_M1_6685
timestamp 1745462530
transform 1 0 2972 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_6686
timestamp 1745462530
transform 1 0 2956 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_6687
timestamp 1745462530
transform 1 0 2980 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_6688
timestamp 1745462530
transform 1 0 2956 0 1 3515
box -2 -2 2 2
use M2_M1  M2_M1_6689
timestamp 1745462530
transform 1 0 3764 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_6690
timestamp 1745462530
transform 1 0 3740 0 1 4005
box -2 -2 2 2
use M2_M1  M2_M1_6691
timestamp 1745462530
transform 1 0 3708 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_6692
timestamp 1745462530
transform 1 0 3700 0 1 3595
box -2 -2 2 2
use M2_M1  M2_M1_6693
timestamp 1745462530
transform 1 0 3700 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_6694
timestamp 1745462530
transform 1 0 3748 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_6695
timestamp 1745462530
transform 1 0 3716 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_6696
timestamp 1745462530
transform 1 0 3700 0 1 3515
box -2 -2 2 2
use M2_M1  M2_M1_6697
timestamp 1745462530
transform 1 0 3564 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_6698
timestamp 1745462530
transform 1 0 3892 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_6699
timestamp 1745462530
transform 1 0 3860 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_6700
timestamp 1745462530
transform 1 0 3796 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_6701
timestamp 1745462530
transform 1 0 3764 0 1 3745
box -2 -2 2 2
use M2_M1  M2_M1_6702
timestamp 1745462530
transform 1 0 3700 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_6703
timestamp 1745462530
transform 1 0 3780 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_6704
timestamp 1745462530
transform 1 0 3764 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_6705
timestamp 1745462530
transform 1 0 3684 0 1 3625
box -2 -2 2 2
use M2_M1  M2_M1_6706
timestamp 1745462530
transform 1 0 3572 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_6707
timestamp 1745462530
transform 1 0 3724 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_6708
timestamp 1745462530
transform 1 0 3684 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_6709
timestamp 1745462530
transform 1 0 3668 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_6710
timestamp 1745462530
transform 1 0 3708 0 1 3545
box -2 -2 2 2
use M2_M1  M2_M1_6711
timestamp 1745462530
transform 1 0 3628 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_6712
timestamp 1745462530
transform 1 0 3772 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_6713
timestamp 1745462530
transform 1 0 3732 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_6714
timestamp 1745462530
transform 1 0 3620 0 1 3515
box -2 -2 2 2
use M2_M1  M2_M1_6715
timestamp 1745462530
transform 1 0 3516 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_6716
timestamp 1745462530
transform 1 0 3716 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_6717
timestamp 1745462530
transform 1 0 3700 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_6718
timestamp 1745462530
transform 1 0 3692 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_6719
timestamp 1745462530
transform 1 0 3692 0 1 3745
box -2 -2 2 2
use M2_M1  M2_M1_6720
timestamp 1745462530
transform 1 0 3668 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_6721
timestamp 1745462530
transform 1 0 3708 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_6722
timestamp 1745462530
transform 1 0 3692 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_6723
timestamp 1745462530
transform 1 0 3660 0 1 3515
box -2 -2 2 2
use M2_M1  M2_M1_6724
timestamp 1745462530
transform 1 0 3476 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_6725
timestamp 1745462530
transform 1 0 2524 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_6726
timestamp 1745462530
transform 1 0 2516 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_6727
timestamp 1745462530
transform 1 0 2492 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_6728
timestamp 1745462530
transform 1 0 2612 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_6729
timestamp 1745462530
transform 1 0 2500 0 1 3745
box -2 -2 2 2
use M2_M1  M2_M1_6730
timestamp 1745462530
transform 1 0 2524 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_6731
timestamp 1745462530
transform 1 0 2508 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_6732
timestamp 1745462530
transform 1 0 2620 0 1 3595
box -2 -2 2 2
use M2_M1  M2_M1_6733
timestamp 1745462530
transform 1 0 2620 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_6734
timestamp 1745462530
transform 1 0 2324 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_6735
timestamp 1745462530
transform 1 0 2316 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_6736
timestamp 1745462530
transform 1 0 2292 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_6737
timestamp 1745462530
transform 1 0 2316 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_6738
timestamp 1745462530
transform 1 0 2284 0 1 3595
box -2 -2 2 2
use M2_M1  M2_M1_6739
timestamp 1745462530
transform 1 0 2308 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_6740
timestamp 1745462530
transform 1 0 2284 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_6741
timestamp 1745462530
transform 1 0 2564 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_6742
timestamp 1745462530
transform 1 0 2324 0 1 3515
box -2 -2 2 2
use M2_M1  M2_M1_6743
timestamp 1745462530
transform 1 0 2684 0 1 3105
box -2 -2 2 2
use M2_M1  M2_M1_6744
timestamp 1745462530
transform 1 0 2684 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_6745
timestamp 1745462530
transform 1 0 2628 0 1 3035
box -2 -2 2 2
use M2_M1  M2_M1_6746
timestamp 1745462530
transform 1 0 2684 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_6747
timestamp 1745462530
transform 1 0 2636 0 1 4005
box -2 -2 2 2
use M2_M1  M2_M1_6748
timestamp 1745462530
transform 1 0 2596 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_6749
timestamp 1745462530
transform 1 0 2708 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_6750
timestamp 1745462530
transform 1 0 2668 0 1 3595
box -2 -2 2 2
use M2_M1  M2_M1_6751
timestamp 1745462530
transform 1 0 2748 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_6752
timestamp 1745462530
transform 1 0 2708 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_6753
timestamp 1745462530
transform 1 0 3852 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_6754
timestamp 1745462530
transform 1 0 3804 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_6755
timestamp 1745462530
transform 1 0 3780 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_6756
timestamp 1745462530
transform 1 0 3780 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_6757
timestamp 1745462530
transform 1 0 2884 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_6758
timestamp 1745462530
transform 1 0 2716 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_6759
timestamp 1745462530
transform 1 0 2004 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_6760
timestamp 1745462530
transform 1 0 1884 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_6761
timestamp 1745462530
transform 1 0 1812 0 1 3515
box -2 -2 2 2
use M2_M1  M2_M1_6762
timestamp 1745462530
transform 1 0 3708 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_6763
timestamp 1745462530
transform 1 0 3676 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_6764
timestamp 1745462530
transform 1 0 3636 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_6765
timestamp 1745462530
transform 1 0 3604 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_6766
timestamp 1745462530
transform 1 0 2940 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_6767
timestamp 1745462530
transform 1 0 2692 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_6768
timestamp 1745462530
transform 1 0 2444 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_6769
timestamp 1745462530
transform 1 0 2324 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_6770
timestamp 1745462530
transform 1 0 2300 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_6771
timestamp 1745462530
transform 1 0 2180 0 1 3425
box -2 -2 2 2
use M2_M1  M2_M1_6772
timestamp 1745462530
transform 1 0 2740 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_6773
timestamp 1745462530
transform 1 0 2716 0 1 3425
box -2 -2 2 2
use M2_M1  M2_M1_6774
timestamp 1745462530
transform 1 0 3588 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_6775
timestamp 1745462530
transform 1 0 3548 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_6776
timestamp 1745462530
transform 1 0 3508 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_6777
timestamp 1745462530
transform 1 0 3460 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_6778
timestamp 1745462530
transform 1 0 2924 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_6779
timestamp 1745462530
transform 1 0 2756 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_6780
timestamp 1745462530
transform 1 0 2604 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_6781
timestamp 1745462530
transform 1 0 2564 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_6782
timestamp 1745462530
transform 1 0 2524 0 1 3425
box -2 -2 2 2
use M2_M1  M2_M1_6783
timestamp 1745462530
transform 1 0 2956 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_6784
timestamp 1745462530
transform 1 0 2956 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_6785
timestamp 1745462530
transform 1 0 2924 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_6786
timestamp 1745462530
transform 1 0 2956 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_6787
timestamp 1745462530
transform 1 0 2932 0 1 3595
box -2 -2 2 2
use M2_M1  M2_M1_6788
timestamp 1745462530
transform 1 0 2948 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_6789
timestamp 1745462530
transform 1 0 2932 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_6790
timestamp 1745462530
transform 1 0 2956 0 1 3425
box -2 -2 2 2
use M2_M1  M2_M1_6791
timestamp 1745462530
transform 1 0 2908 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_6792
timestamp 1745462530
transform 1 0 4300 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_6793
timestamp 1745462530
transform 1 0 4284 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_6794
timestamp 1745462530
transform 1 0 4268 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_6795
timestamp 1745462530
transform 1 0 3876 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_6796
timestamp 1745462530
transform 1 0 3844 0 1 3595
box -2 -2 2 2
use M2_M1  M2_M1_6797
timestamp 1745462530
transform 1 0 3700 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_6798
timestamp 1745462530
transform 1 0 3868 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_6799
timestamp 1745462530
transform 1 0 3852 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_6800
timestamp 1745462530
transform 1 0 3692 0 1 3425
box -2 -2 2 2
use M2_M1  M2_M1_6801
timestamp 1745462530
transform 1 0 3532 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_6802
timestamp 1745462530
transform 1 0 4212 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_6803
timestamp 1745462530
transform 1 0 4196 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_6804
timestamp 1745462530
transform 1 0 3900 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_6805
timestamp 1745462530
transform 1 0 3876 0 1 3595
box -2 -2 2 2
use M2_M1  M2_M1_6806
timestamp 1745462530
transform 1 0 3732 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_6807
timestamp 1745462530
transform 1 0 3892 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_6808
timestamp 1745462530
transform 1 0 3796 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_6809
timestamp 1745462530
transform 1 0 3724 0 1 3425
box -2 -2 2 2
use M2_M1  M2_M1_6810
timestamp 1745462530
transform 1 0 3572 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_6811
timestamp 1745462530
transform 1 0 4228 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_6812
timestamp 1745462530
transform 1 0 4204 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_6813
timestamp 1745462530
transform 1 0 3900 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_6814
timestamp 1745462530
transform 1 0 3892 0 1 3545
box -2 -2 2 2
use M2_M1  M2_M1_6815
timestamp 1745462530
transform 1 0 3620 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_6816
timestamp 1745462530
transform 1 0 3908 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_6817
timestamp 1745462530
transform 1 0 3892 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_6818
timestamp 1745462530
transform 1 0 3620 0 1 3425
box -2 -2 2 2
use M2_M1  M2_M1_6819
timestamp 1745462530
transform 1 0 3492 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_6820
timestamp 1745462530
transform 1 0 3964 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_6821
timestamp 1745462530
transform 1 0 3908 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_6822
timestamp 1745462530
transform 1 0 3852 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_6823
timestamp 1745462530
transform 1 0 3820 0 1 3545
box -2 -2 2 2
use M2_M1  M2_M1_6824
timestamp 1745462530
transform 1 0 3652 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_6825
timestamp 1745462530
transform 1 0 3836 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_6826
timestamp 1745462530
transform 1 0 3820 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_6827
timestamp 1745462530
transform 1 0 3660 0 1 3425
box -2 -2 2 2
use M2_M1  M2_M1_6828
timestamp 1745462530
transform 1 0 3444 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_6829
timestamp 1745462530
transform 1 0 1988 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_6830
timestamp 1745462530
transform 1 0 1980 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_6831
timestamp 1745462530
transform 1 0 1964 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_6832
timestamp 1745462530
transform 1 0 2460 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_6833
timestamp 1745462530
transform 1 0 1956 0 1 3545
box -2 -2 2 2
use M2_M1  M2_M1_6834
timestamp 1745462530
transform 1 0 1972 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_6835
timestamp 1745462530
transform 1 0 1948 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_6836
timestamp 1745462530
transform 1 0 2500 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_6837
timestamp 1745462530
transform 1 0 2476 0 1 3425
box -2 -2 2 2
use M2_M1  M2_M1_6838
timestamp 1745462530
transform 1 0 2060 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_6839
timestamp 1745462530
transform 1 0 2020 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_6840
timestamp 1745462530
transform 1 0 1996 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_6841
timestamp 1745462530
transform 1 0 2340 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_6842
timestamp 1745462530
transform 1 0 2044 0 1 3545
box -2 -2 2 2
use M2_M1  M2_M1_6843
timestamp 1745462530
transform 1 0 2068 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_6844
timestamp 1745462530
transform 1 0 2052 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_6845
timestamp 1745462530
transform 1 0 1772 0 1 3505
box -2 -2 2 2
use M2_M1  M2_M1_6846
timestamp 1745462530
transform 1 0 1756 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_6847
timestamp 1745462530
transform 1 0 2548 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_6848
timestamp 1745462530
transform 1 0 2356 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_6849
timestamp 1745462530
transform 1 0 2596 0 1 3025
box -2 -2 2 2
use M2_M1  M2_M1_6850
timestamp 1745462530
transform 1 0 2572 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_6851
timestamp 1745462530
transform 1 0 2604 0 1 3105
box -2 -2 2 2
use M2_M1  M2_M1_6852
timestamp 1745462530
transform 1 0 2588 0 1 3035
box -2 -2 2 2
use M2_M1  M2_M1_6853
timestamp 1745462530
transform 1 0 2564 0 1 3035
box -2 -2 2 2
use M2_M1  M2_M1_6854
timestamp 1745462530
transform 1 0 2540 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_6855
timestamp 1745462530
transform 1 0 2164 0 1 3435
box -2 -2 2 2
use M2_M1  M2_M1_6856
timestamp 1745462530
transform 1 0 2164 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_6857
timestamp 1745462530
transform 1 0 2716 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_6858
timestamp 1745462530
transform 1 0 2684 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_6859
timestamp 1745462530
transform 1 0 2676 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_6860
timestamp 1745462530
transform 1 0 2668 0 1 3885
box -2 -2 2 2
use M2_M1  M2_M1_6861
timestamp 1745462530
transform 1 0 2740 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_6862
timestamp 1745462530
transform 1 0 2668 0 1 3345
box -2 -2 2 2
use M2_M1  M2_M1_6863
timestamp 1745462530
transform 1 0 2684 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_6864
timestamp 1745462530
transform 1 0 2668 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_6865
timestamp 1745462530
transform 1 0 3836 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_6866
timestamp 1745462530
transform 1 0 3820 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_6867
timestamp 1745462530
transform 1 0 3780 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_6868
timestamp 1745462530
transform 1 0 3740 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_6869
timestamp 1745462530
transform 1 0 3004 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_6870
timestamp 1745462530
transform 1 0 2620 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_6871
timestamp 1745462530
transform 1 0 1972 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_6872
timestamp 1745462530
transform 1 0 1900 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_6873
timestamp 1745462530
transform 1 0 3644 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_6874
timestamp 1745462530
transform 1 0 3628 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_6875
timestamp 1745462530
transform 1 0 3588 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_6876
timestamp 1745462530
transform 1 0 3564 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_6877
timestamp 1745462530
transform 1 0 3548 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_6878
timestamp 1745462530
transform 1 0 2980 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_6879
timestamp 1745462530
transform 1 0 2700 0 1 3295
box -2 -2 2 2
use M2_M1  M2_M1_6880
timestamp 1745462530
transform 1 0 2452 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_6881
timestamp 1745462530
transform 1 0 2364 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_6882
timestamp 1745462530
transform 1 0 2116 0 1 3315
box -2 -2 2 2
use M2_M1  M2_M1_6883
timestamp 1745462530
transform 1 0 2772 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_6884
timestamp 1745462530
transform 1 0 2748 0 1 3315
box -2 -2 2 2
use M2_M1  M2_M1_6885
timestamp 1745462530
transform 1 0 3524 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_6886
timestamp 1745462530
transform 1 0 3476 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_6887
timestamp 1745462530
transform 1 0 3428 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_6888
timestamp 1745462530
transform 1 0 3380 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_6889
timestamp 1745462530
transform 1 0 2964 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_6890
timestamp 1745462530
transform 1 0 2788 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_6891
timestamp 1745462530
transform 1 0 2660 0 1 3715
box -2 -2 2 2
use M2_M1  M2_M1_6892
timestamp 1745462530
transform 1 0 2596 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_6893
timestamp 1745462530
transform 1 0 2556 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_6894
timestamp 1745462530
transform 1 0 2964 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_6895
timestamp 1745462530
transform 1 0 2892 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_6896
timestamp 1745462530
transform 1 0 2860 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_6897
timestamp 1745462530
transform 1 0 2996 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_6898
timestamp 1745462530
transform 1 0 2964 0 1 3395
box -2 -2 2 2
use M2_M1  M2_M1_6899
timestamp 1745462530
transform 1 0 3020 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_6900
timestamp 1745462530
transform 1 0 2996 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_6901
timestamp 1745462530
transform 1 0 2996 0 1 3315
box -2 -2 2 2
use M2_M1  M2_M1_6902
timestamp 1745462530
transform 1 0 2948 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_6903
timestamp 1745462530
transform 1 0 4076 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_6904
timestamp 1745462530
transform 1 0 3996 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_6905
timestamp 1745462530
transform 1 0 3892 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_6906
timestamp 1745462530
transform 1 0 3868 0 1 3345
box -2 -2 2 2
use M2_M1  M2_M1_6907
timestamp 1745462530
transform 1 0 3644 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_6908
timestamp 1745462530
transform 1 0 3892 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_6909
timestamp 1745462530
transform 1 0 3804 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_6910
timestamp 1745462530
transform 1 0 3644 0 1 3315
box -2 -2 2 2
use M2_M1  M2_M1_6911
timestamp 1745462530
transform 1 0 3460 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_6912
timestamp 1745462530
transform 1 0 4044 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_6913
timestamp 1745462530
transform 1 0 4020 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_6914
timestamp 1745462530
transform 1 0 3924 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_6915
timestamp 1745462530
transform 1 0 3876 0 1 3395
box -2 -2 2 2
use M2_M1  M2_M1_6916
timestamp 1745462530
transform 1 0 3692 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_6917
timestamp 1745462530
transform 1 0 3916 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_6918
timestamp 1745462530
transform 1 0 3836 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_6919
timestamp 1745462530
transform 1 0 3676 0 1 3315
box -2 -2 2 2
use M2_M1  M2_M1_6920
timestamp 1745462530
transform 1 0 3508 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_6921
timestamp 1745462530
transform 1 0 4172 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_6922
timestamp 1745462530
transform 1 0 4140 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_6923
timestamp 1745462530
transform 1 0 3932 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_6924
timestamp 1745462530
transform 1 0 3924 0 1 3395
box -2 -2 2 2
use M2_M1  M2_M1_6925
timestamp 1745462530
transform 1 0 3572 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_6926
timestamp 1745462530
transform 1 0 3940 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_6927
timestamp 1745462530
transform 1 0 3900 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_6928
timestamp 1745462530
transform 1 0 3564 0 1 3315
box -2 -2 2 2
use M2_M1  M2_M1_6929
timestamp 1745462530
transform 1 0 3412 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_6930
timestamp 1745462530
transform 1 0 3964 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_6931
timestamp 1745462530
transform 1 0 3940 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_6932
timestamp 1745462530
transform 1 0 3804 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_6933
timestamp 1745462530
transform 1 0 3772 0 1 3395
box -2 -2 2 2
use M2_M1  M2_M1_6934
timestamp 1745462530
transform 1 0 3612 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_6935
timestamp 1745462530
transform 1 0 3804 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_6936
timestamp 1745462530
transform 1 0 3772 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_6937
timestamp 1745462530
transform 1 0 3604 0 1 3315
box -2 -2 2 2
use M2_M1  M2_M1_6938
timestamp 1745462530
transform 1 0 3364 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_6939
timestamp 1745462530
transform 1 0 2052 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_6940
timestamp 1745462530
transform 1 0 2012 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_6941
timestamp 1745462530
transform 1 0 2004 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_6942
timestamp 1745462530
transform 1 0 2468 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_6943
timestamp 1745462530
transform 1 0 2020 0 1 3395
box -2 -2 2 2
use M2_M1  M2_M1_6944
timestamp 1745462530
transform 1 0 2044 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_6945
timestamp 1745462530
transform 1 0 2020 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_6946
timestamp 1745462530
transform 1 0 2516 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_6947
timestamp 1745462530
transform 1 0 2492 0 1 3315
box -2 -2 2 2
use M2_M1  M2_M1_6948
timestamp 1745462530
transform 1 0 1964 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_6949
timestamp 1745462530
transform 1 0 1964 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_6950
timestamp 1745462530
transform 1 0 1932 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_6951
timestamp 1745462530
transform 1 0 2412 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_6952
timestamp 1745462530
transform 1 0 1932 0 1 3395
box -2 -2 2 2
use M2_M1  M2_M1_6953
timestamp 1745462530
transform 1 0 1948 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_6954
timestamp 1745462530
transform 1 0 1932 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_6955
timestamp 1745462530
transform 1 0 2580 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_6956
timestamp 1745462530
transform 1 0 2428 0 1 3355
box -2 -2 2 2
use M2_M1  M2_M1_6957
timestamp 1745462530
transform 1 0 2428 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_6958
timestamp 1745462530
transform 1 0 2428 0 1 3315
box -2 -2 2 2
use M2_M1  M2_M1_6959
timestamp 1745462530
transform 1 0 2748 0 1 3025
box -2 -2 2 2
use M2_M1  M2_M1_6960
timestamp 1745462530
transform 1 0 2740 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_6961
timestamp 1745462530
transform 1 0 2796 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_6962
timestamp 1745462530
transform 1 0 2740 0 1 3035
box -2 -2 2 2
use M2_M1  M2_M1_6963
timestamp 1745462530
transform 1 0 2044 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_6964
timestamp 1745462530
transform 1 0 1900 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_6965
timestamp 1745462530
transform 1 0 1868 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_6966
timestamp 1745462530
transform 1 0 2684 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_6967
timestamp 1745462530
transform 1 0 2020 0 1 3195
box -2 -2 2 2
use M2_M1  M2_M1_6968
timestamp 1745462530
transform 1 0 2036 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_6969
timestamp 1745462530
transform 1 0 2020 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_6970
timestamp 1745462530
transform 1 0 3812 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_6971
timestamp 1745462530
transform 1 0 3812 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_6972
timestamp 1745462530
transform 1 0 3796 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_6973
timestamp 1745462530
transform 1 0 3708 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_6974
timestamp 1745462530
transform 1 0 1980 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_6975
timestamp 1745462530
transform 1 0 1972 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_6976
timestamp 1745462530
transform 1 0 1948 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_6977
timestamp 1745462530
transform 1 0 1924 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_6978
timestamp 1745462530
transform 1 0 1828 0 1 3425
box -2 -2 2 2
use M2_M1  M2_M1_6979
timestamp 1745462530
transform 1 0 1812 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_6980
timestamp 1745462530
transform 1 0 3564 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_6981
timestamp 1745462530
transform 1 0 3556 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_6982
timestamp 1745462530
transform 1 0 3540 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_6983
timestamp 1745462530
transform 1 0 3532 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_6984
timestamp 1745462530
transform 1 0 2812 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_6985
timestamp 1745462530
transform 1 0 2660 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_6986
timestamp 1745462530
transform 1 0 2476 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_6987
timestamp 1745462530
transform 1 0 2308 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_6988
timestamp 1745462530
transform 1 0 2268 0 1 3315
box -2 -2 2 2
use M2_M1  M2_M1_6989
timestamp 1745462530
transform 1 0 2780 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_6990
timestamp 1745462530
transform 1 0 2700 0 1 3225
box -2 -2 2 2
use M2_M1  M2_M1_6991
timestamp 1745462530
transform 1 0 3516 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_6992
timestamp 1745462530
transform 1 0 3508 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_6993
timestamp 1745462530
transform 1 0 3460 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_6994
timestamp 1745462530
transform 1 0 3404 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_6995
timestamp 1745462530
transform 1 0 2876 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_6996
timestamp 1745462530
transform 1 0 2804 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_6997
timestamp 1745462530
transform 1 0 2572 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_6998
timestamp 1745462530
transform 1 0 2564 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_6999
timestamp 1745462530
transform 1 0 1900 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_7000
timestamp 1745462530
transform 1 0 1916 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_7001
timestamp 1745462530
transform 1 0 1820 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_7002
timestamp 1745462530
transform 1 0 1788 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_7003
timestamp 1745462530
transform 1 0 2852 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_7004
timestamp 1745462530
transform 1 0 1932 0 1 3345
box -2 -2 2 2
use M2_M1  M2_M1_7005
timestamp 1745462530
transform 1 0 2004 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_7006
timestamp 1745462530
transform 1 0 1972 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_7007
timestamp 1745462530
transform 1 0 2860 0 1 3225
box -2 -2 2 2
use M2_M1  M2_M1_7008
timestamp 1745462530
transform 1 0 2860 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_7009
timestamp 1745462530
transform 1 0 4220 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_7010
timestamp 1745462530
transform 1 0 4204 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_7011
timestamp 1745462530
transform 1 0 3900 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_7012
timestamp 1745462530
transform 1 0 3860 0 1 3195
box -2 -2 2 2
use M2_M1  M2_M1_7013
timestamp 1745462530
transform 1 0 3636 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_7014
timestamp 1745462530
transform 1 0 3892 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_7015
timestamp 1745462530
transform 1 0 3820 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_7016
timestamp 1745462530
transform 1 0 3612 0 1 3115
box -2 -2 2 2
use M2_M1  M2_M1_7017
timestamp 1745462530
transform 1 0 3500 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_7018
timestamp 1745462530
transform 1 0 4212 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_7019
timestamp 1745462530
transform 1 0 4188 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_7020
timestamp 1745462530
transform 1 0 3876 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_7021
timestamp 1745462530
transform 1 0 3844 0 1 3345
box -2 -2 2 2
use M2_M1  M2_M1_7022
timestamp 1745462530
transform 1 0 3612 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_7023
timestamp 1745462530
transform 1 0 3868 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_7024
timestamp 1745462530
transform 1 0 3852 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_7025
timestamp 1745462530
transform 1 0 3596 0 1 3225
box -2 -2 2 2
use M2_M1  M2_M1_7026
timestamp 1745462530
transform 1 0 3492 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_7027
timestamp 1745462530
transform 1 0 4036 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_7028
timestamp 1745462530
transform 1 0 3988 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_7029
timestamp 1745462530
transform 1 0 3924 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_7030
timestamp 1745462530
transform 1 0 3892 0 1 3195
box -2 -2 2 2
use M2_M1  M2_M1_7031
timestamp 1745462530
transform 1 0 3580 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_7032
timestamp 1745462530
transform 1 0 3916 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_7033
timestamp 1745462530
transform 1 0 3852 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_7034
timestamp 1745462530
transform 1 0 3564 0 1 3115
box -2 -2 2 2
use M2_M1  M2_M1_7035
timestamp 1745462530
transform 1 0 3444 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_7036
timestamp 1745462530
transform 1 0 3956 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_7037
timestamp 1745462530
transform 1 0 3932 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_7038
timestamp 1745462530
transform 1 0 3708 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_7039
timestamp 1745462530
transform 1 0 3676 0 1 3195
box -2 -2 2 2
use M2_M1  M2_M1_7040
timestamp 1745462530
transform 1 0 3556 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_7041
timestamp 1745462530
transform 1 0 3724 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_7042
timestamp 1745462530
transform 1 0 3716 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_7043
timestamp 1745462530
transform 1 0 3564 0 1 3225
box -2 -2 2 2
use M2_M1  M2_M1_7044
timestamp 1745462530
transform 1 0 3388 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_7045
timestamp 1745462530
transform 1 0 1876 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_7046
timestamp 1745462530
transform 1 0 1700 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_7047
timestamp 1745462530
transform 1 0 1668 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_7048
timestamp 1745462530
transform 1 0 2508 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_7049
timestamp 1745462530
transform 1 0 1868 0 1 3195
box -2 -2 2 2
use M2_M1  M2_M1_7050
timestamp 1745462530
transform 1 0 1940 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_7051
timestamp 1745462530
transform 1 0 1916 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_7052
timestamp 1745462530
transform 1 0 2556 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_7053
timestamp 1745462530
transform 1 0 2532 0 1 3225
box -2 -2 2 2
use M2_M1  M2_M1_7054
timestamp 1745462530
transform 1 0 1828 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_7055
timestamp 1745462530
transform 1 0 1684 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_7056
timestamp 1745462530
transform 1 0 1652 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_7057
timestamp 1745462530
transform 1 0 2364 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_7058
timestamp 1745462530
transform 1 0 1812 0 1 3145
box -2 -2 2 2
use M2_M1  M2_M1_7059
timestamp 1745462530
transform 1 0 1844 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_7060
timestamp 1745462530
transform 1 0 1836 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_7061
timestamp 1745462530
transform 1 0 2524 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_7062
timestamp 1745462530
transform 1 0 2364 0 1 3115
box -2 -2 2 2
use M2_M1  M2_M1_7063
timestamp 1745462530
transform 1 0 2780 0 1 3025
box -2 -2 2 2
use M2_M1  M2_M1_7064
timestamp 1745462530
transform 1 0 2772 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_7065
timestamp 1745462530
transform 1 0 2756 0 1 3035
box -2 -2 2 2
use M2_M1  M2_M1_7066
timestamp 1745462530
transform 1 0 2716 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_7067
timestamp 1745462530
transform 1 0 2308 0 1 3305
box -2 -2 2 2
use M2_M1  M2_M1_7068
timestamp 1745462530
transform 1 0 2212 0 1 3305
box -2 -2 2 2
use M2_M1  M2_M1_7069
timestamp 1745462530
transform 1 0 2156 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_7070
timestamp 1745462530
transform 1 0 1764 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_7071
timestamp 1745462530
transform 1 0 1748 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_7072
timestamp 1745462530
transform 1 0 1716 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_7073
timestamp 1745462530
transform 1 0 2628 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_7074
timestamp 1745462530
transform 1 0 1756 0 1 3345
box -2 -2 2 2
use M2_M1  M2_M1_7075
timestamp 1745462530
transform 1 0 1828 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_7076
timestamp 1745462530
transform 1 0 1780 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_7077
timestamp 1745462530
transform 1 0 3756 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_7078
timestamp 1745462530
transform 1 0 3732 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_7079
timestamp 1745462530
transform 1 0 3652 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_7080
timestamp 1745462530
transform 1 0 3084 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_7081
timestamp 1745462530
transform 1 0 2156 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_7082
timestamp 1745462530
transform 1 0 2140 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_7083
timestamp 1745462530
transform 1 0 1860 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_7084
timestamp 1745462530
transform 1 0 1804 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_7085
timestamp 1745462530
transform 1 0 1756 0 1 3425
box -2 -2 2 2
use M2_M1  M2_M1_7086
timestamp 1745462530
transform 1 0 3420 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_7087
timestamp 1745462530
transform 1 0 3404 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_7088
timestamp 1745462530
transform 1 0 3332 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_7089
timestamp 1745462530
transform 1 0 3228 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_7090
timestamp 1745462530
transform 1 0 2828 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_7091
timestamp 1745462530
transform 1 0 2580 0 1 3225
box -2 -2 2 2
use M2_M1  M2_M1_7092
timestamp 1745462530
transform 1 0 2372 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_7093
timestamp 1745462530
transform 1 0 2300 0 1 3315
box -2 -2 2 2
use M2_M1  M2_M1_7094
timestamp 1745462530
transform 1 0 2284 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_7095
timestamp 1745462530
transform 1 0 2724 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_7096
timestamp 1745462530
transform 1 0 2652 0 1 3225
box -2 -2 2 2
use M2_M1  M2_M1_7097
timestamp 1745462530
transform 1 0 3380 0 1 3235
box -2 -2 2 2
use M2_M1  M2_M1_7098
timestamp 1745462530
transform 1 0 3324 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_7099
timestamp 1745462530
transform 1 0 3300 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_7100
timestamp 1745462530
transform 1 0 3260 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_7101
timestamp 1745462530
transform 1 0 2908 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_7102
timestamp 1745462530
transform 1 0 2740 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_7103
timestamp 1745462530
transform 1 0 2460 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_7104
timestamp 1745462530
transform 1 0 2452 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_7105
timestamp 1745462530
transform 1 0 1804 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_7106
timestamp 1745462530
transform 1 0 1908 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_7107
timestamp 1745462530
transform 1 0 1740 0 1 4005
box -2 -2 2 2
use M2_M1  M2_M1_7108
timestamp 1745462530
transform 1 0 1692 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_7109
timestamp 1745462530
transform 1 0 2844 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_7110
timestamp 1745462530
transform 1 0 1900 0 1 3345
box -2 -2 2 2
use M2_M1  M2_M1_7111
timestamp 1745462530
transform 1 0 1916 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_7112
timestamp 1745462530
transform 1 0 1900 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_7113
timestamp 1745462530
transform 1 0 2892 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_7114
timestamp 1745462530
transform 1 0 2860 0 1 3315
box -2 -2 2 2
use M2_M1  M2_M1_7115
timestamp 1745462530
transform 1 0 3004 0 1 3115
box -2 -2 2 2
use M2_M1  M2_M1_7116
timestamp 1745462530
transform 1 0 2956 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_7117
timestamp 1745462530
transform 1 0 3084 0 1 3105
box -2 -2 2 2
use M2_M1  M2_M1_7118
timestamp 1745462530
transform 1 0 3036 0 1 3025
box -2 -2 2 2
use M2_M1  M2_M1_7119
timestamp 1745462530
transform 1 0 2972 0 1 3115
box -2 -2 2 2
use M2_M1  M2_M1_7120
timestamp 1745462530
transform 1 0 2948 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_7121
timestamp 1745462530
transform 1 0 2948 0 1 2855
box -2 -2 2 2
use M2_M1  M2_M1_7122
timestamp 1745462530
transform 1 0 2932 0 1 2855
box -2 -2 2 2
use M2_M1  M2_M1_7123
timestamp 1745462530
transform 1 0 2924 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_7124
timestamp 1745462530
transform 1 0 2900 0 1 2995
box -2 -2 2 2
use M2_M1  M2_M1_7125
timestamp 1745462530
transform 1 0 2556 0 1 1745
box -2 -2 2 2
use M2_M1  M2_M1_7126
timestamp 1745462530
transform 1 0 3020 0 1 3105
box -2 -2 2 2
use M2_M1  M2_M1_7127
timestamp 1745462530
transform 1 0 3004 0 1 3025
box -2 -2 2 2
use M2_M1  M2_M1_7128
timestamp 1745462530
transform 1 0 2996 0 1 3105
box -2 -2 2 2
use M2_M1  M2_M1_7129
timestamp 1745462530
transform 1 0 2964 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_7130
timestamp 1745462530
transform 1 0 2900 0 1 3025
box -2 -2 2 2
use M2_M1  M2_M1_7131
timestamp 1745462530
transform 1 0 2460 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_7132
timestamp 1745462530
transform 1 0 4204 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_7133
timestamp 1745462530
transform 1 0 4172 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_7134
timestamp 1745462530
transform 1 0 3804 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_7135
timestamp 1745462530
transform 1 0 3740 0 1 3145
box -2 -2 2 2
use M2_M1  M2_M1_7136
timestamp 1745462530
transform 1 0 3372 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_7137
timestamp 1745462530
transform 1 0 3780 0 1 3185
box -2 -2 2 2
use M2_M1  M2_M1_7138
timestamp 1745462530
transform 1 0 3780 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_7139
timestamp 1745462530
transform 1 0 3348 0 1 3115
box -2 -2 2 2
use M2_M1  M2_M1_7140
timestamp 1745462530
transform 1 0 3284 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_7141
timestamp 1745462530
transform 1 0 3156 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_7142
timestamp 1745462530
transform 1 0 3068 0 1 3025
box -2 -2 2 2
use M2_M1  M2_M1_7143
timestamp 1745462530
transform 1 0 3052 0 1 3035
box -2 -2 2 2
use M2_M1  M2_M1_7144
timestamp 1745462530
transform 1 0 2996 0 1 3035
box -2 -2 2 2
use M2_M1  M2_M1_7145
timestamp 1745462530
transform 1 0 2980 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_7146
timestamp 1745462530
transform 1 0 2892 0 1 3035
box -2 -2 2 2
use M2_M1  M2_M1_7147
timestamp 1745462530
transform 1 0 2852 0 1 3035
box -2 -2 2 2
use M2_M1  M2_M1_7148
timestamp 1745462530
transform 1 0 2596 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_7149
timestamp 1745462530
transform 1 0 4212 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_7150
timestamp 1745462530
transform 1 0 4188 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_7151
timestamp 1745462530
transform 1 0 3740 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_7152
timestamp 1745462530
transform 1 0 3716 0 1 3195
box -2 -2 2 2
use M2_M1  M2_M1_7153
timestamp 1745462530
transform 1 0 3460 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_7154
timestamp 1745462530
transform 1 0 3756 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_7155
timestamp 1745462530
transform 1 0 3748 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_7156
timestamp 1745462530
transform 1 0 3460 0 1 3225
box -2 -2 2 2
use M2_M1  M2_M1_7157
timestamp 1745462530
transform 1 0 3356 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_7158
timestamp 1745462530
transform 1 0 3188 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_7159
timestamp 1745462530
transform 1 0 3108 0 1 3115
box -2 -2 2 2
use M2_M1  M2_M1_7160
timestamp 1745462530
transform 1 0 4068 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_7161
timestamp 1745462530
transform 1 0 4028 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_7162
timestamp 1745462530
transform 1 0 3636 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_7163
timestamp 1745462530
transform 1 0 3604 0 1 3195
box -2 -2 2 2
use M2_M1  M2_M1_7164
timestamp 1745462530
transform 1 0 3428 0 1 3195
box -2 -2 2 2
use M2_M1  M2_M1_7165
timestamp 1745462530
transform 1 0 3668 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_7166
timestamp 1745462530
transform 1 0 3644 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_7167
timestamp 1745462530
transform 1 0 3428 0 1 3225
box -2 -2 2 2
use M2_M1  M2_M1_7168
timestamp 1745462530
transform 1 0 3308 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_7169
timestamp 1745462530
transform 1 0 3172 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_7170
timestamp 1745462530
transform 1 0 3028 0 1 3025
box -2 -2 2 2
use M2_M1  M2_M1_7171
timestamp 1745462530
transform 1 0 3820 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_7172
timestamp 1745462530
transform 1 0 3804 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_7173
timestamp 1745462530
transform 1 0 3260 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_7174
timestamp 1745462530
transform 1 0 3268 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_7175
timestamp 1745462530
transform 1 0 3116 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_7176
timestamp 1745462530
transform 1 0 3244 0 1 3225
box -2 -2 2 2
use M2_M1  M2_M1_7177
timestamp 1745462530
transform 1 0 3228 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_7178
timestamp 1745462530
transform 1 0 3100 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_7179
timestamp 1745462530
transform 1 0 3060 0 1 3115
box -2 -2 2 2
use M2_M1  M2_M1_7180
timestamp 1745462530
transform 1 0 2100 0 1 3345
box -2 -2 2 2
use M2_M1  M2_M1_7181
timestamp 1745462530
transform 1 0 2100 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_7182
timestamp 1745462530
transform 1 0 2100 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_7183
timestamp 1745462530
transform 1 0 1596 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_7184
timestamp 1745462530
transform 1 0 1564 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_7185
timestamp 1745462530
transform 1 0 2388 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_7186
timestamp 1745462530
transform 1 0 2092 0 1 3195
box -2 -2 2 2
use M2_M1  M2_M1_7187
timestamp 1745462530
transform 1 0 2156 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_7188
timestamp 1745462530
transform 1 0 2124 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_7189
timestamp 1745462530
transform 1 0 2436 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_7190
timestamp 1745462530
transform 1 0 2412 0 1 3225
box -2 -2 2 2
use M2_M1  M2_M1_7191
timestamp 1745462530
transform 1 0 2860 0 1 3025
box -2 -2 2 2
use M2_M1  M2_M1_7192
timestamp 1745462530
transform 1 0 2788 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_7193
timestamp 1745462530
transform 1 0 2828 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_7194
timestamp 1745462530
transform 1 0 2820 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_7195
timestamp 1745462530
transform 1 0 2788 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_7196
timestamp 1745462530
transform 1 0 2876 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_7197
timestamp 1745462530
transform 1 0 2820 0 1 3395
box -2 -2 2 2
use M2_M1  M2_M1_7198
timestamp 1745462530
transform 1 0 2836 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_7199
timestamp 1745462530
transform 1 0 2820 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_7200
timestamp 1745462530
transform 1 0 1700 0 1 3505
box -2 -2 2 2
use M2_M1  M2_M1_7201
timestamp 1745462530
transform 1 0 1684 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_7202
timestamp 1745462530
transform 1 0 2884 0 1 3425
box -2 -2 2 2
use M2_M1  M2_M1_7203
timestamp 1745462530
transform 1 0 2884 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_7204
timestamp 1745462530
transform 1 0 2652 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_7205
timestamp 1745462530
transform 1 0 2652 0 1 3025
box -2 -2 2 2
use M2_M1  M2_M1_7206
timestamp 1745462530
transform 1 0 2916 0 1 3025
box -2 -2 2 2
use M2_M1  M2_M1_7207
timestamp 1745462530
transform 1 0 2876 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_7208
timestamp 1745462530
transform 1 0 2260 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_7209
timestamp 1745462530
transform 1 0 1628 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_7210
timestamp 1745462530
transform 1 0 1596 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_7211
timestamp 1745462530
transform 1 0 2300 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_7212
timestamp 1745462530
transform 1 0 2236 0 1 3195
box -2 -2 2 2
use M2_M1  M2_M1_7213
timestamp 1745462530
transform 1 0 2252 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_7214
timestamp 1745462530
transform 1 0 2236 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_7215
timestamp 1745462530
transform 1 0 2444 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_7216
timestamp 1745462530
transform 1 0 2332 0 1 3115
box -2 -2 2 2
use M2_M1  M2_M1_7217
timestamp 1745462530
transform 1 0 2932 0 1 3115
box -2 -2 2 2
use M2_M1  M2_M1_7218
timestamp 1745462530
transform 1 0 2804 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_7219
timestamp 1745462530
transform 1 0 2556 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_7220
timestamp 1745462530
transform 1 0 2532 0 1 1745
box -2 -2 2 2
use M2_M1  M2_M1_7221
timestamp 1745462530
transform 1 0 2548 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_7222
timestamp 1745462530
transform 1 0 2532 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_7223
timestamp 1745462530
transform 1 0 3724 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_7224
timestamp 1745462530
transform 1 0 2484 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_7225
timestamp 1745462530
transform 1 0 2492 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_7226
timestamp 1745462530
transform 1 0 2068 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_7227
timestamp 1745462530
transform 1 0 2036 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_7228
timestamp 1745462530
transform 1 0 1012 0 1 1795
box -2 -2 2 2
use M2_M1  M2_M1_7229
timestamp 1745462530
transform 1 0 2060 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_7230
timestamp 1745462530
transform 1 0 828 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_7231
timestamp 1745462530
transform 1 0 2092 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_7232
timestamp 1745462530
transform 1 0 2092 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_7233
timestamp 1745462530
transform 1 0 2084 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_7234
timestamp 1745462530
transform 1 0 2060 0 1 1035
box -2 -2 2 2
use M2_M1  M2_M1_7235
timestamp 1745462530
transform 1 0 2084 0 1 995
box -2 -2 2 2
use M2_M1  M2_M1_7236
timestamp 1745462530
transform 1 0 2084 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_7237
timestamp 1745462530
transform 1 0 2140 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_7238
timestamp 1745462530
transform 1 0 2124 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7239
timestamp 1745462530
transform 1 0 2596 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_7240
timestamp 1745462530
transform 1 0 2596 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_7241
timestamp 1745462530
transform 1 0 2564 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_7242
timestamp 1745462530
transform 1 0 2540 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_7243
timestamp 1745462530
transform 1 0 2452 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_7244
timestamp 1745462530
transform 1 0 2548 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_7245
timestamp 1745462530
transform 1 0 2516 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_7246
timestamp 1745462530
transform 1 0 2492 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_7247
timestamp 1745462530
transform 1 0 2460 0 1 2295
box -2 -2 2 2
use M2_M1  M2_M1_7248
timestamp 1745462530
transform 1 0 2500 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_7249
timestamp 1745462530
transform 1 0 2468 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_7250
timestamp 1745462530
transform 1 0 2436 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_7251
timestamp 1745462530
transform 1 0 2412 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_7252
timestamp 1745462530
transform 1 0 2412 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_7253
timestamp 1745462530
transform 1 0 2068 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_7254
timestamp 1745462530
transform 1 0 2020 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_7255
timestamp 1745462530
transform 1 0 2492 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_7256
timestamp 1745462530
transform 1 0 2484 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_7257
timestamp 1745462530
transform 1 0 2460 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_7258
timestamp 1745462530
transform 1 0 2436 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_7259
timestamp 1745462530
transform 1 0 2636 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_7260
timestamp 1745462530
transform 1 0 2596 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_7261
timestamp 1745462530
transform 1 0 2572 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_7262
timestamp 1745462530
transform 1 0 2548 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_7263
timestamp 1745462530
transform 1 0 2532 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_7264
timestamp 1745462530
transform 1 0 2108 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_7265
timestamp 1745462530
transform 1 0 2100 0 1 1395
box -2 -2 2 2
use M2_M1  M2_M1_7266
timestamp 1745462530
transform 1 0 2116 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_7267
timestamp 1745462530
transform 1 0 2116 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_7268
timestamp 1745462530
transform 1 0 2492 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_7269
timestamp 1745462530
transform 1 0 2484 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_7270
timestamp 1745462530
transform 1 0 2452 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_7271
timestamp 1745462530
transform 1 0 2452 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_7272
timestamp 1745462530
transform 1 0 2444 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_7273
timestamp 1745462530
transform 1 0 2164 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_7274
timestamp 1745462530
transform 1 0 2092 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_7275
timestamp 1745462530
transform 1 0 2356 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_7276
timestamp 1745462530
transform 1 0 2348 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_7277
timestamp 1745462530
transform 1 0 2348 0 1 2105
box -2 -2 2 2
use M2_M1  M2_M1_7278
timestamp 1745462530
transform 1 0 2332 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_7279
timestamp 1745462530
transform 1 0 2324 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_7280
timestamp 1745462530
transform 1 0 2300 0 1 2035
box -2 -2 2 2
use M2_M1  M2_M1_7281
timestamp 1745462530
transform 1 0 2420 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_7282
timestamp 1745462530
transform 1 0 2404 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_7283
timestamp 1745462530
transform 1 0 2388 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_7284
timestamp 1745462530
transform 1 0 2380 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_7285
timestamp 1745462530
transform 1 0 2380 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_7286
timestamp 1745462530
transform 1 0 836 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_7287
timestamp 1745462530
transform 1 0 732 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_7288
timestamp 1745462530
transform 1 0 812 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_7289
timestamp 1745462530
transform 1 0 804 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_7290
timestamp 1745462530
transform 1 0 956 0 1 1795
box -2 -2 2 2
use M2_M1  M2_M1_7291
timestamp 1745462530
transform 1 0 948 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_7292
timestamp 1745462530
transform 1 0 980 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_7293
timestamp 1745462530
transform 1 0 964 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_7294
timestamp 1745462530
transform 1 0 2116 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_7295
timestamp 1745462530
transform 1 0 2068 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_7296
timestamp 1745462530
transform 1 0 3724 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_7297
timestamp 1745462530
transform 1 0 3700 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_7298
timestamp 1745462530
transform 1 0 3732 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_7299
timestamp 1745462530
transform 1 0 3692 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_7300
timestamp 1745462530
transform 1 0 3780 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_7301
timestamp 1745462530
transform 1 0 3764 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_7302
timestamp 1745462530
transform 1 0 3732 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_7303
timestamp 1745462530
transform 1 0 3708 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_7304
timestamp 1745462530
transform 1 0 3788 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_7305
timestamp 1745462530
transform 1 0 3708 0 1 2545
box -2 -2 2 2
use M2_M1  M2_M1_7306
timestamp 1745462530
transform 1 0 3740 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_7307
timestamp 1745462530
transform 1 0 3684 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_7308
timestamp 1745462530
transform 1 0 3804 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_7309
timestamp 1745462530
transform 1 0 3780 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_7310
timestamp 1745462530
transform 1 0 3820 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_7311
timestamp 1745462530
transform 1 0 3772 0 1 2345
box -2 -2 2 2
use M2_M1  M2_M1_7312
timestamp 1745462530
transform 1 0 3788 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_7313
timestamp 1745462530
transform 1 0 3116 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_7314
timestamp 1745462530
transform 1 0 3780 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_7315
timestamp 1745462530
transform 1 0 3700 0 1 945
box -2 -2 2 2
use M2_M1  M2_M1_7316
timestamp 1745462530
transform 1 0 3724 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_7317
timestamp 1745462530
transform 1 0 3660 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_7318
timestamp 1745462530
transform 1 0 3772 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_7319
timestamp 1745462530
transform 1 0 3692 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_7320
timestamp 1745462530
transform 1 0 3820 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_7321
timestamp 1745462530
transform 1 0 3716 0 1 1195
box -2 -2 2 2
use M2_M1  M2_M1_7322
timestamp 1745462530
transform 1 0 3740 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7323
timestamp 1745462530
transform 1 0 3716 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_7324
timestamp 1745462530
transform 1 0 2220 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_7325
timestamp 1745462530
transform 1 0 2212 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_7326
timestamp 1745462530
transform 1 0 2508 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_7327
timestamp 1745462530
transform 1 0 2508 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_7328
timestamp 1745462530
transform 1 0 2492 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_7329
timestamp 1745462530
transform 1 0 2492 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_7330
timestamp 1745462530
transform 1 0 2508 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_7331
timestamp 1745462530
transform 1 0 1908 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_7332
timestamp 1745462530
transform 1 0 1892 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_7333
timestamp 1745462530
transform 1 0 1892 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_7334
timestamp 1745462530
transform 1 0 1916 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_7335
timestamp 1745462530
transform 1 0 1900 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_7336
timestamp 1745462530
transform 1 0 1924 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_7337
timestamp 1745462530
transform 1 0 1148 0 1 1555
box -2 -2 2 2
use M2_M1  M2_M1_7338
timestamp 1745462530
transform 1 0 1916 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_7339
timestamp 1745462530
transform 1 0 796 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_7340
timestamp 1745462530
transform 1 0 828 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_7341
timestamp 1745462530
transform 1 0 780 0 1 995
box -2 -2 2 2
use M2_M1  M2_M1_7342
timestamp 1745462530
transform 1 0 804 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7343
timestamp 1745462530
transform 1 0 732 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_7344
timestamp 1745462530
transform 1 0 828 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_7345
timestamp 1745462530
transform 1 0 788 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_7346
timestamp 1745462530
transform 1 0 1108 0 1 1545
box -2 -2 2 2
use M2_M1  M2_M1_7347
timestamp 1745462530
transform 1 0 1020 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_7348
timestamp 1745462530
transform 1 0 1124 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_7349
timestamp 1745462530
transform 1 0 1100 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_7350
timestamp 1745462530
transform 1 0 1964 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_7351
timestamp 1745462530
transform 1 0 1924 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_7352
timestamp 1745462530
transform 1 0 1884 0 1 2515
box -2 -2 2 2
use M2_M1  M2_M1_7353
timestamp 1745462530
transform 1 0 1836 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_7354
timestamp 1745462530
transform 1 0 1932 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_7355
timestamp 1745462530
transform 1 0 1868 0 1 1795
box -2 -2 2 2
use M2_M1  M2_M1_7356
timestamp 1745462530
transform 1 0 1956 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_7357
timestamp 1745462530
transform 1 0 1924 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_7358
timestamp 1745462530
transform 1 0 2492 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_7359
timestamp 1745462530
transform 1 0 2492 0 1 1355
box -2 -2 2 2
use M2_M1  M2_M1_7360
timestamp 1745462530
transform 1 0 2468 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_7361
timestamp 1745462530
transform 1 0 2460 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7362
timestamp 1745462530
transform 1 0 2628 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_7363
timestamp 1745462530
transform 1 0 2548 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_7364
timestamp 1745462530
transform 1 0 3148 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_7365
timestamp 1745462530
transform 1 0 2540 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_7366
timestamp 1745462530
transform 1 0 3740 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_7367
timestamp 1745462530
transform 1 0 3132 0 1 1395
box -2 -2 2 2
use M2_M1  M2_M1_7368
timestamp 1745462530
transform 1 0 3212 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_7369
timestamp 1745462530
transform 1 0 3172 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_7370
timestamp 1745462530
transform 1 0 3756 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_7371
timestamp 1745462530
transform 1 0 3748 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_7372
timestamp 1745462530
transform 1 0 3724 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_7373
timestamp 1745462530
transform 1 0 2620 0 1 1595
box -2 -2 2 2
use M2_M1  M2_M1_7374
timestamp 1745462530
transform 1 0 2692 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_7375
timestamp 1745462530
transform 1 0 2684 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_7376
timestamp 1745462530
transform 1 0 2548 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_7377
timestamp 1745462530
transform 1 0 2484 0 1 1145
box -2 -2 2 2
use M2_M1  M2_M1_7378
timestamp 1745462530
transform 1 0 2516 0 1 1105
box -2 -2 2 2
use M2_M1  M2_M1_7379
timestamp 1745462530
transform 1 0 2516 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_7380
timestamp 1745462530
transform 1 0 2548 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_7381
timestamp 1745462530
transform 1 0 2532 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_7382
timestamp 1745462530
transform 1 0 2444 0 1 1345
box -2 -2 2 2
use M2_M1  M2_M1_7383
timestamp 1745462530
transform 1 0 2420 0 1 985
box -2 -2 2 2
use M2_M1  M2_M1_7384
timestamp 1745462530
transform 1 0 2404 0 1 985
box -2 -2 2 2
use M2_M1  M2_M1_7385
timestamp 1745462530
transform 1 0 2404 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_7386
timestamp 1745462530
transform 1 0 2540 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_7387
timestamp 1745462530
transform 1 0 2508 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_7388
timestamp 1745462530
transform 1 0 2564 0 1 1745
box -2 -2 2 2
use M2_M1  M2_M1_7389
timestamp 1745462530
transform 1 0 2492 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_7390
timestamp 1745462530
transform 1 0 2588 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_7391
timestamp 1745462530
transform 1 0 2468 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_7392
timestamp 1745462530
transform 1 0 3516 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_7393
timestamp 1745462530
transform 1 0 2428 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_7394
timestamp 1745462530
transform 1 0 2420 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_7395
timestamp 1745462530
transform 1 0 1060 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_7396
timestamp 1745462530
transform 1 0 996 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_7397
timestamp 1745462530
transform 1 0 972 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_7398
timestamp 1745462530
transform 1 0 1052 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_7399
timestamp 1745462530
transform 1 0 828 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_7400
timestamp 1745462530
transform 1 0 1140 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_7401
timestamp 1745462530
transform 1 0 1100 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_7402
timestamp 1745462530
transform 1 0 1068 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_7403
timestamp 1745462530
transform 1 0 1068 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_7404
timestamp 1745462530
transform 1 0 1084 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_7405
timestamp 1745462530
transform 1 0 1068 0 1 995
box -2 -2 2 2
use M2_M1  M2_M1_7406
timestamp 1745462530
transform 1 0 1084 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7407
timestamp 1745462530
transform 1 0 1028 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_7408
timestamp 1745462530
transform 1 0 1100 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_7409
timestamp 1745462530
transform 1 0 1100 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_7410
timestamp 1745462530
transform 1 0 1084 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_7411
timestamp 1745462530
transform 1 0 1076 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_7412
timestamp 1745462530
transform 1 0 1148 0 1 1545
box -2 -2 2 2
use M2_M1  M2_M1_7413
timestamp 1745462530
transform 1 0 1132 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_7414
timestamp 1745462530
transform 1 0 1244 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_7415
timestamp 1745462530
transform 1 0 1212 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_7416
timestamp 1745462530
transform 1 0 796 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_7417
timestamp 1745462530
transform 1 0 796 0 1 2395
box -2 -2 2 2
use M2_M1  M2_M1_7418
timestamp 1745462530
transform 1 0 820 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_7419
timestamp 1745462530
transform 1 0 764 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_7420
timestamp 1745462530
transform 1 0 788 0 1 2515
box -2 -2 2 2
use M2_M1  M2_M1_7421
timestamp 1745462530
transform 1 0 764 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_7422
timestamp 1745462530
transform 1 0 996 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_7423
timestamp 1745462530
transform 1 0 940 0 1 1745
box -2 -2 2 2
use M2_M1  M2_M1_7424
timestamp 1745462530
transform 1 0 956 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_7425
timestamp 1745462530
transform 1 0 916 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_7426
timestamp 1745462530
transform 1 0 3484 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_7427
timestamp 1745462530
transform 1 0 3476 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_7428
timestamp 1745462530
transform 1 0 3532 0 1 1555
box -2 -2 2 2
use M2_M1  M2_M1_7429
timestamp 1745462530
transform 1 0 3532 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_7430
timestamp 1745462530
transform 1 0 3508 0 1 1555
box -2 -2 2 2
use M2_M1  M2_M1_7431
timestamp 1745462530
transform 1 0 3492 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_7432
timestamp 1745462530
transform 1 0 3540 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_7433
timestamp 1745462530
transform 1 0 3516 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_7434
timestamp 1745462530
transform 1 0 3556 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_7435
timestamp 1745462530
transform 1 0 3524 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_7436
timestamp 1745462530
transform 1 0 3492 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_7437
timestamp 1745462530
transform 1 0 3492 0 1 2385
box -2 -2 2 2
use M2_M1  M2_M1_7438
timestamp 1745462530
transform 1 0 3644 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_7439
timestamp 1745462530
transform 1 0 3556 0 1 2545
box -2 -2 2 2
use M2_M1  M2_M1_7440
timestamp 1745462530
transform 1 0 3588 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_7441
timestamp 1745462530
transform 1 0 3516 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_7442
timestamp 1745462530
transform 1 0 3660 0 1 2515
box -2 -2 2 2
use M2_M1  M2_M1_7443
timestamp 1745462530
transform 1 0 3596 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_7444
timestamp 1745462530
transform 1 0 3564 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_7445
timestamp 1745462530
transform 1 0 3508 0 1 2345
box -2 -2 2 2
use M2_M1  M2_M1_7446
timestamp 1745462530
transform 1 0 3532 0 1 2305
box -2 -2 2 2
use M2_M1  M2_M1_7447
timestamp 1745462530
transform 1 0 3068 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_7448
timestamp 1745462530
transform 1 0 3636 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_7449
timestamp 1745462530
transform 1 0 3540 0 1 945
box -2 -2 2 2
use M2_M1  M2_M1_7450
timestamp 1745462530
transform 1 0 3596 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_7451
timestamp 1745462530
transform 1 0 3572 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_7452
timestamp 1745462530
transform 1 0 3636 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_7453
timestamp 1745462530
transform 1 0 3636 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_7454
timestamp 1745462530
transform 1 0 3708 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_7455
timestamp 1745462530
transform 1 0 3508 0 1 1195
box -2 -2 2 2
use M2_M1  M2_M1_7456
timestamp 1745462530
transform 1 0 3564 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_7457
timestamp 1745462530
transform 1 0 3524 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7458
timestamp 1745462530
transform 1 0 2812 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_7459
timestamp 1745462530
transform 1 0 2428 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_7460
timestamp 1745462530
transform 1 0 2404 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_7461
timestamp 1745462530
transform 1 0 1396 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_7462
timestamp 1745462530
transform 1 0 1412 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_7463
timestamp 1745462530
transform 1 0 1380 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_7464
timestamp 1745462530
transform 1 0 1428 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_7465
timestamp 1745462530
transform 1 0 1388 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_7466
timestamp 1745462530
transform 1 0 1420 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_7467
timestamp 1745462530
transform 1 0 1188 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_7468
timestamp 1745462530
transform 1 0 1404 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_7469
timestamp 1745462530
transform 1 0 932 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_7470
timestamp 1745462530
transform 1 0 924 0 1 1195
box -2 -2 2 2
use M2_M1  M2_M1_7471
timestamp 1745462530
transform 1 0 812 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_7472
timestamp 1745462530
transform 1 0 956 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7473
timestamp 1745462530
transform 1 0 892 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_7474
timestamp 1745462530
transform 1 0 812 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_7475
timestamp 1745462530
transform 1 0 564 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_7476
timestamp 1745462530
transform 1 0 1156 0 1 1395
box -2 -2 2 2
use M2_M1  M2_M1_7477
timestamp 1745462530
transform 1 0 1028 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_7478
timestamp 1745462530
transform 1 0 1172 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_7479
timestamp 1745462530
transform 1 0 1156 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_7480
timestamp 1745462530
transform 1 0 1500 0 1 2732
box -2 -2 2 2
use M2_M1  M2_M1_7481
timestamp 1745462530
transform 1 0 1412 0 1 2595
box -2 -2 2 2
use M2_M1  M2_M1_7482
timestamp 1745462530
transform 1 0 1484 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_7483
timestamp 1745462530
transform 1 0 1444 0 1 2595
box -2 -2 2 2
use M2_M1  M2_M1_7484
timestamp 1745462530
transform 1 0 1532 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_7485
timestamp 1745462530
transform 1 0 1508 0 1 2755
box -2 -2 2 2
use M2_M1  M2_M1_7486
timestamp 1745462530
transform 1 0 1467 0 1 1804
box -2 -2 2 2
use M2_M1  M2_M1_7487
timestamp 1745462530
transform 1 0 1388 0 1 1595
box -2 -2 2 2
use M2_M1  M2_M1_7488
timestamp 1745462530
transform 1 0 1420 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_7489
timestamp 1745462530
transform 1 0 1404 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_7490
timestamp 1745462530
transform 1 0 2788 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_7491
timestamp 1745462530
transform 1 0 2772 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_7492
timestamp 1745462530
transform 1 0 2820 0 1 1145
box -2 -2 2 2
use M2_M1  M2_M1_7493
timestamp 1745462530
transform 1 0 2804 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_7494
timestamp 1745462530
transform 1 0 2828 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_7495
timestamp 1745462530
transform 1 0 2796 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_7496
timestamp 1745462530
transform 1 0 3244 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_7497
timestamp 1745462530
transform 1 0 2820 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_7498
timestamp 1745462530
transform 1 0 3420 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_7499
timestamp 1745462530
transform 1 0 3252 0 1 1945
box -2 -2 2 2
use M2_M1  M2_M1_7500
timestamp 1745462530
transform 1 0 3268 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_7501
timestamp 1745462530
transform 1 0 3212 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_7502
timestamp 1745462530
transform 1 0 3596 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_7503
timestamp 1745462530
transform 1 0 3444 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_7504
timestamp 1745462530
transform 1 0 3380 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_7505
timestamp 1745462530
transform 1 0 2780 0 1 1995
box -2 -2 2 2
use M2_M1  M2_M1_7506
timestamp 1745462530
transform 1 0 2796 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_7507
timestamp 1745462530
transform 1 0 2788 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_7508
timestamp 1745462530
transform 1 0 2812 0 1 835
box -2 -2 2 2
use M2_M1  M2_M1_7509
timestamp 1745462530
transform 1 0 2780 0 1 1145
box -2 -2 2 2
use M2_M1  M2_M1_7510
timestamp 1745462530
transform 1 0 2804 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_7511
timestamp 1745462530
transform 1 0 2756 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7512
timestamp 1745462530
transform 1 0 2812 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_7513
timestamp 1745462530
transform 1 0 2716 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_7514
timestamp 1745462530
transform 1 0 2804 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_7515
timestamp 1745462530
transform 1 0 2764 0 1 1395
box -2 -2 2 2
use M2_M1  M2_M1_7516
timestamp 1745462530
transform 1 0 2796 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_7517
timestamp 1745462530
transform 1 0 2780 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_7518
timestamp 1745462530
transform 1 0 2492 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_7519
timestamp 1745462530
transform 1 0 2484 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_7520
timestamp 1745462530
transform 1 0 3380 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_7521
timestamp 1745462530
transform 1 0 2468 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_7522
timestamp 1745462530
transform 1 0 2444 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_7523
timestamp 1745462530
transform 1 0 1108 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_7524
timestamp 1745462530
transform 1 0 1100 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_7525
timestamp 1745462530
transform 1 0 900 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_7526
timestamp 1745462530
transform 1 0 1196 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_7527
timestamp 1745462530
transform 1 0 1140 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_7528
timestamp 1745462530
transform 1 0 1180 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7529
timestamp 1745462530
transform 1 0 1156 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_7530
timestamp 1745462530
transform 1 0 1124 0 1 1145
box -2 -2 2 2
use M2_M1  M2_M1_7531
timestamp 1745462530
transform 1 0 1100 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_7532
timestamp 1745462530
transform 1 0 1164 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_7533
timestamp 1745462530
transform 1 0 1100 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7534
timestamp 1745462530
transform 1 0 1132 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_7535
timestamp 1745462530
transform 1 0 1100 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_7536
timestamp 1745462530
transform 1 0 1196 0 1 1395
box -2 -2 2 2
use M2_M1  M2_M1_7537
timestamp 1745462530
transform 1 0 1172 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_7538
timestamp 1745462530
transform 1 0 1284 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_7539
timestamp 1745462530
transform 1 0 1252 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_7540
timestamp 1745462530
transform 1 0 892 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_7541
timestamp 1745462530
transform 1 0 892 0 1 1995
box -2 -2 2 2
use M2_M1  M2_M1_7542
timestamp 1745462530
transform 1 0 916 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_7543
timestamp 1745462530
transform 1 0 868 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_7544
timestamp 1745462530
transform 1 0 876 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_7545
timestamp 1745462530
transform 1 0 852 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_7546
timestamp 1745462530
transform 1 0 1036 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_7547
timestamp 1745462530
transform 1 0 1036 0 1 1745
box -2 -2 2 2
use M2_M1  M2_M1_7548
timestamp 1745462530
transform 1 0 1060 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_7549
timestamp 1745462530
transform 1 0 1044 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_7550
timestamp 1745462530
transform 1 0 3452 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_7551
timestamp 1745462530
transform 1 0 3444 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_7552
timestamp 1745462530
transform 1 0 3420 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_7553
timestamp 1745462530
transform 1 0 3356 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_7554
timestamp 1745462530
transform 1 0 3356 0 1 1255
box -2 -2 2 2
use M2_M1  M2_M1_7555
timestamp 1745462530
transform 1 0 3356 0 1 1235
box -2 -2 2 2
use M2_M1  M2_M1_7556
timestamp 1745462530
transform 1 0 3356 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7557
timestamp 1745462530
transform 1 0 3340 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_7558
timestamp 1745462530
transform 1 0 3404 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_7559
timestamp 1745462530
transform 1 0 3316 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_7560
timestamp 1745462530
transform 1 0 3412 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_7561
timestamp 1745462530
transform 1 0 3356 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_7562
timestamp 1745462530
transform 1 0 3452 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_7563
timestamp 1745462530
transform 1 0 3380 0 1 2595
box -2 -2 2 2
use M2_M1  M2_M1_7564
timestamp 1745462530
transform 1 0 3396 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_7565
timestamp 1745462530
transform 1 0 3284 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_7566
timestamp 1745462530
transform 1 0 3532 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_7567
timestamp 1745462530
transform 1 0 3468 0 1 2625
box -2 -2 2 2
use M2_M1  M2_M1_7568
timestamp 1745462530
transform 1 0 3316 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_7569
timestamp 1745462530
transform 1 0 3292 0 1 2195
box -2 -2 2 2
use M2_M1  M2_M1_7570
timestamp 1745462530
transform 1 0 3316 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_7571
timestamp 1745462530
transform 1 0 2892 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_7572
timestamp 1745462530
transform 1 0 3404 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_7573
timestamp 1745462530
transform 1 0 3348 0 1 1145
box -2 -2 2 2
use M2_M1  M2_M1_7574
timestamp 1745462530
transform 1 0 3364 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_7575
timestamp 1745462530
transform 1 0 3300 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7576
timestamp 1745462530
transform 1 0 3436 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_7577
timestamp 1745462530
transform 1 0 3428 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_7578
timestamp 1745462530
transform 1 0 3380 0 1 1355
box -2 -2 2 2
use M2_M1  M2_M1_7579
timestamp 1745462530
transform 1 0 3380 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_7580
timestamp 1745462530
transform 1 0 3404 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_7581
timestamp 1745462530
transform 1 0 3380 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_7582
timestamp 1745462530
transform 1 0 2508 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_7583
timestamp 1745462530
transform 1 0 2396 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_7584
timestamp 1745462530
transform 1 0 2404 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_7585
timestamp 1745462530
transform 1 0 1188 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_7586
timestamp 1745462530
transform 1 0 1148 0 1 1795
box -2 -2 2 2
use M2_M1  M2_M1_7587
timestamp 1745462530
transform 1 0 1148 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_7588
timestamp 1745462530
transform 1 0 1180 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_7589
timestamp 1745462530
transform 1 0 1124 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_7590
timestamp 1745462530
transform 1 0 1236 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_7591
timestamp 1745462530
transform 1 0 1228 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_7592
timestamp 1745462530
transform 1 0 1196 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_7593
timestamp 1745462530
transform 1 0 940 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7594
timestamp 1745462530
transform 1 0 932 0 1 1155
box -2 -2 2 2
use M2_M1  M2_M1_7595
timestamp 1745462530
transform 1 0 916 0 1 1155
box -2 -2 2 2
use M2_M1  M2_M1_7596
timestamp 1745462530
transform 1 0 916 0 1 1145
box -2 -2 2 2
use M2_M1  M2_M1_7597
timestamp 1745462530
transform 1 0 860 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_7598
timestamp 1745462530
transform 1 0 956 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_7599
timestamp 1745462530
transform 1 0 892 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7600
timestamp 1745462530
transform 1 0 860 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_7601
timestamp 1745462530
transform 1 0 628 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_7602
timestamp 1745462530
transform 1 0 1188 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_7603
timestamp 1745462530
transform 1 0 964 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_7604
timestamp 1745462530
transform 1 0 1220 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_7605
timestamp 1745462530
transform 1 0 1188 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_7606
timestamp 1745462530
transform 1 0 1196 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_7607
timestamp 1745462530
transform 1 0 1108 0 1 2595
box -2 -2 2 2
use M2_M1  M2_M1_7608
timestamp 1745462530
transform 1 0 1164 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_7609
timestamp 1745462530
transform 1 0 1140 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_7610
timestamp 1745462530
transform 1 0 1196 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_7611
timestamp 1745462530
transform 1 0 1196 0 1 2715
box -2 -2 2 2
use M2_M1  M2_M1_7612
timestamp 1745462530
transform 1 0 1108 0 1 1795
box -2 -2 2 2
use M2_M1  M2_M1_7613
timestamp 1745462530
transform 1 0 1100 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_7614
timestamp 1745462530
transform 1 0 1188 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_7615
timestamp 1745462530
transform 1 0 1156 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_7616
timestamp 1745462530
transform 1 0 2508 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_7617
timestamp 1745462530
transform 1 0 2468 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_7618
timestamp 1745462530
transform 1 0 2500 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_7619
timestamp 1745462530
transform 1 0 2452 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7620
timestamp 1745462530
transform 1 0 2532 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_7621
timestamp 1745462530
transform 1 0 2532 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_7622
timestamp 1745462530
transform 1 0 3068 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_7623
timestamp 1745462530
transform 1 0 2516 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_7624
timestamp 1745462530
transform 1 0 3468 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_7625
timestamp 1745462530
transform 1 0 3092 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_7626
timestamp 1745462530
transform 1 0 3092 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_7627
timestamp 1745462530
transform 1 0 3076 0 1 1955
box -2 -2 2 2
use M2_M1  M2_M1_7628
timestamp 1745462530
transform 1 0 3108 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_7629
timestamp 1745462530
transform 1 0 3044 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_7630
timestamp 1745462530
transform 1 0 3588 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_7631
timestamp 1745462530
transform 1 0 3500 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_7632
timestamp 1745462530
transform 1 0 3316 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_7633
timestamp 1745462530
transform 1 0 2516 0 1 1995
box -2 -2 2 2
use M2_M1  M2_M1_7634
timestamp 1745462530
transform 1 0 2564 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_7635
timestamp 1745462530
transform 1 0 2548 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_7636
timestamp 1745462530
transform 1 0 2476 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_7637
timestamp 1745462530
transform 1 0 2468 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_7638
timestamp 1745462530
transform 1 0 2452 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_7639
timestamp 1745462530
transform 1 0 2444 0 1 1145
box -2 -2 2 2
use M2_M1  M2_M1_7640
timestamp 1745462530
transform 1 0 2484 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_7641
timestamp 1745462530
transform 1 0 2380 0 1 1004
box -2 -2 2 2
use M2_M1  M2_M1_7642
timestamp 1745462530
transform 1 0 2484 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_7643
timestamp 1745462530
transform 1 0 2388 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_7644
timestamp 1745462530
transform 1 0 2484 0 1 1545
box -2 -2 2 2
use M2_M1  M2_M1_7645
timestamp 1745462530
transform 1 0 2444 0 1 1004
box -2 -2 2 2
use M2_M1  M2_M1_7646
timestamp 1745462530
transform 1 0 2532 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_7647
timestamp 1745462530
transform 1 0 2492 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_7648
timestamp 1745462530
transform 1 0 2628 0 1 3115
box -2 -2 2 2
use M2_M1  M2_M1_7649
timestamp 1745462530
transform 1 0 2588 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_7650
timestamp 1745462530
transform 1 0 2388 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_7651
timestamp 1745462530
transform 1 0 2388 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_7652
timestamp 1745462530
transform 1 0 4060 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_7653
timestamp 1745462530
transform 1 0 2356 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_7654
timestamp 1745462530
transform 1 0 2332 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_7655
timestamp 1745462530
transform 1 0 1676 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_7656
timestamp 1745462530
transform 1 0 1644 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_7657
timestamp 1745462530
transform 1 0 1084 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_7658
timestamp 1745462530
transform 1 0 1652 0 1 1845
box -2 -2 2 2
use M2_M1  M2_M1_7659
timestamp 1745462530
transform 1 0 1652 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_7660
timestamp 1745462530
transform 1 0 1636 0 1 1845
box -2 -2 2 2
use M2_M1  M2_M1_7661
timestamp 1745462530
transform 1 0 548 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_7662
timestamp 1745462530
transform 1 0 1748 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_7663
timestamp 1745462530
transform 1 0 1708 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_7664
timestamp 1745462530
transform 1 0 1692 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_7665
timestamp 1745462530
transform 1 0 1676 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7666
timestamp 1745462530
transform 1 0 1660 0 1 855
box -2 -2 2 2
use M2_M1  M2_M1_7667
timestamp 1745462530
transform 1 0 1644 0 1 1145
box -2 -2 2 2
use M2_M1  M2_M1_7668
timestamp 1745462530
transform 1 0 1732 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7669
timestamp 1745462530
transform 1 0 1708 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_7670
timestamp 1745462530
transform 1 0 1652 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_7671
timestamp 1745462530
transform 1 0 1636 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_7672
timestamp 1745462530
transform 1 0 1724 0 1 1545
box -2 -2 2 2
use M2_M1  M2_M1_7673
timestamp 1745462530
transform 1 0 1716 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_7674
timestamp 1745462530
transform 1 0 1748 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_7675
timestamp 1745462530
transform 1 0 1748 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_7676
timestamp 1745462530
transform 1 0 572 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_7677
timestamp 1745462530
transform 1 0 564 0 1 2195
box -2 -2 2 2
use M2_M1  M2_M1_7678
timestamp 1745462530
transform 1 0 580 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_7679
timestamp 1745462530
transform 1 0 524 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_7680
timestamp 1745462530
transform 1 0 636 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_7681
timestamp 1745462530
transform 1 0 564 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_7682
timestamp 1745462530
transform 1 0 1020 0 1 1945
box -2 -2 2 2
use M2_M1  M2_M1_7683
timestamp 1745462530
transform 1 0 924 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_7684
timestamp 1745462530
transform 1 0 1052 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_7685
timestamp 1745462530
transform 1 0 1036 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_7686
timestamp 1745462530
transform 1 0 4036 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_7687
timestamp 1745462530
transform 1 0 3996 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_7688
timestamp 1745462530
transform 1 0 4044 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7689
timestamp 1745462530
transform 1 0 4036 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_7690
timestamp 1745462530
transform 1 0 4084 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_7691
timestamp 1745462530
transform 1 0 4076 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_7692
timestamp 1745462530
transform 1 0 4092 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_7693
timestamp 1745462530
transform 1 0 4068 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_7694
timestamp 1745462530
transform 1 0 4148 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_7695
timestamp 1745462530
transform 1 0 4084 0 1 2545
box -2 -2 2 2
use M2_M1  M2_M1_7696
timestamp 1745462530
transform 1 0 4100 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_7697
timestamp 1745462530
transform 1 0 4012 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_7698
timestamp 1745462530
transform 1 0 4140 0 1 2515
box -2 -2 2 2
use M2_M1  M2_M1_7699
timestamp 1745462530
transform 1 0 4124 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_7700
timestamp 1745462530
transform 1 0 4116 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_7701
timestamp 1745462530
transform 1 0 4076 0 1 2345
box -2 -2 2 2
use M2_M1  M2_M1_7702
timestamp 1745462530
transform 1 0 4092 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_7703
timestamp 1745462530
transform 1 0 3012 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_7704
timestamp 1745462530
transform 1 0 4028 0 1 1145
box -2 -2 2 2
use M2_M1  M2_M1_7705
timestamp 1745462530
transform 1 0 4020 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_7706
timestamp 1745462530
transform 1 0 4060 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_7707
timestamp 1745462530
transform 1 0 3948 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7708
timestamp 1745462530
transform 1 0 4004 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_7709
timestamp 1745462530
transform 1 0 3924 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_7710
timestamp 1745462530
transform 1 0 3996 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_7711
timestamp 1745462530
transform 1 0 3980 0 1 1345
box -2 -2 2 2
use M2_M1  M2_M1_7712
timestamp 1745462530
transform 1 0 3996 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_7713
timestamp 1745462530
transform 1 0 3916 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_7714
timestamp 1745462530
transform 1 0 3148 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_7715
timestamp 1745462530
transform 1 0 2292 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_7716
timestamp 1745462530
transform 1 0 2284 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_7717
timestamp 1745462530
transform 1 0 2004 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_7718
timestamp 1745462530
transform 1 0 2028 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_7719
timestamp 1745462530
transform 1 0 1988 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_7720
timestamp 1745462530
transform 1 0 2084 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_7721
timestamp 1745462530
transform 1 0 1996 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_7722
timestamp 1745462530
transform 1 0 2052 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_7723
timestamp 1745462530
transform 1 0 1012 0 1 1395
box -2 -2 2 2
use M2_M1  M2_M1_7724
timestamp 1745462530
transform 1 0 2012 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_7725
timestamp 1745462530
transform 1 0 596 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_7726
timestamp 1745462530
transform 1 0 676 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_7727
timestamp 1745462530
transform 1 0 556 0 1 1195
box -2 -2 2 2
use M2_M1  M2_M1_7728
timestamp 1745462530
transform 1 0 588 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7729
timestamp 1745462530
transform 1 0 524 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_7730
timestamp 1745462530
transform 1 0 660 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_7731
timestamp 1745462530
transform 1 0 588 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_7732
timestamp 1745462530
transform 1 0 972 0 1 1395
box -2 -2 2 2
use M2_M1  M2_M1_7733
timestamp 1745462530
transform 1 0 884 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_7734
timestamp 1745462530
transform 1 0 988 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_7735
timestamp 1745462530
transform 1 0 964 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_7736
timestamp 1745462530
transform 1 0 2076 0 1 2395
box -2 -2 2 2
use M2_M1  M2_M1_7737
timestamp 1745462530
transform 1 0 2068 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_7738
timestamp 1745462530
transform 1 0 2124 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_7739
timestamp 1745462530
transform 1 0 2044 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_7740
timestamp 1745462530
transform 1 0 2060 0 1 2515
box -2 -2 2 2
use M2_M1  M2_M1_7741
timestamp 1745462530
transform 1 0 1964 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_7742
timestamp 1745462530
transform 1 0 2052 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_7743
timestamp 1745462530
transform 1 0 2044 0 1 1945
box -2 -2 2 2
use M2_M1  M2_M1_7744
timestamp 1745462530
transform 1 0 2076 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_7745
timestamp 1745462530
transform 1 0 2060 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_7746
timestamp 1745462530
transform 1 0 3180 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_7747
timestamp 1745462530
transform 1 0 3116 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_7748
timestamp 1745462530
transform 1 0 3180 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7749
timestamp 1745462530
transform 1 0 3140 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_7750
timestamp 1745462530
transform 1 0 3164 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_7751
timestamp 1745462530
transform 1 0 3132 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_7752
timestamp 1745462530
transform 1 0 3948 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_7753
timestamp 1745462530
transform 1 0 3180 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_7754
timestamp 1745462530
transform 1 0 4020 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_7755
timestamp 1745462530
transform 1 0 3964 0 1 2145
box -2 -2 2 2
use M2_M1  M2_M1_7756
timestamp 1745462530
transform 1 0 3980 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_7757
timestamp 1745462530
transform 1 0 3924 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_7758
timestamp 1745462530
transform 1 0 4060 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_7759
timestamp 1745462530
transform 1 0 4036 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_7760
timestamp 1745462530
transform 1 0 3956 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_7761
timestamp 1745462530
transform 1 0 3092 0 1 1995
box -2 -2 2 2
use M2_M1  M2_M1_7762
timestamp 1745462530
transform 1 0 3132 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_7763
timestamp 1745462530
transform 1 0 3116 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_7764
timestamp 1745462530
transform 1 0 3172 0 1 1145
box -2 -2 2 2
use M2_M1  M2_M1_7765
timestamp 1745462530
transform 1 0 3172 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_7766
timestamp 1745462530
transform 1 0 3188 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_7767
timestamp 1745462530
transform 1 0 3148 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7768
timestamp 1745462530
transform 1 0 3140 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_7769
timestamp 1745462530
transform 1 0 2972 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_7770
timestamp 1745462530
transform 1 0 3132 0 1 1345
box -2 -2 2 2
use M2_M1  M2_M1_7771
timestamp 1745462530
transform 1 0 3052 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_7772
timestamp 1745462530
transform 1 0 3172 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_7773
timestamp 1745462530
transform 1 0 3156 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_7774
timestamp 1745462530
transform 1 0 2284 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_7775
timestamp 1745462530
transform 1 0 2260 0 1 1745
box -2 -2 2 2
use M2_M1  M2_M1_7776
timestamp 1745462530
transform 1 0 2316 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_7777
timestamp 1745462530
transform 1 0 2284 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_7778
timestamp 1745462530
transform 1 0 4068 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_7779
timestamp 1745462530
transform 1 0 2292 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_7780
timestamp 1745462530
transform 1 0 2300 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_7781
timestamp 1745462530
transform 1 0 1804 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_7782
timestamp 1745462530
transform 1 0 1756 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_7783
timestamp 1745462530
transform 1 0 988 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_7784
timestamp 1745462530
transform 1 0 1796 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_7785
timestamp 1745462530
transform 1 0 676 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_7786
timestamp 1745462530
transform 1 0 1836 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_7787
timestamp 1745462530
transform 1 0 1836 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_7788
timestamp 1745462530
transform 1 0 1812 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_7789
timestamp 1745462530
transform 1 0 1812 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_7790
timestamp 1745462530
transform 1 0 1812 0 1 1395
box -2 -2 2 2
use M2_M1  M2_M1_7791
timestamp 1745462530
transform 1 0 1812 0 1 1155
box -2 -2 2 2
use M2_M1  M2_M1_7792
timestamp 1745462530
transform 1 0 1796 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_7793
timestamp 1745462530
transform 1 0 1772 0 1 1145
box -2 -2 2 2
use M2_M1  M2_M1_7794
timestamp 1745462530
transform 1 0 1836 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7795
timestamp 1745462530
transform 1 0 1812 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_7796
timestamp 1745462530
transform 1 0 1804 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_7797
timestamp 1745462530
transform 1 0 1756 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_7798
timestamp 1745462530
transform 1 0 1860 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_7799
timestamp 1745462530
transform 1 0 1820 0 1 1545
box -2 -2 2 2
use M2_M1  M2_M1_7800
timestamp 1745462530
transform 1 0 1916 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_7801
timestamp 1745462530
transform 1 0 1892 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_7802
timestamp 1745462530
transform 1 0 668 0 1 1995
box -2 -2 2 2
use M2_M1  M2_M1_7803
timestamp 1745462530
transform 1 0 620 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_7804
timestamp 1745462530
transform 1 0 684 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_7805
timestamp 1745462530
transform 1 0 596 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_7806
timestamp 1745462530
transform 1 0 604 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_7807
timestamp 1745462530
transform 1 0 596 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_7808
timestamp 1745462530
transform 1 0 956 0 1 1595
box -2 -2 2 2
use M2_M1  M2_M1_7809
timestamp 1745462530
transform 1 0 900 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_7810
timestamp 1745462530
transform 1 0 1020 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_7811
timestamp 1745462530
transform 1 0 940 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_7812
timestamp 1745462530
transform 1 0 4052 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_7813
timestamp 1745462530
transform 1 0 4052 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_7814
timestamp 1745462530
transform 1 0 4060 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_7815
timestamp 1745462530
transform 1 0 4060 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7816
timestamp 1745462530
transform 1 0 4084 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_7817
timestamp 1745462530
transform 1 0 4052 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_7818
timestamp 1745462530
transform 1 0 4092 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_7819
timestamp 1745462530
transform 1 0 4068 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_7820
timestamp 1745462530
transform 1 0 4108 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_7821
timestamp 1745462530
transform 1 0 4052 0 1 2395
box -2 -2 2 2
use M2_M1  M2_M1_7822
timestamp 1745462530
transform 1 0 4068 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_7823
timestamp 1745462530
transform 1 0 4004 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_7824
timestamp 1745462530
transform 1 0 4132 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_7825
timestamp 1745462530
transform 1 0 4132 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_7826
timestamp 1745462530
transform 1 0 4108 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_7827
timestamp 1745462530
transform 1 0 4060 0 1 2195
box -2 -2 2 2
use M2_M1  M2_M1_7828
timestamp 1745462530
transform 1 0 4076 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_7829
timestamp 1745462530
transform 1 0 2948 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_7830
timestamp 1745462530
transform 1 0 4068 0 1 1145
box -2 -2 2 2
use M2_M1  M2_M1_7831
timestamp 1745462530
transform 1 0 4060 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_7832
timestamp 1745462530
transform 1 0 4084 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_7833
timestamp 1745462530
transform 1 0 3996 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7834
timestamp 1745462530
transform 1 0 4060 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_7835
timestamp 1745462530
transform 1 0 3860 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_7836
timestamp 1745462530
transform 1 0 4060 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_7837
timestamp 1745462530
transform 1 0 4012 0 1 1345
box -2 -2 2 2
use M2_M1  M2_M1_7838
timestamp 1745462530
transform 1 0 4036 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_7839
timestamp 1745462530
transform 1 0 3972 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_7840
timestamp 1745462530
transform 1 0 2284 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_7841
timestamp 1745462530
transform 1 0 2260 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_7842
timestamp 1745462530
transform 1 0 2268 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_7843
timestamp 1745462530
transform 1 0 1572 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_7844
timestamp 1745462530
transform 1 0 1556 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_7845
timestamp 1745462530
transform 1 0 1556 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_7846
timestamp 1745462530
transform 1 0 1620 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_7847
timestamp 1745462530
transform 1 0 1532 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_7848
timestamp 1745462530
transform 1 0 1588 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_7849
timestamp 1745462530
transform 1 0 1012 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_7850
timestamp 1745462530
transform 1 0 1580 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_7851
timestamp 1745462530
transform 1 0 668 0 1 1145
box -2 -2 2 2
use M2_M1  M2_M1_7852
timestamp 1745462530
transform 1 0 612 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_7853
timestamp 1745462530
transform 1 0 604 0 1 1145
box -2 -2 2 2
use M2_M1  M2_M1_7854
timestamp 1745462530
transform 1 0 644 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_7855
timestamp 1745462530
transform 1 0 580 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7856
timestamp 1745462530
transform 1 0 596 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_7857
timestamp 1745462530
transform 1 0 524 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_7858
timestamp 1745462530
transform 1 0 996 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_7859
timestamp 1745462530
transform 1 0 980 0 1 1545
box -2 -2 2 2
use M2_M1  M2_M1_7860
timestamp 1745462530
transform 1 0 1020 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_7861
timestamp 1745462530
transform 1 0 996 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_7862
timestamp 1745462530
transform 1 0 1652 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_7863
timestamp 1745462530
transform 1 0 1596 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_7864
timestamp 1745462530
transform 1 0 1644 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_7865
timestamp 1745462530
transform 1 0 1620 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_7866
timestamp 1745462530
transform 1 0 1676 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_7867
timestamp 1745462530
transform 1 0 1644 0 1 2715
box -2 -2 2 2
use M2_M1  M2_M1_7868
timestamp 1745462530
transform 1 0 1652 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_7869
timestamp 1745462530
transform 1 0 1580 0 1 1745
box -2 -2 2 2
use M2_M1  M2_M1_7870
timestamp 1745462530
transform 1 0 1604 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_7871
timestamp 1745462530
transform 1 0 1572 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_7872
timestamp 1745462530
transform 1 0 2268 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_7873
timestamp 1745462530
transform 1 0 2268 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_7874
timestamp 1745462530
transform 1 0 2276 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_7875
timestamp 1745462530
transform 1 0 2268 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_7876
timestamp 1745462530
transform 1 0 2612 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_7877
timestamp 1745462530
transform 1 0 2300 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_7878
timestamp 1745462530
transform 1 0 2916 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_7879
timestamp 1745462530
transform 1 0 2292 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_7880
timestamp 1745462530
transform 1 0 3268 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_7881
timestamp 1745462530
transform 1 0 2948 0 1 1545
box -2 -2 2 2
use M2_M1  M2_M1_7882
timestamp 1745462530
transform 1 0 3020 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_7883
timestamp 1745462530
transform 1 0 2996 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_7884
timestamp 1745462530
transform 1 0 3404 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_7885
timestamp 1745462530
transform 1 0 3300 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_7886
timestamp 1745462530
transform 1 0 3212 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_7887
timestamp 1745462530
transform 1 0 2604 0 1 1595
box -2 -2 2 2
use M2_M1  M2_M1_7888
timestamp 1745462530
transform 1 0 2628 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_7889
timestamp 1745462530
transform 1 0 2620 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_7890
timestamp 1745462530
transform 1 0 2276 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_7891
timestamp 1745462530
transform 1 0 2244 0 1 995
box -2 -2 2 2
use M2_M1  M2_M1_7892
timestamp 1745462530
transform 1 0 2276 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7893
timestamp 1745462530
transform 1 0 2212 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_7894
timestamp 1745462530
transform 1 0 2284 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_7895
timestamp 1745462530
transform 1 0 2236 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_7896
timestamp 1745462530
transform 1 0 2340 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_7897
timestamp 1745462530
transform 1 0 2260 0 1 1395
box -2 -2 2 2
use M2_M1  M2_M1_7898
timestamp 1745462530
transform 1 0 2348 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_7899
timestamp 1745462530
transform 1 0 2308 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_7900
timestamp 1745462530
transform 1 0 2396 0 1 1745
box -2 -2 2 2
use M2_M1  M2_M1_7901
timestamp 1745462530
transform 1 0 2396 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_7902
timestamp 1745462530
transform 1 0 2412 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_7903
timestamp 1745462530
transform 1 0 2388 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_7904
timestamp 1745462530
transform 1 0 3148 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_7905
timestamp 1745462530
transform 1 0 2348 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_7906
timestamp 1745462530
transform 1 0 2324 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_7907
timestamp 1745462530
transform 1 0 1460 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_7908
timestamp 1745462530
transform 1 0 1436 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_7909
timestamp 1745462530
transform 1 0 1076 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_7910
timestamp 1745462530
transform 1 0 1452 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_7911
timestamp 1745462530
transform 1 0 716 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_7912
timestamp 1745462530
transform 1 0 1476 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_7913
timestamp 1745462530
transform 1 0 1476 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_7914
timestamp 1745462530
transform 1 0 1524 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7915
timestamp 1745462530
transform 1 0 1508 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_7916
timestamp 1745462530
transform 1 0 1524 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_7917
timestamp 1745462530
transform 1 0 1508 0 1 1145
box -2 -2 2 2
use M2_M1  M2_M1_7918
timestamp 1745462530
transform 1 0 1540 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_7919
timestamp 1745462530
transform 1 0 1540 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_7920
timestamp 1745462530
transform 1 0 1532 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_7921
timestamp 1745462530
transform 1 0 1380 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_7922
timestamp 1745462530
transform 1 0 1452 0 1 1545
box -2 -2 2 2
use M2_M1  M2_M1_7923
timestamp 1745462530
transform 1 0 1420 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_7924
timestamp 1745462530
transform 1 0 1532 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_7925
timestamp 1745462530
transform 1 0 1492 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_7926
timestamp 1745462530
transform 1 0 668 0 1 2345
box -2 -2 2 2
use M2_M1  M2_M1_7927
timestamp 1745462530
transform 1 0 644 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_7928
timestamp 1745462530
transform 1 0 700 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_7929
timestamp 1745462530
transform 1 0 644 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_7930
timestamp 1745462530
transform 1 0 644 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_7931
timestamp 1745462530
transform 1 0 596 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_7932
timestamp 1745462530
transform 1 0 1060 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_7933
timestamp 1745462530
transform 1 0 1052 0 1 1795
box -2 -2 2 2
use M2_M1  M2_M1_7934
timestamp 1745462530
transform 1 0 1084 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_7935
timestamp 1745462530
transform 1 0 1060 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_7936
timestamp 1745462530
transform 1 0 3180 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_7937
timestamp 1745462530
transform 1 0 3116 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_7938
timestamp 1745462530
transform 1 0 3204 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_7939
timestamp 1745462530
transform 1 0 3108 0 1 1745
box -2 -2 2 2
use M2_M1  M2_M1_7940
timestamp 1745462530
transform 1 0 3076 0 1 1555
box -2 -2 2 2
use M2_M1  M2_M1_7941
timestamp 1745462530
transform 1 0 3044 0 1 1505
box -2 -2 2 2
use M2_M1  M2_M1_7942
timestamp 1745462530
transform 1 0 3172 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_7943
timestamp 1745462530
transform 1 0 3164 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_7944
timestamp 1745462530
transform 1 0 3156 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_7945
timestamp 1745462530
transform 1 0 3140 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_7946
timestamp 1745462530
transform 1 0 3132 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_7947
timestamp 1745462530
transform 1 0 3108 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_7948
timestamp 1745462530
transform 1 0 3236 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_7949
timestamp 1745462530
transform 1 0 3132 0 1 2545
box -2 -2 2 2
use M2_M1  M2_M1_7950
timestamp 1745462530
transform 1 0 3148 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_7951
timestamp 1745462530
transform 1 0 3084 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_7952
timestamp 1745462530
transform 1 0 3244 0 1 2515
box -2 -2 2 2
use M2_M1  M2_M1_7953
timestamp 1745462530
transform 1 0 3228 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_7954
timestamp 1745462530
transform 1 0 3220 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_7955
timestamp 1745462530
transform 1 0 3148 0 1 1995
box -2 -2 2 2
use M2_M1  M2_M1_7956
timestamp 1745462530
transform 1 0 3180 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_7957
timestamp 1745462530
transform 1 0 2780 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_7958
timestamp 1745462530
transform 1 0 3316 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_7959
timestamp 1745462530
transform 1 0 3204 0 1 995
box -2 -2 2 2
use M2_M1  M2_M1_7960
timestamp 1745462530
transform 1 0 3228 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7961
timestamp 1745462530
transform 1 0 3116 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_7962
timestamp 1745462530
transform 1 0 3308 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_7963
timestamp 1745462530
transform 1 0 3220 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_7964
timestamp 1745462530
transform 1 0 3204 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_7965
timestamp 1745462530
transform 1 0 3148 0 1 1195
box -2 -2 2 2
use M2_M1  M2_M1_7966
timestamp 1745462530
transform 1 0 3172 0 1 1245
box -2 -2 2 2
use M2_M1  M2_M1_7967
timestamp 1745462530
transform 1 0 3148 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_7968
timestamp 1745462530
transform 1 0 3052 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_7969
timestamp 1745462530
transform 1 0 2364 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_7970
timestamp 1745462530
transform 1 0 2356 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_7971
timestamp 1745462530
transform 1 0 1164 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_7972
timestamp 1745462530
transform 1 0 1244 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_7973
timestamp 1745462530
transform 1 0 1148 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_7974
timestamp 1745462530
transform 1 0 1332 0 1 2595
box -2 -2 2 2
use M2_M1  M2_M1_7975
timestamp 1745462530
transform 1 0 1156 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_7976
timestamp 1745462530
transform 1 0 1188 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_7977
timestamp 1745462530
transform 1 0 1100 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_7978
timestamp 1745462530
transform 1 0 1172 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_7979
timestamp 1745462530
transform 1 0 628 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_7980
timestamp 1745462530
transform 1 0 644 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_7981
timestamp 1745462530
transform 1 0 620 0 1 995
box -2 -2 2 2
use M2_M1  M2_M1_7982
timestamp 1745462530
transform 1 0 652 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7983
timestamp 1745462530
transform 1 0 588 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_7984
timestamp 1745462530
transform 1 0 644 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_7985
timestamp 1745462530
transform 1 0 588 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_7986
timestamp 1745462530
transform 1 0 1060 0 1 1395
box -2 -2 2 2
use M2_M1  M2_M1_7987
timestamp 1745462530
transform 1 0 1060 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_7988
timestamp 1745462530
transform 1 0 1076 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_7989
timestamp 1745462530
transform 1 0 1052 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_7990
timestamp 1745462530
transform 1 0 1364 0 1 2705
box -2 -2 2 2
use M2_M1  M2_M1_7991
timestamp 1745462530
transform 1 0 1308 0 1 2595
box -2 -2 2 2
use M2_M1  M2_M1_7992
timestamp 1745462530
transform 1 0 1356 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_7993
timestamp 1745462530
transform 1 0 1332 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_7994
timestamp 1745462530
transform 1 0 1356 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_7995
timestamp 1745462530
transform 1 0 1356 0 1 2715
box -2 -2 2 2
use M2_M1  M2_M1_7996
timestamp 1745462530
transform 1 0 1324 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_7997
timestamp 1745462530
transform 1 0 1260 0 1 1595
box -2 -2 2 2
use M2_M1  M2_M1_7998
timestamp 1745462530
transform 1 0 1276 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_7999
timestamp 1745462530
transform 1 0 1276 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_8000
timestamp 1745462530
transform 1 0 3028 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_8001
timestamp 1745462530
transform 1 0 3028 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_8002
timestamp 1745462530
transform 1 0 3060 0 1 1145
box -2 -2 2 2
use M2_M1  M2_M1_8003
timestamp 1745462530
transform 1 0 3012 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_8004
timestamp 1745462530
transform 1 0 3068 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_8005
timestamp 1745462530
transform 1 0 2972 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_8006
timestamp 1745462530
transform 1 0 3188 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_8007
timestamp 1745462530
transform 1 0 3108 0 1 1395
box -2 -2 2 2
use M2_M1  M2_M1_8008
timestamp 1745462530
transform 1 0 3132 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_8009
timestamp 1745462530
transform 1 0 3100 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_8010
timestamp 1745462530
transform 1 0 3324 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_8011
timestamp 1745462530
transform 1 0 3212 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_8012
timestamp 1745462530
transform 1 0 3132 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_8013
timestamp 1745462530
transform 1 0 2956 0 1 1595
box -2 -2 2 2
use M2_M1  M2_M1_8014
timestamp 1745462530
transform 1 0 2980 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_8015
timestamp 1745462530
transform 1 0 2964 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_8016
timestamp 1745462530
transform 1 0 3044 0 1 1145
box -2 -2 2 2
use M2_M1  M2_M1_8017
timestamp 1745462530
transform 1 0 3036 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8018
timestamp 1745462530
transform 1 0 3083 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_8019
timestamp 1745462530
transform 1 0 3060 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_8020
timestamp 1745462530
transform 1 0 2444 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_8021
timestamp 1745462530
transform 1 0 2436 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_8022
timestamp 1745462530
transform 1 0 2428 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_8023
timestamp 1745462530
transform 1 0 2460 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_8024
timestamp 1745462530
transform 1 0 2436 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_8025
timestamp 1745462530
transform 1 0 3036 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_8026
timestamp 1745462530
transform 1 0 2892 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_8027
timestamp 1745462530
transform 1 0 2492 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_8028
timestamp 1745462530
transform 1 0 2428 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_8029
timestamp 1745462530
transform 1 0 2412 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_8030
timestamp 1745462530
transform 1 0 2388 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_8031
timestamp 1745462530
transform 1 0 2388 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_8032
timestamp 1745462530
transform 1 0 2372 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_8033
timestamp 1745462530
transform 1 0 3116 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_8034
timestamp 1745462530
transform 1 0 3052 0 1 1345
box -2 -2 2 2
use M2_M1  M2_M1_8035
timestamp 1745462530
transform 1 0 3068 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_8036
timestamp 1745462530
transform 1 0 3044 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_8037
timestamp 1745462530
transform 1 0 2228 0 1 3825
box -2 -2 2 2
use M2_M1  M2_M1_8038
timestamp 1745462530
transform 1 0 2172 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_8039
timestamp 1745462530
transform 1 0 2380 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_8040
timestamp 1745462530
transform 1 0 2212 0 1 3835
box -2 -2 2 2
use M2_M1  M2_M1_8041
timestamp 1745462530
transform 1 0 2732 0 1 3825
box -2 -2 2 2
use M2_M1  M2_M1_8042
timestamp 1745462530
transform 1 0 2356 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_8043
timestamp 1745462530
transform 1 0 2004 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_8044
timestamp 1745462530
transform 1 0 1596 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_8045
timestamp 1745462530
transform 1 0 1164 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_8046
timestamp 1745462530
transform 1 0 2308 0 1 3825
box -2 -2 2 2
use M2_M1  M2_M1_8047
timestamp 1745462530
transform 1 0 2132 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_8048
timestamp 1745462530
transform 1 0 3476 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_8049
timestamp 1745462530
transform 1 0 2332 0 1 3835
box -2 -2 2 2
use M2_M1  M2_M1_8050
timestamp 1745462530
transform 1 0 3580 0 1 3715
box -2 -2 2 2
use M2_M1  M2_M1_8051
timestamp 1745462530
transform 1 0 3468 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_8052
timestamp 1745462530
transform 1 0 3484 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_8053
timestamp 1745462530
transform 1 0 3468 0 1 3825
box -2 -2 2 2
use M2_M1  M2_M1_8054
timestamp 1745462530
transform 1 0 3444 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_8055
timestamp 1745462530
transform 1 0 3436 0 1 3825
box -2 -2 2 2
use M2_M1  M2_M1_8056
timestamp 1745462530
transform 1 0 3444 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_8057
timestamp 1745462530
transform 1 0 3260 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_8058
timestamp 1745462530
transform 1 0 3924 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_8059
timestamp 1745462530
transform 1 0 3452 0 1 3835
box -2 -2 2 2
use M2_M1  M2_M1_8060
timestamp 1745462530
transform 1 0 3988 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_8061
timestamp 1745462530
transform 1 0 3940 0 1 3795
box -2 -2 2 2
use M2_M1  M2_M1_8062
timestamp 1745462530
transform 1 0 4044 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_8063
timestamp 1745462530
transform 1 0 3964 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_8064
timestamp 1745462530
transform 1 0 4236 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_8065
timestamp 1745462530
transform 1 0 4164 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_8066
timestamp 1745462530
transform 1 0 4156 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_8067
timestamp 1745462530
transform 1 0 4036 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_8068
timestamp 1745462530
transform 1 0 1732 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_8069
timestamp 1745462530
transform 1 0 1724 0 1 3625
box -2 -2 2 2
use M2_M1  M2_M1_8070
timestamp 1745462530
transform 1 0 4252 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_8071
timestamp 1745462530
transform 1 0 4180 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_8072
timestamp 1745462530
transform 1 0 4172 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_8073
timestamp 1745462530
transform 1 0 4052 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_8074
timestamp 1745462530
transform 1 0 1868 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_8075
timestamp 1745462530
transform 1 0 1868 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_8076
timestamp 1745462530
transform 1 0 4084 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_8077
timestamp 1745462530
transform 1 0 4084 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_8078
timestamp 1745462530
transform 1 0 4052 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_8079
timestamp 1745462530
transform 1 0 3980 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_8080
timestamp 1745462530
transform 1 0 2468 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_8081
timestamp 1745462530
transform 1 0 1932 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_8082
timestamp 1745462530
transform 1 0 4124 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_8083
timestamp 1745462530
transform 1 0 4100 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_8084
timestamp 1745462530
transform 1 0 4068 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_8085
timestamp 1745462530
transform 1 0 3996 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_8086
timestamp 1745462530
transform 1 0 2492 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_8087
timestamp 1745462530
transform 1 0 1684 0 1 3715
box -2 -2 2 2
use M2_M1  M2_M1_8088
timestamp 1745462530
transform 1 0 1908 0 1 3145
box -2 -2 2 2
use M2_M1  M2_M1_8089
timestamp 1745462530
transform 1 0 1868 0 1 3145
box -2 -2 2 2
use M2_M1  M2_M1_8090
timestamp 1745462530
transform 1 0 1652 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_8091
timestamp 1745462530
transform 1 0 1644 0 1 3225
box -2 -2 2 2
use M2_M1  M2_M1_8092
timestamp 1745462530
transform 1 0 3564 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_8093
timestamp 1745462530
transform 1 0 3556 0 1 3715
box -2 -2 2 2
use M2_M1  M2_M1_8094
timestamp 1745462530
transform 1 0 3564 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_8095
timestamp 1745462530
transform 1 0 3540 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_8096
timestamp 1745462530
transform 1 0 3996 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_8097
timestamp 1745462530
transform 1 0 3572 0 1 3705
box -2 -2 2 2
use M2_M1  M2_M1_8098
timestamp 1745462530
transform 1 0 4060 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_8099
timestamp 1745462530
transform 1 0 4012 0 1 3745
box -2 -2 2 2
use M2_M1  M2_M1_8100
timestamp 1745462530
transform 1 0 4164 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_8101
timestamp 1745462530
transform 1 0 4044 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_8102
timestamp 1745462530
transform 1 0 3132 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_8103
timestamp 1745462530
transform 1 0 1708 0 1 3115
box -2 -2 2 2
use M2_M1  M2_M1_8104
timestamp 1745462530
transform 1 0 2300 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_8105
timestamp 1745462530
transform 1 0 2268 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_8106
timestamp 1745462530
transform 1 0 2276 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_8107
timestamp 1745462530
transform 1 0 2100 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_8108
timestamp 1745462530
transform 1 0 1972 0 1 3145
box -2 -2 2 2
use M2_M1  M2_M1_8109
timestamp 1745462530
transform 1 0 1956 0 1 3145
box -2 -2 2 2
use M2_M1  M2_M1_8110
timestamp 1745462530
transform 1 0 1612 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_8111
timestamp 1745462530
transform 1 0 2092 0 1 3715
box -2 -2 2 2
use M2_M1  M2_M1_8112
timestamp 1745462530
transform 1 0 1716 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_8113
timestamp 1745462530
transform 1 0 2116 0 1 3715
box -2 -2 2 2
use M2_M1  M2_M1_8114
timestamp 1745462530
transform 1 0 2068 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_8115
timestamp 1745462530
transform 1 0 2356 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_8116
timestamp 1745462530
transform 1 0 2300 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_8117
timestamp 1745462530
transform 1 0 2340 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_8118
timestamp 1745462530
transform 1 0 2324 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_8119
timestamp 1745462530
transform 1 0 2116 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_8120
timestamp 1745462530
transform 1 0 2100 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_8121
timestamp 1745462530
transform 1 0 2164 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_8122
timestamp 1745462530
transform 1 0 1532 0 1 3315
box -2 -2 2 2
use M2_M1  M2_M1_8123
timestamp 1745462530
transform 1 0 1492 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_8124
timestamp 1745462530
transform 1 0 2060 0 1 3825
box -2 -2 2 2
use M2_M1  M2_M1_8125
timestamp 1745462530
transform 1 0 1740 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_8126
timestamp 1745462530
transform 1 0 2084 0 1 3825
box -2 -2 2 2
use M2_M1  M2_M1_8127
timestamp 1745462530
transform 1 0 2036 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_8128
timestamp 1745462530
transform 1 0 2244 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_8129
timestamp 1745462530
transform 1 0 2108 0 1 4005
box -2 -2 2 2
use M2_M1  M2_M1_8130
timestamp 1745462530
transform 1 0 2172 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_8131
timestamp 1745462530
transform 1 0 2124 0 1 4025
box -2 -2 2 2
use M2_M1  M2_M1_8132
timestamp 1745462530
transform 1 0 2764 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_8133
timestamp 1745462530
transform 1 0 2716 0 1 3825
box -2 -2 2 2
use M2_M1  M2_M1_8134
timestamp 1745462530
transform 1 0 3524 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_8135
timestamp 1745462530
transform 1 0 2708 0 1 3835
box -2 -2 2 2
use M2_M1  M2_M1_8136
timestamp 1745462530
transform 1 0 3596 0 1 3825
box -2 -2 2 2
use M2_M1  M2_M1_8137
timestamp 1745462530
transform 1 0 3516 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_8138
timestamp 1745462530
transform 1 0 3532 0 1 3915
box -2 -2 2 2
use M2_M1  M2_M1_8139
timestamp 1745462530
transform 1 0 3532 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_8140
timestamp 1745462530
transform 1 0 3540 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_8141
timestamp 1745462530
transform 1 0 3508 0 1 3915
box -2 -2 2 2
use M2_M1  M2_M1_8142
timestamp 1745462530
transform 1 0 3516 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_8143
timestamp 1745462530
transform 1 0 3476 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_8144
timestamp 1745462530
transform 1 0 4116 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_8145
timestamp 1745462530
transform 1 0 3524 0 1 3905
box -2 -2 2 2
use M2_M1  M2_M1_8146
timestamp 1745462530
transform 1 0 4116 0 1 3795
box -2 -2 2 2
use M2_M1  M2_M1_8147
timestamp 1745462530
transform 1 0 4092 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_8148
timestamp 1745462530
transform 1 0 4172 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_8149
timestamp 1745462530
transform 1 0 4156 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_8150
timestamp 1745462530
transform 1 0 1636 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_8151
timestamp 1745462530
transform 1 0 1564 0 1 3315
box -2 -2 2 2
use M2_M1  M2_M1_8152
timestamp 1745462530
transform 1 0 1500 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_8153
timestamp 1745462530
transform 1 0 3580 0 1 3825
box -2 -2 2 2
use M2_M1  M2_M1_8154
timestamp 1745462530
transform 1 0 3564 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_8155
timestamp 1745462530
transform 1 0 3580 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_8156
timestamp 1745462530
transform 1 0 3492 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_8157
timestamp 1745462530
transform 1 0 4212 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_8158
timestamp 1745462530
transform 1 0 3588 0 1 3835
box -2 -2 2 2
use M2_M1  M2_M1_8159
timestamp 1745462530
transform 1 0 4196 0 1 3745
box -2 -2 2 2
use M2_M1  M2_M1_8160
timestamp 1745462530
transform 1 0 4116 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_8161
timestamp 1745462530
transform 1 0 4244 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_8162
timestamp 1745462530
transform 1 0 4228 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_8163
timestamp 1745462530
transform 1 0 2732 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_8164
timestamp 1745462530
transform 1 0 2668 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_8165
timestamp 1745462530
transform 1 0 2660 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_8166
timestamp 1745462530
transform 1 0 2524 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_8167
timestamp 1745462530
transform 1 0 2508 0 1 3825
box -2 -2 2 2
use M2_M1  M2_M1_8168
timestamp 1745462530
transform 1 0 1844 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_8169
timestamp 1745462530
transform 1 0 2556 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_8170
timestamp 1745462530
transform 1 0 2532 0 1 3825
box -2 -2 2 2
use M2_M1  M2_M1_8171
timestamp 1745462530
transform 1 0 2732 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_8172
timestamp 1745462530
transform 1 0 2684 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_8173
timestamp 1745462530
transform 1 0 2780 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_8174
timestamp 1745462530
transform 1 0 2756 0 1 3915
box -2 -2 2 2
use M2_M1  M2_M1_8175
timestamp 1745462530
transform 1 0 3004 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_8176
timestamp 1745462530
transform 1 0 2740 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_8177
timestamp 1745462530
transform 1 0 2748 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_8178
timestamp 1745462530
transform 1 0 2612 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_8179
timestamp 1745462530
transform 1 0 2572 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_8180
timestamp 1745462530
transform 1 0 1796 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_8181
timestamp 1745462530
transform 1 0 2636 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_8182
timestamp 1745462530
transform 1 0 2612 0 1 3825
box -2 -2 2 2
use M2_M1  M2_M1_8183
timestamp 1745462530
transform 1 0 1908 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_8184
timestamp 1745462530
transform 1 0 1860 0 1 3745
box -2 -2 2 2
use M2_M1  M2_M1_8185
timestamp 1745462530
transform 1 0 1652 0 1 3715
box -2 -2 2 2
use M2_M1  M2_M1_8186
timestamp 1745462530
transform 1 0 1652 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_8187
timestamp 1745462530
transform 1 0 1788 0 1 3745
box -2 -2 2 2
use M2_M1  M2_M1_8188
timestamp 1745462530
transform 1 0 1772 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_8189
timestamp 1745462530
transform 1 0 1756 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_8190
timestamp 1745462530
transform 1 0 1628 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_8191
timestamp 1745462530
transform 1 0 1628 0 1 3625
box -2 -2 2 2
use M2_M1  M2_M1_8192
timestamp 1745462530
transform 1 0 3060 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_8193
timestamp 1745462530
transform 1 0 2996 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_8194
timestamp 1745462530
transform 1 0 3052 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_8195
timestamp 1745462530
transform 1 0 3012 0 1 3915
box -2 -2 2 2
use M2_M1  M2_M1_8196
timestamp 1745462530
transform 1 0 1820 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_8197
timestamp 1745462530
transform 1 0 1612 0 1 3625
box -2 -2 2 2
use M2_M1  M2_M1_8198
timestamp 1745462530
transform 1 0 1428 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_8199
timestamp 1745462530
transform 1 0 2068 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_8200
timestamp 1745462530
transform 1 0 1572 0 1 3625
box -2 -2 2 2
use M2_M1  M2_M1_8201
timestamp 1745462530
transform 1 0 1540 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_8202
timestamp 1745462530
transform 1 0 988 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_8203
timestamp 1745462530
transform 1 0 956 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_8204
timestamp 1745462530
transform 1 0 1108 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_8205
timestamp 1745462530
transform 1 0 1068 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_8206
timestamp 1745462530
transform 1 0 988 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_8207
timestamp 1745462530
transform 1 0 844 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_8208
timestamp 1745462530
transform 1 0 836 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_8209
timestamp 1745462530
transform 1 0 812 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_8210
timestamp 1745462530
transform 1 0 948 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_8211
timestamp 1745462530
transform 1 0 844 0 1 3515
box -2 -2 2 2
use M2_M1  M2_M1_8212
timestamp 1745462530
transform 1 0 916 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_8213
timestamp 1745462530
transform 1 0 884 0 1 3515
box -2 -2 2 2
use M2_M1  M2_M1_8214
timestamp 1745462530
transform 1 0 1020 0 1 3625
box -2 -2 2 2
use M2_M1  M2_M1_8215
timestamp 1745462530
transform 1 0 964 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_8216
timestamp 1745462530
transform 1 0 1140 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_8217
timestamp 1745462530
transform 1 0 1132 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_8218
timestamp 1745462530
transform 1 0 908 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_8219
timestamp 1745462530
transform 1 0 876 0 1 3425
box -2 -2 2 2
use M2_M1  M2_M1_8220
timestamp 1745462530
transform 1 0 1604 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_8221
timestamp 1745462530
transform 1 0 1564 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_8222
timestamp 1745462530
transform 1 0 1428 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_8223
timestamp 1745462530
transform 1 0 1364 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_8224
timestamp 1745462530
transform 1 0 1316 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_8225
timestamp 1745462530
transform 1 0 1300 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_8226
timestamp 1745462530
transform 1 0 1292 0 1 3115
box -2 -2 2 2
use M2_M1  M2_M1_8227
timestamp 1745462530
transform 1 0 1260 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_8228
timestamp 1745462530
transform 1 0 1292 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_8229
timestamp 1745462530
transform 1 0 1276 0 1 3225
box -2 -2 2 2
use M2_M1  M2_M1_8230
timestamp 1745462530
transform 1 0 1444 0 1 3115
box -2 -2 2 2
use M2_M1  M2_M1_8231
timestamp 1745462530
transform 1 0 1420 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_8232
timestamp 1745462530
transform 1 0 1636 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_8233
timestamp 1745462530
transform 1 0 1588 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_8234
timestamp 1745462530
transform 1 0 1356 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_8235
timestamp 1745462530
transform 1 0 1332 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_8236
timestamp 1745462530
transform 1 0 1308 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_8237
timestamp 1745462530
transform 1 0 1380 0 1 3225
box -2 -2 2 2
use M2_M1  M2_M1_8238
timestamp 1745462530
transform 1 0 1356 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_8239
timestamp 1745462530
transform 1 0 1860 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_8240
timestamp 1745462530
transform 1 0 1796 0 1 2845
box -2 -2 2 2
use M2_M1  M2_M1_8241
timestamp 1745462530
transform 1 0 1732 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_8242
timestamp 1745462530
transform 1 0 1636 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_8243
timestamp 1745462530
transform 1 0 1580 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_8244
timestamp 1745462530
transform 1 0 1492 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_8245
timestamp 1745462530
transform 1 0 1292 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_8246
timestamp 1745462530
transform 1 0 1236 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_8247
timestamp 1745462530
transform 1 0 2452 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_8248
timestamp 1745462530
transform 1 0 1844 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_8249
timestamp 1745462530
transform 1 0 1836 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_8250
timestamp 1745462530
transform 1 0 1972 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_8251
timestamp 1745462530
transform 1 0 1892 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_8252
timestamp 1745462530
transform 1 0 1692 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_8253
timestamp 1745462530
transform 1 0 1636 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_8254
timestamp 1745462530
transform 1 0 1548 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_8255
timestamp 1745462530
transform 1 0 1548 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_8256
timestamp 1745462530
transform 1 0 1276 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_8257
timestamp 1745462530
transform 1 0 1220 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_8258
timestamp 1745462530
transform 1 0 1884 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_8259
timestamp 1745462530
transform 1 0 1820 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_8260
timestamp 1745462530
transform 1 0 1812 0 1 2595
box -2 -2 2 2
use M2_M1  M2_M1_8261
timestamp 1745462530
transform 1 0 1668 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_8262
timestamp 1745462530
transform 1 0 1668 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_8263
timestamp 1745462530
transform 1 0 1540 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_8264
timestamp 1745462530
transform 1 0 1484 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_8265
timestamp 1745462530
transform 1 0 1268 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_8266
timestamp 1745462530
transform 1 0 1220 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_8267
timestamp 1745462530
transform 1 0 1852 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_8268
timestamp 1745462530
transform 1 0 1812 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_8269
timestamp 1745462530
transform 1 0 1796 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_8270
timestamp 1745462530
transform 1 0 1604 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_8271
timestamp 1745462530
transform 1 0 1444 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_8272
timestamp 1745462530
transform 1 0 1420 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_8273
timestamp 1745462530
transform 1 0 1244 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_8274
timestamp 1745462530
transform 1 0 1220 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_8275
timestamp 1745462530
transform 1 0 1796 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_8276
timestamp 1745462530
transform 1 0 1732 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_8277
timestamp 1745462530
transform 1 0 1540 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_8278
timestamp 1745462530
transform 1 0 1404 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_8279
timestamp 1745462530
transform 1 0 1340 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_8280
timestamp 1745462530
transform 1 0 1260 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_8281
timestamp 1745462530
transform 1 0 1204 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_8282
timestamp 1745462530
transform 1 0 1812 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_8283
timestamp 1745462530
transform 1 0 1740 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_8284
timestamp 1745462530
transform 1 0 1580 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_8285
timestamp 1745462530
transform 1 0 1484 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_8286
timestamp 1745462530
transform 1 0 1484 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_8287
timestamp 1745462530
transform 1 0 1372 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_8288
timestamp 1745462530
transform 1 0 1364 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_8289
timestamp 1745462530
transform 1 0 1348 0 1 1945
box -2 -2 2 2
use M2_M1  M2_M1_8290
timestamp 1745462530
transform 1 0 1252 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_8291
timestamp 1745462530
transform 1 0 1180 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_8292
timestamp 1745462530
transform 1 0 1020 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_8293
timestamp 1745462530
transform 1 0 852 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_8294
timestamp 1745462530
transform 1 0 772 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_8295
timestamp 1745462530
transform 1 0 444 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_8296
timestamp 1745462530
transform 1 0 404 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_8297
timestamp 1745462530
transform 1 0 388 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_8298
timestamp 1745462530
transform 1 0 332 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_8299
timestamp 1745462530
transform 1 0 284 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_8300
timestamp 1745462530
transform 1 0 796 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_8301
timestamp 1745462530
transform 1 0 764 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_8302
timestamp 1745462530
transform 1 0 740 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_8303
timestamp 1745462530
transform 1 0 700 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_8304
timestamp 1745462530
transform 1 0 604 0 1 2524
box -2 -2 2 2
use M2_M1  M2_M1_8305
timestamp 1745462530
transform 1 0 596 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_8306
timestamp 1745462530
transform 1 0 548 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_8307
timestamp 1745462530
transform 1 0 532 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_8308
timestamp 1745462530
transform 1 0 508 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_8309
timestamp 1745462530
transform 1 0 540 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_8310
timestamp 1745462530
transform 1 0 460 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_8311
timestamp 1745462530
transform 1 0 356 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_8312
timestamp 1745462530
transform 1 0 308 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_8313
timestamp 1745462530
transform 1 0 260 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_8314
timestamp 1745462530
transform 1 0 236 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_8315
timestamp 1745462530
transform 1 0 236 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_8316
timestamp 1745462530
transform 1 0 228 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_8317
timestamp 1745462530
transform 1 0 980 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_8318
timestamp 1745462530
transform 1 0 972 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_8319
timestamp 1745462530
transform 1 0 972 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_8320
timestamp 1745462530
transform 1 0 972 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_8321
timestamp 1745462530
transform 1 0 972 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_8322
timestamp 1745462530
transform 1 0 940 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_8323
timestamp 1745462530
transform 1 0 924 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_8324
timestamp 1745462530
transform 1 0 924 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_8325
timestamp 1745462530
transform 1 0 476 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_8326
timestamp 1745462530
transform 1 0 412 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_8327
timestamp 1745462530
transform 1 0 372 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_8328
timestamp 1745462530
transform 1 0 340 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_8329
timestamp 1745462530
transform 1 0 292 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_8330
timestamp 1745462530
transform 1 0 228 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_8331
timestamp 1745462530
transform 1 0 220 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_8332
timestamp 1745462530
transform 1 0 180 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_8333
timestamp 1745462530
transform 1 0 556 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_8334
timestamp 1745462530
transform 1 0 444 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_8335
timestamp 1745462530
transform 1 0 404 0 1 1985
box -2 -2 2 2
use M2_M1  M2_M1_8336
timestamp 1745462530
transform 1 0 340 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_8337
timestamp 1745462530
transform 1 0 268 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_8338
timestamp 1745462530
transform 1 0 252 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_8339
timestamp 1745462530
transform 1 0 204 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_8340
timestamp 1745462530
transform 1 0 196 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_8341
timestamp 1745462530
transform 1 0 668 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_8342
timestamp 1745462530
transform 1 0 396 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_8343
timestamp 1745462530
transform 1 0 396 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_8344
timestamp 1745462530
transform 1 0 316 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_8345
timestamp 1745462530
transform 1 0 244 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_8346
timestamp 1745462530
transform 1 0 228 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_8347
timestamp 1745462530
transform 1 0 212 0 1 1785
box -2 -2 2 2
use M2_M1  M2_M1_8348
timestamp 1745462530
transform 1 0 204 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_8349
timestamp 1745462530
transform 1 0 180 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_8350
timestamp 1745462530
transform 1 0 172 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_8351
timestamp 1745462530
transform 1 0 740 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_8352
timestamp 1745462530
transform 1 0 708 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_8353
timestamp 1745462530
transform 1 0 652 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_8354
timestamp 1745462530
transform 1 0 652 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_8355
timestamp 1745462530
transform 1 0 620 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_8356
timestamp 1745462530
transform 1 0 596 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_8357
timestamp 1745462530
transform 1 0 596 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_8358
timestamp 1745462530
transform 1 0 564 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_8359
timestamp 1745462530
transform 1 0 500 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_8360
timestamp 1745462530
transform 1 0 508 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_8361
timestamp 1745462530
transform 1 0 452 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_8362
timestamp 1745462530
transform 1 0 388 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_8363
timestamp 1745462530
transform 1 0 388 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_8364
timestamp 1745462530
transform 1 0 324 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_8365
timestamp 1745462530
transform 1 0 324 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_8366
timestamp 1745462530
transform 1 0 284 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_8367
timestamp 1745462530
transform 1 0 212 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_8368
timestamp 1745462530
transform 1 0 460 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_8369
timestamp 1745462530
transform 1 0 396 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_8370
timestamp 1745462530
transform 1 0 388 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_8371
timestamp 1745462530
transform 1 0 388 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8372
timestamp 1745462530
transform 1 0 260 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_8373
timestamp 1745462530
transform 1 0 220 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_8374
timestamp 1745462530
transform 1 0 220 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8375
timestamp 1745462530
transform 1 0 212 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_8376
timestamp 1745462530
transform 1 0 444 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8377
timestamp 1745462530
transform 1 0 412 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_8378
timestamp 1745462530
transform 1 0 340 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_8379
timestamp 1745462530
transform 1 0 268 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8380
timestamp 1745462530
transform 1 0 268 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_8381
timestamp 1745462530
transform 1 0 252 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_8382
timestamp 1745462530
transform 1 0 220 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_8383
timestamp 1745462530
transform 1 0 212 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_8384
timestamp 1745462530
transform 1 0 500 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_8385
timestamp 1745462530
transform 1 0 484 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_8386
timestamp 1745462530
transform 1 0 444 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_8387
timestamp 1745462530
transform 1 0 420 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_8388
timestamp 1745462530
transform 1 0 340 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_8389
timestamp 1745462530
transform 1 0 260 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_8390
timestamp 1745462530
transform 1 0 228 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_8391
timestamp 1745462530
transform 1 0 220 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8392
timestamp 1745462530
transform 1 0 724 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_8393
timestamp 1745462530
transform 1 0 724 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_8394
timestamp 1745462530
transform 1 0 700 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_8395
timestamp 1745462530
transform 1 0 692 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_8396
timestamp 1745462530
transform 1 0 652 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_8397
timestamp 1745462530
transform 1 0 644 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_8398
timestamp 1745462530
transform 1 0 556 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_8399
timestamp 1745462530
transform 1 0 556 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_8400
timestamp 1745462530
transform 1 0 948 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_8401
timestamp 1745462530
transform 1 0 908 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_8402
timestamp 1745462530
transform 1 0 892 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_8403
timestamp 1745462530
transform 1 0 876 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_8404
timestamp 1745462530
transform 1 0 860 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_8405
timestamp 1745462530
transform 1 0 836 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_8406
timestamp 1745462530
transform 1 0 820 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_8407
timestamp 1745462530
transform 1 0 812 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_8408
timestamp 1745462530
transform 1 0 1004 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_8409
timestamp 1745462530
transform 1 0 460 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_8410
timestamp 1745462530
transform 1 0 380 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_8411
timestamp 1745462530
transform 1 0 372 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_8412
timestamp 1745462530
transform 1 0 268 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_8413
timestamp 1745462530
transform 1 0 252 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_8414
timestamp 1745462530
transform 1 0 220 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_8415
timestamp 1745462530
transform 1 0 204 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_8416
timestamp 1745462530
transform 1 0 204 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_8417
timestamp 1745462530
transform 1 0 172 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_8418
timestamp 1745462530
transform 1 0 1076 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_8419
timestamp 1745462530
transform 1 0 940 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_8420
timestamp 1745462530
transform 1 0 836 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_8421
timestamp 1745462530
transform 1 0 820 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_8422
timestamp 1745462530
transform 1 0 804 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_8423
timestamp 1745462530
transform 1 0 740 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_8424
timestamp 1745462530
transform 1 0 676 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_8425
timestamp 1745462530
transform 1 0 676 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_8426
timestamp 1745462530
transform 1 0 1668 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_8427
timestamp 1745462530
transform 1 0 1588 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_8428
timestamp 1745462530
transform 1 0 1492 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_8429
timestamp 1745462530
transform 1 0 1484 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_8430
timestamp 1745462530
transform 1 0 1460 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_8431
timestamp 1745462530
transform 1 0 1148 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_8432
timestamp 1745462530
transform 1 0 1140 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_8433
timestamp 1745462530
transform 1 0 1108 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_8434
timestamp 1745462530
transform 1 0 1100 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_8435
timestamp 1745462530
transform 1 0 1940 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_8436
timestamp 1745462530
transform 1 0 1852 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_8437
timestamp 1745462530
transform 1 0 1692 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_8438
timestamp 1745462530
transform 1 0 1452 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_8439
timestamp 1745462530
transform 1 0 1444 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_8440
timestamp 1745462530
transform 1 0 1260 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_8441
timestamp 1745462530
transform 1 0 1172 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_8442
timestamp 1745462530
transform 1 0 1044 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_8443
timestamp 1745462530
transform 1 0 1908 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_8444
timestamp 1745462530
transform 1 0 1812 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_8445
timestamp 1745462530
transform 1 0 1676 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_8446
timestamp 1745462530
transform 1 0 1532 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_8447
timestamp 1745462530
transform 1 0 1468 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_8448
timestamp 1745462530
transform 1 0 1380 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_8449
timestamp 1745462530
transform 1 0 1340 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_8450
timestamp 1745462530
transform 1 0 1324 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_8451
timestamp 1745462530
transform 1 0 1916 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8452
timestamp 1745462530
transform 1 0 1908 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_8453
timestamp 1745462530
transform 1 0 1844 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_8454
timestamp 1745462530
transform 1 0 1748 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_8455
timestamp 1745462530
transform 1 0 1596 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8456
timestamp 1745462530
transform 1 0 1436 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_8457
timestamp 1745462530
transform 1 0 1364 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_8458
timestamp 1745462530
transform 1 0 1276 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_8459
timestamp 1745462530
transform 1 0 2036 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_8460
timestamp 1745462530
transform 1 0 1916 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_8461
timestamp 1745462530
transform 1 0 1916 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_8462
timestamp 1745462530
transform 1 0 1740 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_8463
timestamp 1745462530
transform 1 0 1524 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_8464
timestamp 1745462530
transform 1 0 1508 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_8465
timestamp 1745462530
transform 1 0 1436 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_8466
timestamp 1745462530
transform 1 0 1332 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_8467
timestamp 1745462530
transform 1 0 2020 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_8468
timestamp 1745462530
transform 1 0 1988 0 1 955
box -2 -2 2 2
use M2_M1  M2_M1_8469
timestamp 1745462530
transform 1 0 1940 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_8470
timestamp 1745462530
transform 1 0 1780 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_8471
timestamp 1745462530
transform 1 0 1588 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_8472
timestamp 1745462530
transform 1 0 1500 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_8473
timestamp 1745462530
transform 1 0 1396 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_8474
timestamp 1745462530
transform 1 0 1396 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_8475
timestamp 1745462530
transform 1 0 1980 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_8476
timestamp 1745462530
transform 1 0 1972 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_8477
timestamp 1745462530
transform 1 0 1820 0 1 1185
box -2 -2 2 2
use M2_M1  M2_M1_8478
timestamp 1745462530
transform 1 0 1620 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_8479
timestamp 1745462530
transform 1 0 1580 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_8480
timestamp 1745462530
transform 1 0 1556 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_8481
timestamp 1745462530
transform 1 0 1500 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_8482
timestamp 1745462530
transform 1 0 1428 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_8483
timestamp 1745462530
transform 1 0 1404 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_8484
timestamp 1745462530
transform 1 0 2020 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_8485
timestamp 1745462530
transform 1 0 1956 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_8486
timestamp 1745462530
transform 1 0 1908 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_8487
timestamp 1745462530
transform 1 0 1828 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_8488
timestamp 1745462530
transform 1 0 1620 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_8489
timestamp 1745462530
transform 1 0 1604 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_8490
timestamp 1745462530
transform 1 0 1556 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_8491
timestamp 1745462530
transform 1 0 1508 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_8492
timestamp 1745462530
transform 1 0 2884 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_8493
timestamp 1745462530
transform 1 0 2812 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_8494
timestamp 1745462530
transform 1 0 2708 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_8495
timestamp 1745462530
transform 1 0 2564 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_8496
timestamp 1745462530
transform 1 0 2340 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_8497
timestamp 1745462530
transform 1 0 2324 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_8498
timestamp 1745462530
transform 1 0 2268 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_8499
timestamp 1745462530
transform 1 0 2228 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_8500
timestamp 1745462530
transform 1 0 3092 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_8501
timestamp 1745462530
transform 1 0 3060 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_8502
timestamp 1745462530
transform 1 0 3044 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_8503
timestamp 1745462530
transform 1 0 3044 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8504
timestamp 1745462530
transform 1 0 2764 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_8505
timestamp 1745462530
transform 1 0 2700 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8506
timestamp 1745462530
transform 1 0 2628 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8507
timestamp 1745462530
transform 1 0 2300 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_8508
timestamp 1745462530
transform 1 0 2212 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_8509
timestamp 1745462530
transform 1 0 2212 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8510
timestamp 1745462530
transform 1 0 2828 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_8511
timestamp 1745462530
transform 1 0 2684 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_8512
timestamp 1745462530
transform 1 0 2676 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_8513
timestamp 1745462530
transform 1 0 2628 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_8514
timestamp 1745462530
transform 1 0 2604 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_8515
timestamp 1745462530
transform 1 0 2532 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_8516
timestamp 1745462530
transform 1 0 2316 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_8517
timestamp 1745462530
transform 1 0 2244 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_8518
timestamp 1745462530
transform 1 0 3020 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_8519
timestamp 1745462530
transform 1 0 2948 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_8520
timestamp 1745462530
transform 1 0 2788 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_8521
timestamp 1745462530
transform 1 0 2692 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_8522
timestamp 1745462530
transform 1 0 2644 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_8523
timestamp 1745462530
transform 1 0 2316 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_8524
timestamp 1745462530
transform 1 0 2308 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_8525
timestamp 1745462530
transform 1 0 2252 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_8526
timestamp 1745462530
transform 1 0 3124 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_8527
timestamp 1745462530
transform 1 0 3052 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_8528
timestamp 1745462530
transform 1 0 2980 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_8529
timestamp 1745462530
transform 1 0 2676 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_8530
timestamp 1745462530
transform 1 0 2660 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_8531
timestamp 1745462530
transform 1 0 2620 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_8532
timestamp 1745462530
transform 1 0 2516 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_8533
timestamp 1745462530
transform 1 0 2468 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_8534
timestamp 1745462530
transform 1 0 2876 0 1 985
box -2 -2 2 2
use M2_M1  M2_M1_8535
timestamp 1745462530
transform 1 0 2876 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_8536
timestamp 1745462530
transform 1 0 2764 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_8537
timestamp 1745462530
transform 1 0 2716 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_8538
timestamp 1745462530
transform 1 0 2548 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_8539
timestamp 1745462530
transform 1 0 2316 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_8540
timestamp 1745462530
transform 1 0 2276 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_8541
timestamp 1745462530
transform 1 0 2836 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_8542
timestamp 1745462530
transform 1 0 2828 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_8543
timestamp 1745462530
transform 1 0 2820 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_8544
timestamp 1745462530
transform 1 0 2820 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_8545
timestamp 1745462530
transform 1 0 2668 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_8546
timestamp 1745462530
transform 1 0 2636 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_8547
timestamp 1745462530
transform 1 0 2596 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_8548
timestamp 1745462530
transform 1 0 2348 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_8549
timestamp 1745462530
transform 1 0 2292 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_8550
timestamp 1745462530
transform 1 0 2796 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_8551
timestamp 1745462530
transform 1 0 2772 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_8552
timestamp 1745462530
transform 1 0 2684 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_8553
timestamp 1745462530
transform 1 0 2604 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_8554
timestamp 1745462530
transform 1 0 2580 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_8555
timestamp 1745462530
transform 1 0 2372 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_8556
timestamp 1745462530
transform 1 0 2364 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_8557
timestamp 1745462530
transform 1 0 3396 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_8558
timestamp 1745462530
transform 1 0 3364 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_8559
timestamp 1745462530
transform 1 0 3356 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_8560
timestamp 1745462530
transform 1 0 3300 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_8561
timestamp 1745462530
transform 1 0 3300 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_8562
timestamp 1745462530
transform 1 0 3244 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_8563
timestamp 1745462530
transform 1 0 3180 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_8564
timestamp 1745462530
transform 1 0 3180 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_8565
timestamp 1745462530
transform 1 0 3900 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_8566
timestamp 1745462530
transform 1 0 3828 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_8567
timestamp 1745462530
transform 1 0 3804 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_8568
timestamp 1745462530
transform 1 0 3756 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_8569
timestamp 1745462530
transform 1 0 3556 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_8570
timestamp 1745462530
transform 1 0 3540 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_8571
timestamp 1745462530
transform 1 0 3540 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_8572
timestamp 1745462530
transform 1 0 3372 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_8573
timestamp 1745462530
transform 1 0 4236 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_8574
timestamp 1745462530
transform 1 0 4236 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_8575
timestamp 1745462530
transform 1 0 4164 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_8576
timestamp 1745462530
transform 1 0 4092 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_8577
timestamp 1745462530
transform 1 0 4076 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_8578
timestamp 1745462530
transform 1 0 4028 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_8579
timestamp 1745462530
transform 1 0 3764 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_8580
timestamp 1745462530
transform 1 0 3620 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_8581
timestamp 1745462530
transform 1 0 4004 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_8582
timestamp 1745462530
transform 1 0 4004 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_8583
timestamp 1745462530
transform 1 0 3796 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8584
timestamp 1745462530
transform 1 0 3708 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_8585
timestamp 1745462530
transform 1 0 3660 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_8586
timestamp 1745462530
transform 1 0 3572 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_8587
timestamp 1745462530
transform 1 0 3532 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8588
timestamp 1745462530
transform 1 0 3388 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8589
timestamp 1745462530
transform 1 0 4340 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8590
timestamp 1745462530
transform 1 0 4324 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_8591
timestamp 1745462530
transform 1 0 4268 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_8592
timestamp 1745462530
transform 1 0 4236 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_8593
timestamp 1745462530
transform 1 0 4172 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_8594
timestamp 1745462530
transform 1 0 4164 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8595
timestamp 1745462530
transform 1 0 4108 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8596
timestamp 1745462530
transform 1 0 3820 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_8597
timestamp 1745462530
transform 1 0 4276 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_8598
timestamp 1745462530
transform 1 0 4220 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_8599
timestamp 1745462530
transform 1 0 4212 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_8600
timestamp 1745462530
transform 1 0 4196 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_8601
timestamp 1745462530
transform 1 0 4124 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_8602
timestamp 1745462530
transform 1 0 4044 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_8603
timestamp 1745462530
transform 1 0 3932 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_8604
timestamp 1745462530
transform 1 0 3292 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_8605
timestamp 1745462530
transform 1 0 4188 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_8606
timestamp 1745462530
transform 1 0 4148 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_8607
timestamp 1745462530
transform 1 0 4124 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_8608
timestamp 1745462530
transform 1 0 4084 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_8609
timestamp 1745462530
transform 1 0 3780 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_8610
timestamp 1745462530
transform 1 0 3428 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_8611
timestamp 1745462530
transform 1 0 3404 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_8612
timestamp 1745462530
transform 1 0 3380 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_8613
timestamp 1745462530
transform 1 0 3916 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_8614
timestamp 1745462530
transform 1 0 3860 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_8615
timestamp 1745462530
transform 1 0 3812 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_8616
timestamp 1745462530
transform 1 0 3772 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_8617
timestamp 1745462530
transform 1 0 3604 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_8618
timestamp 1745462530
transform 1 0 3460 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_8619
timestamp 1745462530
transform 1 0 3444 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_8620
timestamp 1745462530
transform 1 0 3364 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_8621
timestamp 1745462530
transform 1 0 4204 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_8622
timestamp 1745462530
transform 1 0 4204 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_8623
timestamp 1745462530
transform 1 0 4140 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_8624
timestamp 1745462530
transform 1 0 4116 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_8625
timestamp 1745462530
transform 1 0 4092 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_8626
timestamp 1745462530
transform 1 0 4084 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_8627
timestamp 1745462530
transform 1 0 4076 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_8628
timestamp 1745462530
transform 1 0 3492 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_8629
timestamp 1745462530
transform 1 0 3844 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_8630
timestamp 1745462530
transform 1 0 3820 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_8631
timestamp 1745462530
transform 1 0 3812 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_8632
timestamp 1745462530
transform 1 0 3700 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_8633
timestamp 1745462530
transform 1 0 3692 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_8634
timestamp 1745462530
transform 1 0 3692 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_8635
timestamp 1745462530
transform 1 0 3524 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_8636
timestamp 1745462530
transform 1 0 3492 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_8637
timestamp 1745462530
transform 1 0 4236 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_8638
timestamp 1745462530
transform 1 0 4236 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_8639
timestamp 1745462530
transform 1 0 4228 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_8640
timestamp 1745462530
transform 1 0 4196 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_8641
timestamp 1745462530
transform 1 0 4188 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_8642
timestamp 1745462530
transform 1 0 4132 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_8643
timestamp 1745462530
transform 1 0 4084 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_8644
timestamp 1745462530
transform 1 0 4028 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_8645
timestamp 1745462530
transform 1 0 3868 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_8646
timestamp 1745462530
transform 1 0 3852 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_8647
timestamp 1745462530
transform 1 0 3836 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_8648
timestamp 1745462530
transform 1 0 3828 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_8649
timestamp 1745462530
transform 1 0 3796 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_8650
timestamp 1745462530
transform 1 0 3700 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_8651
timestamp 1745462530
transform 1 0 3668 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_8652
timestamp 1745462530
transform 1 0 3588 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_8653
timestamp 1745462530
transform 1 0 4332 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_8654
timestamp 1745462530
transform 1 0 4308 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_8655
timestamp 1745462530
transform 1 0 4236 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_8656
timestamp 1745462530
transform 1 0 4180 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_8657
timestamp 1745462530
transform 1 0 4164 0 1 1795
box -2 -2 2 2
use M2_M1  M2_M1_8658
timestamp 1745462530
transform 1 0 4156 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_8659
timestamp 1745462530
transform 1 0 4004 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_8660
timestamp 1745462530
transform 1 0 3988 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_8661
timestamp 1745462530
transform 1 0 3860 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_8662
timestamp 1745462530
transform 1 0 3844 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_8663
timestamp 1745462530
transform 1 0 3732 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_8664
timestamp 1745462530
transform 1 0 3564 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_8665
timestamp 1745462530
transform 1 0 3340 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_8666
timestamp 1745462530
transform 1 0 3276 0 1 1895
box -2 -2 2 2
use M2_M1  M2_M1_8667
timestamp 1745462530
transform 1 0 3276 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_8668
timestamp 1745462530
transform 1 0 3268 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_8669
timestamp 1745462530
transform 1 0 3268 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_8670
timestamp 1745462530
transform 1 0 3196 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_8671
timestamp 1745462530
transform 1 0 3100 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_8672
timestamp 1745462530
transform 1 0 3100 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_8673
timestamp 1745462530
transform 1 0 2980 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_8674
timestamp 1745462530
transform 1 0 2956 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_8675
timestamp 1745462530
transform 1 0 2836 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_8676
timestamp 1745462530
transform 1 0 2828 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_8677
timestamp 1745462530
transform 1 0 2780 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_8678
timestamp 1745462530
transform 1 0 2764 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_8679
timestamp 1745462530
transform 1 0 2956 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_8680
timestamp 1745462530
transform 1 0 2924 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_8681
timestamp 1745462530
transform 1 0 2732 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_8682
timestamp 1745462530
transform 1 0 2700 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_8683
timestamp 1745462530
transform 1 0 2668 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_8684
timestamp 1745462530
transform 1 0 2660 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_8685
timestamp 1745462530
transform 1 0 2612 0 1 2185
box -2 -2 2 2
use M2_M1  M2_M1_8686
timestamp 1745462530
transform 1 0 2612 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_8687
timestamp 1745462530
transform 1 0 4188 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_8688
timestamp 1745462530
transform 1 0 4180 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_8689
timestamp 1745462530
transform 1 0 3844 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_8690
timestamp 1745462530
transform 1 0 3740 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_8691
timestamp 1745462530
transform 1 0 3652 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_8692
timestamp 1745462530
transform 1 0 3420 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_8693
timestamp 1745462530
transform 1 0 3268 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_8694
timestamp 1745462530
transform 1 0 3076 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_8695
timestamp 1745462530
transform 1 0 3908 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_8696
timestamp 1745462530
transform 1 0 3892 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_8697
timestamp 1745462530
transform 1 0 3892 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_8698
timestamp 1745462530
transform 1 0 3756 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_8699
timestamp 1745462530
transform 1 0 3692 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_8700
timestamp 1745462530
transform 1 0 3212 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_8701
timestamp 1745462530
transform 1 0 3100 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_8702
timestamp 1745462530
transform 1 0 2996 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_8703
timestamp 1745462530
transform 1 0 4140 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_8704
timestamp 1745462530
transform 1 0 4060 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_8705
timestamp 1745462530
transform 1 0 3996 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_8706
timestamp 1745462530
transform 1 0 3852 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_8707
timestamp 1745462530
transform 1 0 3620 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_8708
timestamp 1745462530
transform 1 0 3388 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_8709
timestamp 1745462530
transform 1 0 3244 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_8710
timestamp 1745462530
transform 1 0 3148 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_8711
timestamp 1745462530
transform 1 0 4220 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_8712
timestamp 1745462530
transform 1 0 4204 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_8713
timestamp 1745462530
transform 1 0 4148 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_8714
timestamp 1745462530
transform 1 0 3724 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_8715
timestamp 1745462530
transform 1 0 3524 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_8716
timestamp 1745462530
transform 1 0 3284 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_8717
timestamp 1745462530
transform 1 0 3196 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_8718
timestamp 1745462530
transform 1 0 2980 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_8719
timestamp 1745462530
transform 1 0 4204 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_8720
timestamp 1745462530
transform 1 0 4204 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_8721
timestamp 1745462530
transform 1 0 3932 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_8722
timestamp 1745462530
transform 1 0 3828 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_8723
timestamp 1745462530
transform 1 0 3628 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_8724
timestamp 1745462530
transform 1 0 3452 0 1 2404
box -2 -2 2 2
use M2_M1  M2_M1_8725
timestamp 1745462530
transform 1 0 3276 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_8726
timestamp 1745462530
transform 1 0 3052 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_8727
timestamp 1745462530
transform 1 0 4244 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_8728
timestamp 1745462530
transform 1 0 4196 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_8729
timestamp 1745462530
transform 1 0 4156 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_8730
timestamp 1745462530
transform 1 0 3948 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_8731
timestamp 1745462530
transform 1 0 3892 0 1 2305
box -2 -2 2 2
use M2_M1  M2_M1_8732
timestamp 1745462530
transform 1 0 3636 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_8733
timestamp 1745462530
transform 1 0 3388 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_8734
timestamp 1745462530
transform 1 0 3260 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_8735
timestamp 1745462530
transform 1 0 4116 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_8736
timestamp 1745462530
transform 1 0 4076 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_8737
timestamp 1745462530
transform 1 0 3860 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_8738
timestamp 1745462530
transform 1 0 3860 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_8739
timestamp 1745462530
transform 1 0 3700 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_8740
timestamp 1745462530
transform 1 0 3484 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_8741
timestamp 1745462530
transform 1 0 3212 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_8742
timestamp 1745462530
transform 1 0 3196 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_8743
timestamp 1745462530
transform 1 0 3020 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_8744
timestamp 1745462530
transform 1 0 2932 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_8745
timestamp 1745462530
transform 1 0 2852 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_8746
timestamp 1745462530
transform 1 0 2852 0 1 2545
box -2 -2 2 2
use M2_M1  M2_M1_8747
timestamp 1745462530
transform 1 0 2836 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_8748
timestamp 1745462530
transform 1 0 2836 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_8749
timestamp 1745462530
transform 1 0 2804 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_8750
timestamp 1745462530
transform 1 0 2748 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_8751
timestamp 1745462530
transform 1 0 2740 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_8752
timestamp 1745462530
transform 1 0 2828 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_8753
timestamp 1745462530
transform 1 0 2788 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_8754
timestamp 1745462530
transform 1 0 2764 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_8755
timestamp 1745462530
transform 1 0 2676 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_8756
timestamp 1745462530
transform 1 0 2612 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_8757
timestamp 1745462530
transform 1 0 2604 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_8758
timestamp 1745462530
transform 1 0 2484 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_8759
timestamp 1745462530
transform 1 0 2420 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_8760
timestamp 1745462530
transform 1 0 1788 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_8761
timestamp 1745462530
transform 1 0 1780 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_8762
timestamp 1745462530
transform 1 0 1756 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_8763
timestamp 1745462530
transform 1 0 1628 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_8764
timestamp 1745462530
transform 1 0 1788 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_8765
timestamp 1745462530
transform 1 0 1764 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_8766
timestamp 1745462530
transform 1 0 3788 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_8767
timestamp 1745462530
transform 1 0 1796 0 1 2235
box -2 -2 2 2
use M2_M1  M2_M1_8768
timestamp 1745462530
transform 1 0 3908 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_8769
timestamp 1745462530
transform 1 0 3764 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_8770
timestamp 1745462530
transform 1 0 3772 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_8771
timestamp 1745462530
transform 1 0 3740 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_8772
timestamp 1745462530
transform 1 0 3500 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_8773
timestamp 1745462530
transform 1 0 3476 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_8774
timestamp 1745462530
transform 1 0 3716 0 1 995
box -2 -2 2 2
use M2_M1  M2_M1_8775
timestamp 1745462530
transform 1 0 3004 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_8776
timestamp 1745462530
transform 1 0 3892 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_8777
timestamp 1745462530
transform 1 0 3748 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_8778
timestamp 1745462530
transform 1 0 3836 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_8779
timestamp 1745462530
transform 1 0 3828 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_8780
timestamp 1745462530
transform 1 0 3932 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_8781
timestamp 1745462530
transform 1 0 3868 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_8782
timestamp 1745462530
transform 1 0 3884 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_8783
timestamp 1745462530
transform 1 0 3852 0 1 1035
box -2 -2 2 2
use M2_M1  M2_M1_8784
timestamp 1745462530
transform 1 0 3852 0 1 345
box -2 -2 2 2
use M2_M1  M2_M1_8785
timestamp 1745462530
transform 1 0 3772 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_8786
timestamp 1745462530
transform 1 0 3924 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_8787
timestamp 1745462530
transform 1 0 3908 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_8788
timestamp 1745462530
transform 1 0 3892 0 1 395
box -2 -2 2 2
use M2_M1  M2_M1_8789
timestamp 1745462530
transform 1 0 3892 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_8790
timestamp 1745462530
transform 1 0 3780 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_8791
timestamp 1745462530
transform 1 0 3692 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8792
timestamp 1745462530
transform 1 0 3636 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_8793
timestamp 1745462530
transform 1 0 3564 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8794
timestamp 1745462530
transform 1 0 3340 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8795
timestamp 1745462530
transform 1 0 3340 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_8796
timestamp 1745462530
transform 1 0 3964 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_8797
timestamp 1745462530
transform 1 0 3948 0 1 385
box -2 -2 2 2
use M2_M1  M2_M1_8798
timestamp 1745462530
transform 1 0 3940 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_8799
timestamp 1745462530
transform 1 0 3740 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8800
timestamp 1745462530
transform 1 0 3700 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_8801
timestamp 1745462530
transform 1 0 3596 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8802
timestamp 1745462530
transform 1 0 3548 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_8803
timestamp 1745462530
transform 1 0 3396 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_8804
timestamp 1745462530
transform 1 0 3300 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8805
timestamp 1745462530
transform 1 0 3772 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_8806
timestamp 1745462530
transform 1 0 3724 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_8807
timestamp 1745462530
transform 1 0 3580 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_8808
timestamp 1745462530
transform 1 0 3580 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_8809
timestamp 1745462530
transform 1 0 3556 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_8810
timestamp 1745462530
transform 1 0 3556 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_8811
timestamp 1745462530
transform 1 0 3436 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_8812
timestamp 1745462530
transform 1 0 3236 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_8813
timestamp 1745462530
transform 1 0 3228 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8814
timestamp 1745462530
transform 1 0 3852 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_8815
timestamp 1745462530
transform 1 0 3788 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_8816
timestamp 1745462530
transform 1 0 3636 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_8817
timestamp 1745462530
transform 1 0 3596 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_8818
timestamp 1745462530
transform 1 0 3476 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_8819
timestamp 1745462530
transform 1 0 3300 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_8820
timestamp 1745462530
transform 1 0 3268 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8821
timestamp 1745462530
transform 1 0 3908 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_8822
timestamp 1745462530
transform 1 0 3908 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_8823
timestamp 1745462530
transform 1 0 3860 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_8824
timestamp 1745462530
transform 1 0 3620 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_8825
timestamp 1745462530
transform 1 0 3484 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_8826
timestamp 1745462530
transform 1 0 3332 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_8827
timestamp 1745462530
transform 1 0 3244 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_8828
timestamp 1745462530
transform 1 0 3244 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_8829
timestamp 1745462530
transform 1 0 3940 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_8830
timestamp 1745462530
transform 1 0 3940 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_8831
timestamp 1745462530
transform 1 0 3884 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_8832
timestamp 1745462530
transform 1 0 3652 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_8833
timestamp 1745462530
transform 1 0 3508 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_8834
timestamp 1745462530
transform 1 0 3380 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_8835
timestamp 1745462530
transform 1 0 3364 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_8836
timestamp 1745462530
transform 1 0 3236 0 1 1115
box -2 -2 2 2
use M2_M1  M2_M1_8837
timestamp 1745462530
transform 1 0 3876 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_8838
timestamp 1745462530
transform 1 0 3820 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_8839
timestamp 1745462530
transform 1 0 3636 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_8840
timestamp 1745462530
transform 1 0 3612 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_8841
timestamp 1745462530
transform 1 0 3540 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_8842
timestamp 1745462530
transform 1 0 3428 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_8843
timestamp 1745462530
transform 1 0 3308 0 1 1035
box -2 -2 2 2
use M2_M1  M2_M1_8844
timestamp 1745462530
transform 1 0 3196 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_8845
timestamp 1745462530
transform 1 0 3892 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_8846
timestamp 1745462530
transform 1 0 3852 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_8847
timestamp 1745462530
transform 1 0 3836 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_8848
timestamp 1745462530
transform 1 0 3692 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_8849
timestamp 1745462530
transform 1 0 3628 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_8850
timestamp 1745462530
transform 1 0 3572 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_8851
timestamp 1745462530
transform 1 0 3412 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_8852
timestamp 1745462530
transform 1 0 3356 0 1 1035
box -2 -2 2 2
use M2_M1  M2_M1_8853
timestamp 1745462530
transform 1 0 3212 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_8854
timestamp 1745462530
transform 1 0 2972 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_8855
timestamp 1745462530
transform 1 0 2940 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_8856
timestamp 1745462530
transform 1 0 3076 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_8857
timestamp 1745462530
transform 1 0 2988 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_8858
timestamp 1745462530
transform 1 0 2996 0 1 1035
box -2 -2 2 2
use M2_M1  M2_M1_8859
timestamp 1745462530
transform 1 0 2956 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8860
timestamp 1745462530
transform 1 0 2908 0 1 595
box -2 -2 2 2
use M2_M1  M2_M1_8861
timestamp 1745462530
transform 1 0 2884 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8862
timestamp 1745462530
transform 1 0 2948 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_8863
timestamp 1745462530
transform 1 0 2940 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8864
timestamp 1745462530
transform 1 0 2908 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_8865
timestamp 1745462530
transform 1 0 2804 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_8866
timestamp 1745462530
transform 1 0 2684 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_8867
timestamp 1745462530
transform 1 0 2644 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_8868
timestamp 1745462530
transform 1 0 2572 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8869
timestamp 1745462530
transform 1 0 2508 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_8870
timestamp 1745462530
transform 1 0 2452 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_8871
timestamp 1745462530
transform 1 0 2372 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_8872
timestamp 1745462530
transform 1 0 2964 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_8873
timestamp 1745462530
transform 1 0 2860 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_8874
timestamp 1745462530
transform 1 0 2724 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_8875
timestamp 1745462530
transform 1 0 2604 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8876
timestamp 1745462530
transform 1 0 2604 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_8877
timestamp 1745462530
transform 1 0 2540 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_8878
timestamp 1745462530
transform 1 0 2484 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_8879
timestamp 1745462530
transform 1 0 2420 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_8880
timestamp 1745462530
transform 1 0 2916 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8881
timestamp 1745462530
transform 1 0 2868 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8882
timestamp 1745462530
transform 1 0 2844 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8883
timestamp 1745462530
transform 1 0 2764 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8884
timestamp 1745462530
transform 1 0 2644 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_8885
timestamp 1745462530
transform 1 0 2572 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_8886
timestamp 1745462530
transform 1 0 2460 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8887
timestamp 1745462530
transform 1 0 2316 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8888
timestamp 1745462530
transform 1 0 2252 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8889
timestamp 1745462530
transform 1 0 2964 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8890
timestamp 1745462530
transform 1 0 2900 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8891
timestamp 1745462530
transform 1 0 2796 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8892
timestamp 1745462530
transform 1 0 2636 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_8893
timestamp 1745462530
transform 1 0 2604 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8894
timestamp 1745462530
transform 1 0 2492 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8895
timestamp 1745462530
transform 1 0 2348 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8896
timestamp 1745462530
transform 1 0 2308 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8897
timestamp 1745462530
transform 1 0 3044 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_8898
timestamp 1745462530
transform 1 0 3036 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_8899
timestamp 1745462530
transform 1 0 2844 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_8900
timestamp 1745462530
transform 1 0 2828 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_8901
timestamp 1745462530
transform 1 0 2676 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_8902
timestamp 1745462530
transform 1 0 2636 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_8903
timestamp 1745462530
transform 1 0 2508 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_8904
timestamp 1745462530
transform 1 0 2484 0 1 835
box -2 -2 2 2
use M2_M1  M2_M1_8905
timestamp 1745462530
transform 1 0 2476 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_8906
timestamp 1745462530
transform 1 0 3100 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_8907
timestamp 1745462530
transform 1 0 3068 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_8908
timestamp 1745462530
transform 1 0 2852 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_8909
timestamp 1745462530
transform 1 0 2788 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_8910
timestamp 1745462530
transform 1 0 2716 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_8911
timestamp 1745462530
transform 1 0 2652 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_8912
timestamp 1745462530
transform 1 0 2524 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_8913
timestamp 1745462530
transform 1 0 2524 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_8914
timestamp 1745462530
transform 1 0 2980 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_8915
timestamp 1745462530
transform 1 0 2916 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_8916
timestamp 1745462530
transform 1 0 2756 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_8917
timestamp 1745462530
transform 1 0 2724 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_8918
timestamp 1745462530
transform 1 0 2508 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_8919
timestamp 1745462530
transform 1 0 2508 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_8920
timestamp 1745462530
transform 1 0 2436 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_8921
timestamp 1745462530
transform 1 0 2436 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_8922
timestamp 1745462530
transform 1 0 3140 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_8923
timestamp 1745462530
transform 1 0 3012 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_8924
timestamp 1745462530
transform 1 0 2948 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_8925
timestamp 1745462530
transform 1 0 2820 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_8926
timestamp 1745462530
transform 1 0 2652 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_8927
timestamp 1745462530
transform 1 0 2548 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_8928
timestamp 1745462530
transform 1 0 2524 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_8929
timestamp 1745462530
transform 1 0 2492 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_8930
timestamp 1745462530
transform 1 0 3908 0 1 2195
box -2 -2 2 2
use M2_M1  M2_M1_8931
timestamp 1745462530
transform 1 0 3900 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_8932
timestamp 1745462530
transform 1 0 4012 0 1 2715
box -2 -2 2 2
use M2_M1  M2_M1_8933
timestamp 1745462530
transform 1 0 3940 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_8934
timestamp 1745462530
transform 1 0 4060 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_8935
timestamp 1745462530
transform 1 0 3988 0 1 2715
box -2 -2 2 2
use M2_M1  M2_M1_8936
timestamp 1745462530
transform 1 0 3972 0 1 2705
box -2 -2 2 2
use M2_M1  M2_M1_8937
timestamp 1745462530
transform 1 0 3948 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_8938
timestamp 1745462530
transform 1 0 4100 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_8939
timestamp 1745462530
transform 1 0 4004 0 1 2705
box -2 -2 2 2
use M2_M1  M2_M1_8940
timestamp 1745462530
transform 1 0 4084 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_8941
timestamp 1745462530
transform 1 0 4060 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_8942
timestamp 1745462530
transform 1 0 3836 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_8943
timestamp 1745462530
transform 1 0 3484 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_8944
timestamp 1745462530
transform 1 0 3308 0 1 2595
box -2 -2 2 2
use M2_M1  M2_M1_8945
timestamp 1745462530
transform 1 0 3172 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_8946
timestamp 1745462530
transform 1 0 2980 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_8947
timestamp 1745462530
transform 1 0 2900 0 1 2345
box -2 -2 2 2
use M2_M1  M2_M1_8948
timestamp 1745462530
transform 1 0 4172 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_8949
timestamp 1745462530
transform 1 0 4108 0 1 2595
box -2 -2 2 2
use M2_M1  M2_M1_8950
timestamp 1745462530
transform 1 0 4148 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_8951
timestamp 1745462530
transform 1 0 4140 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_8952
timestamp 1745462530
transform 1 0 3868 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_8953
timestamp 1745462530
transform 1 0 3804 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_8954
timestamp 1745462530
transform 1 0 3524 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_8955
timestamp 1745462530
transform 1 0 3356 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_8956
timestamp 1745462530
transform 1 0 3188 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_8957
timestamp 1745462530
transform 1 0 2572 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_8958
timestamp 1745462530
transform 1 0 4188 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_8959
timestamp 1745462530
transform 1 0 4172 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_8960
timestamp 1745462530
transform 1 0 3916 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_8961
timestamp 1745462530
transform 1 0 3860 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_8962
timestamp 1745462530
transform 1 0 3556 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_8963
timestamp 1745462530
transform 1 0 3404 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_8964
timestamp 1745462530
transform 1 0 3228 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_8965
timestamp 1745462530
transform 1 0 2668 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_8966
timestamp 1745462530
transform 1 0 3988 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_8967
timestamp 1745462530
transform 1 0 3900 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_8968
timestamp 1745462530
transform 1 0 3724 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_8969
timestamp 1745462530
transform 1 0 3556 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_8970
timestamp 1745462530
transform 1 0 3380 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_8971
timestamp 1745462530
transform 1 0 3100 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_8972
timestamp 1745462530
transform 1 0 3068 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_8973
timestamp 1745462530
transform 1 0 2708 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_8974
timestamp 1745462530
transform 1 0 4004 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_8975
timestamp 1745462530
transform 1 0 3956 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_8976
timestamp 1745462530
transform 1 0 3764 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_8977
timestamp 1745462530
transform 1 0 3612 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_8978
timestamp 1745462530
transform 1 0 3396 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_8979
timestamp 1745462530
transform 1 0 3116 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_8980
timestamp 1745462530
transform 1 0 3108 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_8981
timestamp 1745462530
transform 1 0 2708 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_8982
timestamp 1745462530
transform 1 0 4036 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_8983
timestamp 1745462530
transform 1 0 4036 0 1 2745
box -2 -2 2 2
use M2_M1  M2_M1_8984
timestamp 1745462530
transform 1 0 3780 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_8985
timestamp 1745462530
transform 1 0 3540 0 1 2795
box -2 -2 2 2
use M2_M1  M2_M1_8986
timestamp 1745462530
transform 1 0 3300 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_8987
timestamp 1745462530
transform 1 0 2988 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_8988
timestamp 1745462530
transform 1 0 2956 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_8989
timestamp 1745462530
transform 1 0 2628 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_8990
timestamp 1745462530
transform 1 0 4068 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_8991
timestamp 1745462530
transform 1 0 4052 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_8992
timestamp 1745462530
transform 1 0 3812 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_8993
timestamp 1745462530
transform 1 0 3572 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_8994
timestamp 1745462530
transform 1 0 3340 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_8995
timestamp 1745462530
transform 1 0 3028 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_8996
timestamp 1745462530
transform 1 0 3012 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_8997
timestamp 1745462530
transform 1 0 2676 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_8998
timestamp 1745462530
transform 1 0 3868 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_8999
timestamp 1745462530
transform 1 0 3004 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_9000
timestamp 1745462530
transform 1 0 3852 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_9001
timestamp 1745462530
transform 1 0 3836 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_9002
timestamp 1745462530
transform 1 0 3884 0 1 2105
box -2 -2 2 2
use M2_M1  M2_M1_9003
timestamp 1745462530
transform 1 0 3884 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_9004
timestamp 1745462530
transform 1 0 3892 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_9005
timestamp 1745462530
transform 1 0 3876 0 1 1945
box -2 -2 2 2
use M2_M1  M2_M1_9006
timestamp 1745462530
transform 1 0 3924 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_9007
timestamp 1745462530
transform 1 0 3892 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_9008
timestamp 1745462530
transform 1 0 3964 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_9009
timestamp 1745462530
transform 1 0 3908 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_9010
timestamp 1745462530
transform 1 0 3844 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_9011
timestamp 1745462530
transform 1 0 3732 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_9012
timestamp 1745462530
transform 1 0 3644 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_9013
timestamp 1745462530
transform 1 0 3588 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_9014
timestamp 1745462530
transform 1 0 3460 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_9015
timestamp 1745462530
transform 1 0 3404 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_9016
timestamp 1745462530
transform 1 0 3964 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_9017
timestamp 1745462530
transform 1 0 3940 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_9018
timestamp 1745462530
transform 1 0 3940 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_9019
timestamp 1745462530
transform 1 0 3940 0 1 1795
box -2 -2 2 2
use M2_M1  M2_M1_9020
timestamp 1745462530
transform 1 0 3900 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_9021
timestamp 1745462530
transform 1 0 3828 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_9022
timestamp 1745462530
transform 1 0 3772 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_9023
timestamp 1745462530
transform 1 0 3676 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_9024
timestamp 1745462530
transform 1 0 3668 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_9025
timestamp 1745462530
transform 1 0 3500 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_9026
timestamp 1745462530
transform 1 0 3340 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_9027
timestamp 1745462530
transform 1 0 3988 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_9028
timestamp 1745462530
transform 1 0 3876 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_9029
timestamp 1745462530
transform 1 0 3860 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_9030
timestamp 1745462530
transform 1 0 3748 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_9031
timestamp 1745462530
transform 1 0 3548 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_9032
timestamp 1745462530
transform 1 0 3516 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_9033
timestamp 1745462530
transform 1 0 3396 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_9034
timestamp 1745462530
transform 1 0 3364 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_9035
timestamp 1745462530
transform 1 0 3292 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_9036
timestamp 1745462530
transform 1 0 3932 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_9037
timestamp 1745462530
transform 1 0 3908 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_9038
timestamp 1745462530
transform 1 0 3788 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_9039
timestamp 1745462530
transform 1 0 3764 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_9040
timestamp 1745462530
transform 1 0 3604 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_9041
timestamp 1745462530
transform 1 0 3572 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_9042
timestamp 1745462530
transform 1 0 3452 0 1 1395
box -2 -2 2 2
use M2_M1  M2_M1_9043
timestamp 1745462530
transform 1 0 3268 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_9044
timestamp 1745462530
transform 1 0 3804 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_9045
timestamp 1745462530
transform 1 0 3804 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_9046
timestamp 1745462530
transform 1 0 3548 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_9047
timestamp 1745462530
transform 1 0 3444 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_9048
timestamp 1745462530
transform 1 0 3316 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_9049
timestamp 1745462530
transform 1 0 3260 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_9050
timestamp 1745462530
transform 1 0 3204 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_9051
timestamp 1745462530
transform 1 0 3204 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_9052
timestamp 1745462530
transform 1 0 3172 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_9053
timestamp 1745462530
transform 1 0 3844 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_9054
timestamp 1745462530
transform 1 0 3820 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_9055
timestamp 1745462530
transform 1 0 3564 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_9056
timestamp 1745462530
transform 1 0 3460 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_9057
timestamp 1745462530
transform 1 0 3388 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_9058
timestamp 1745462530
transform 1 0 3244 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_9059
timestamp 1745462530
transform 1 0 3180 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_9060
timestamp 1745462530
transform 1 0 3060 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_9061
timestamp 1745462530
transform 1 0 2980 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_9062
timestamp 1745462530
transform 1 0 2980 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_9063
timestamp 1745462530
transform 1 0 2956 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_9064
timestamp 1745462530
transform 1 0 2948 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_9065
timestamp 1745462530
transform 1 0 2940 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_9066
timestamp 1745462530
transform 1 0 2940 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_9067
timestamp 1745462530
transform 1 0 2924 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_9068
timestamp 1745462530
transform 1 0 2916 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_9069
timestamp 1745462530
transform 1 0 2916 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_9070
timestamp 1745462530
transform 1 0 2908 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_9071
timestamp 1745462530
transform 1 0 2884 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_9072
timestamp 1745462530
transform 1 0 2860 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_9073
timestamp 1745462530
transform 1 0 3020 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_9074
timestamp 1745462530
transform 1 0 3020 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_9075
timestamp 1745462530
transform 1 0 3012 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_9076
timestamp 1745462530
transform 1 0 3004 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_9077
timestamp 1745462530
transform 1 0 2956 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_9078
timestamp 1745462530
transform 1 0 2948 0 1 2395
box -2 -2 2 2
use M2_M1  M2_M1_9079
timestamp 1745462530
transform 1 0 2940 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_9080
timestamp 1745462530
transform 1 0 2876 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_9081
timestamp 1745462530
transform 1 0 1972 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_9082
timestamp 1745462530
transform 1 0 1748 0 1 2195
box -2 -2 2 2
use M2_M1  M2_M1_9083
timestamp 1745462530
transform 1 0 1772 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_9084
timestamp 1745462530
transform 1 0 684 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_9085
timestamp 1745462530
transform 1 0 732 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_9086
timestamp 1745462530
transform 1 0 660 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_9087
timestamp 1745462530
transform 1 0 668 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_9088
timestamp 1745462530
transform 1 0 620 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_9089
timestamp 1745462530
transform 1 0 676 0 1 2395
box -2 -2 2 2
use M2_M1  M2_M1_9090
timestamp 1745462530
transform 1 0 676 0 1 2235
box -2 -2 2 2
use M2_M1  M2_M1_9091
timestamp 1745462530
transform 1 0 692 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_9092
timestamp 1745462530
transform 1 0 652 0 1 2395
box -2 -2 2 2
use M2_M1  M2_M1_9093
timestamp 1745462530
transform 1 0 708 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_9094
timestamp 1745462530
transform 1 0 668 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_9095
timestamp 1745462530
transform 1 0 876 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_9096
timestamp 1745462530
transform 1 0 860 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_9097
timestamp 1745462530
transform 1 0 828 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_9098
timestamp 1745462530
transform 1 0 724 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_9099
timestamp 1745462530
transform 1 0 708 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_9100
timestamp 1745462530
transform 1 0 700 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_9101
timestamp 1745462530
transform 1 0 676 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_9102
timestamp 1745462530
transform 1 0 452 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_9103
timestamp 1745462530
transform 1 0 948 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_9104
timestamp 1745462530
transform 1 0 940 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_9105
timestamp 1745462530
transform 1 0 908 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_9106
timestamp 1745462530
transform 1 0 900 0 1 2795
box -2 -2 2 2
use M2_M1  M2_M1_9107
timestamp 1745462530
transform 1 0 764 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_9108
timestamp 1745462530
transform 1 0 756 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_9109
timestamp 1745462530
transform 1 0 740 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_9110
timestamp 1745462530
transform 1 0 732 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_9111
timestamp 1745462530
transform 1 0 868 0 1 2435
box -2 -2 2 2
use M2_M1  M2_M1_9112
timestamp 1745462530
transform 1 0 828 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_9113
timestamp 1745462530
transform 1 0 772 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_9114
timestamp 1745462530
transform 1 0 676 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_9115
timestamp 1745462530
transform 1 0 660 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_9116
timestamp 1745462530
transform 1 0 652 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_9117
timestamp 1745462530
transform 1 0 628 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_9118
timestamp 1745462530
transform 1 0 628 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_9119
timestamp 1745462530
transform 1 0 516 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_9120
timestamp 1745462530
transform 1 0 900 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_9121
timestamp 1745462530
transform 1 0 876 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_9122
timestamp 1745462530
transform 1 0 812 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_9123
timestamp 1745462530
transform 1 0 716 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_9124
timestamp 1745462530
transform 1 0 700 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_9125
timestamp 1745462530
transform 1 0 684 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_9126
timestamp 1745462530
transform 1 0 684 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_9127
timestamp 1745462530
transform 1 0 660 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_9128
timestamp 1745462530
transform 1 0 660 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_9129
timestamp 1745462530
transform 1 0 964 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_9130
timestamp 1745462530
transform 1 0 788 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_9131
timestamp 1745462530
transform 1 0 788 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_9132
timestamp 1745462530
transform 1 0 692 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_9133
timestamp 1745462530
transform 1 0 644 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_9134
timestamp 1745462530
transform 1 0 588 0 1 2185
box -2 -2 2 2
use M2_M1  M2_M1_9135
timestamp 1745462530
transform 1 0 588 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_9136
timestamp 1745462530
transform 1 0 532 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_9137
timestamp 1745462530
transform 1 0 1012 0 1 2235
box -2 -2 2 2
use M2_M1  M2_M1_9138
timestamp 1745462530
transform 1 0 836 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_9139
timestamp 1745462530
transform 1 0 804 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_9140
timestamp 1745462530
transform 1 0 740 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_9141
timestamp 1745462530
transform 1 0 660 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_9142
timestamp 1745462530
transform 1 0 644 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_9143
timestamp 1745462530
transform 1 0 620 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_9144
timestamp 1745462530
transform 1 0 604 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_9145
timestamp 1745462530
transform 1 0 940 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_9146
timestamp 1745462530
transform 1 0 908 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_9147
timestamp 1745462530
transform 1 0 804 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_9148
timestamp 1745462530
transform 1 0 788 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_9149
timestamp 1745462530
transform 1 0 748 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_9150
timestamp 1745462530
transform 1 0 740 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_9151
timestamp 1745462530
transform 1 0 684 0 1 1995
box -2 -2 2 2
use M2_M1  M2_M1_9152
timestamp 1745462530
transform 1 0 684 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_9153
timestamp 1745462530
transform 1 0 652 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_9154
timestamp 1745462530
transform 1 0 1100 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_9155
timestamp 1745462530
transform 1 0 932 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_9156
timestamp 1745462530
transform 1 0 860 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_9157
timestamp 1745462530
transform 1 0 804 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_9158
timestamp 1745462530
transform 1 0 796 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_9159
timestamp 1745462530
transform 1 0 740 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_9160
timestamp 1745462530
transform 1 0 668 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_9161
timestamp 1745462530
transform 1 0 476 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_9162
timestamp 1745462530
transform 1 0 1980 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_9163
timestamp 1745462530
transform 1 0 1948 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_9164
timestamp 1745462530
transform 1 0 1996 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_9165
timestamp 1745462530
transform 1 0 1956 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_9166
timestamp 1745462530
transform 1 0 1948 0 1 2305
box -2 -2 2 2
use M2_M1  M2_M1_9167
timestamp 1745462530
transform 1 0 1932 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_9168
timestamp 1745462530
transform 1 0 2012 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_9169
timestamp 1745462530
transform 1 0 1924 0 1 2345
box -2 -2 2 2
use M2_M1  M2_M1_9170
timestamp 1745462530
transform 1 0 1940 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_9171
timestamp 1745462530
transform 1 0 1724 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_9172
timestamp 1745462530
transform 1 0 1772 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_9173
timestamp 1745462530
transform 1 0 1708 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_9174
timestamp 1745462530
transform 1 0 1540 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_9175
timestamp 1745462530
transform 1 0 1324 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_9176
timestamp 1745462530
transform 1 0 1180 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_9177
timestamp 1745462530
transform 1 0 1124 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_9178
timestamp 1745462530
transform 1 0 1036 0 1 2505
box -2 -2 2 2
use M2_M1  M2_M1_9179
timestamp 1745462530
transform 1 0 1036 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_9180
timestamp 1745462530
transform 1 0 1020 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_9181
timestamp 1745462530
transform 1 0 996 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_9182
timestamp 1745462530
transform 1 0 2076 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_9183
timestamp 1745462530
transform 1 0 1812 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_9184
timestamp 1745462530
transform 1 0 1748 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_9185
timestamp 1745462530
transform 1 0 1596 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_9186
timestamp 1745462530
transform 1 0 1420 0 1 2235
box -2 -2 2 2
use M2_M1  M2_M1_9187
timestamp 1745462530
transform 1 0 1388 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_9188
timestamp 1745462530
transform 1 0 1236 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_9189
timestamp 1745462530
transform 1 0 1156 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_9190
timestamp 1745462530
transform 1 0 2108 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_9191
timestamp 1745462530
transform 1 0 1980 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_9192
timestamp 1745462530
transform 1 0 1844 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_9193
timestamp 1745462530
transform 1 0 1652 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_9194
timestamp 1745462530
transform 1 0 1444 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_9195
timestamp 1745462530
transform 1 0 1380 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_9196
timestamp 1745462530
transform 1 0 1252 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_9197
timestamp 1745462530
transform 1 0 1244 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_9198
timestamp 1745462530
transform 1 0 1212 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_9199
timestamp 1745462530
transform 1 0 2124 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_9200
timestamp 1745462530
transform 1 0 2028 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_9201
timestamp 1745462530
transform 1 0 1924 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_9202
timestamp 1745462530
transform 1 0 1692 0 1 2305
box -2 -2 2 2
use M2_M1  M2_M1_9203
timestamp 1745462530
transform 1 0 1476 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_9204
timestamp 1745462530
transform 1 0 1388 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_9205
timestamp 1745462530
transform 1 0 1308 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_9206
timestamp 1745462530
transform 1 0 1284 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_9207
timestamp 1745462530
transform 1 0 1284 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_9208
timestamp 1745462530
transform 1 0 2388 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_9209
timestamp 1745462530
transform 1 0 2220 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_9210
timestamp 1745462530
transform 1 0 1980 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_9211
timestamp 1745462530
transform 1 0 1908 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_9212
timestamp 1745462530
transform 1 0 1652 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_9213
timestamp 1745462530
transform 1 0 1500 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_9214
timestamp 1745462530
transform 1 0 1444 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_9215
timestamp 1745462530
transform 1 0 1428 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_9216
timestamp 1745462530
transform 1 0 2076 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_9217
timestamp 1745462530
transform 1 0 2004 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_9218
timestamp 1745462530
transform 1 0 1948 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_9219
timestamp 1745462530
transform 1 0 1692 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_9220
timestamp 1745462530
transform 1 0 1516 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_9221
timestamp 1745462530
transform 1 0 1460 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_9222
timestamp 1745462530
transform 1 0 1460 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_9223
timestamp 1745462530
transform 1 0 2140 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_9224
timestamp 1745462530
transform 1 0 1972 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_9225
timestamp 1745462530
transform 1 0 1908 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_9226
timestamp 1745462530
transform 1 0 1628 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_9227
timestamp 1745462530
transform 1 0 1516 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_9228
timestamp 1745462530
transform 1 0 1508 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_9229
timestamp 1745462530
transform 1 0 1340 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_9230
timestamp 1745462530
transform 1 0 1188 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_9231
timestamp 1745462530
transform 1 0 2156 0 1 2395
box -2 -2 2 2
use M2_M1  M2_M1_9232
timestamp 1745462530
transform 1 0 1988 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_9233
timestamp 1745462530
transform 1 0 1924 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_9234
timestamp 1745462530
transform 1 0 1684 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_9235
timestamp 1745462530
transform 1 0 1572 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_9236
timestamp 1745462530
transform 1 0 1452 0 1 2515
box -2 -2 2 2
use M2_M1  M2_M1_9237
timestamp 1745462530
transform 1 0 1372 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_9238
timestamp 1745462530
transform 1 0 1204 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_9239
timestamp 1745462530
transform 1 0 1620 0 1 995
box -2 -2 2 2
use M2_M1  M2_M1_9240
timestamp 1745462530
transform 1 0 708 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_9241
timestamp 1745462530
transform 1 0 1676 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_9242
timestamp 1745462530
transform 1 0 1636 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_9243
timestamp 1745462530
transform 1 0 1660 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_9244
timestamp 1745462530
transform 1 0 1660 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_9245
timestamp 1745462530
transform 1 0 1668 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_9246
timestamp 1745462530
transform 1 0 1660 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_9247
timestamp 1745462530
transform 1 0 1660 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_9248
timestamp 1745462530
transform 1 0 1652 0 1 1035
box -2 -2 2 2
use M2_M1  M2_M1_9249
timestamp 1745462530
transform 1 0 1644 0 1 745
box -2 -2 2 2
use M2_M1  M2_M1_9250
timestamp 1745462530
transform 1 0 1620 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_9251
timestamp 1745462530
transform 1 0 1700 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_9252
timestamp 1745462530
transform 1 0 1692 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_9253
timestamp 1745462530
transform 1 0 1980 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_9254
timestamp 1745462530
transform 1 0 1924 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_9255
timestamp 1745462530
transform 1 0 1788 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_9256
timestamp 1745462530
transform 1 0 1668 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_9257
timestamp 1745462530
transform 1 0 1500 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_9258
timestamp 1745462530
transform 1 0 1420 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_9259
timestamp 1745462530
transform 1 0 1308 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_9260
timestamp 1745462530
transform 1 0 1244 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_9261
timestamp 1745462530
transform 1 0 1972 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_9262
timestamp 1745462530
transform 1 0 1884 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_9263
timestamp 1745462530
transform 1 0 1828 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_9264
timestamp 1745462530
transform 1 0 1716 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_9265
timestamp 1745462530
transform 1 0 1580 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_9266
timestamp 1745462530
transform 1 0 1452 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_9267
timestamp 1745462530
transform 1 0 1348 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_9268
timestamp 1745462530
transform 1 0 1300 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_9269
timestamp 1745462530
transform 1 0 1908 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_9270
timestamp 1745462530
transform 1 0 1836 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_9271
timestamp 1745462530
transform 1 0 1588 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_9272
timestamp 1745462530
transform 1 0 1588 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_9273
timestamp 1745462530
transform 1 0 1348 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_9274
timestamp 1745462530
transform 1 0 1268 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_9275
timestamp 1745462530
transform 1 0 1164 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_9276
timestamp 1745462530
transform 1 0 1092 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_9277
timestamp 1745462530
transform 1 0 1956 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_9278
timestamp 1745462530
transform 1 0 1900 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_9279
timestamp 1745462530
transform 1 0 1636 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_9280
timestamp 1745462530
transform 1 0 1564 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_9281
timestamp 1745462530
transform 1 0 1380 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_9282
timestamp 1745462530
transform 1 0 1196 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_9283
timestamp 1745462530
transform 1 0 1132 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_9284
timestamp 1745462530
transform 1 0 1956 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_9285
timestamp 1745462530
transform 1 0 1892 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_9286
timestamp 1745462530
transform 1 0 1636 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_9287
timestamp 1745462530
transform 1 0 1612 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_9288
timestamp 1745462530
transform 1 0 1476 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_9289
timestamp 1745462530
transform 1 0 1460 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_9290
timestamp 1745462530
transform 1 0 1228 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_9291
timestamp 1745462530
transform 1 0 1228 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_9292
timestamp 1745462530
transform 1 0 1972 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_9293
timestamp 1745462530
transform 1 0 1916 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_9294
timestamp 1745462530
transform 1 0 1676 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_9295
timestamp 1745462530
transform 1 0 1492 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_9296
timestamp 1745462530
transform 1 0 1380 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_9297
timestamp 1745462530
transform 1 0 1244 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_9298
timestamp 1745462530
transform 1 0 1244 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_9299
timestamp 1745462530
transform 1 0 2068 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_9300
timestamp 1745462530
transform 1 0 1900 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_9301
timestamp 1745462530
transform 1 0 1876 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_9302
timestamp 1745462530
transform 1 0 1644 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_9303
timestamp 1745462530
transform 1 0 1508 0 1 1315
box -2 -2 2 2
use M2_M1  M2_M1_9304
timestamp 1745462530
transform 1 0 1452 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_9305
timestamp 1745462530
transform 1 0 1260 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_9306
timestamp 1745462530
transform 1 0 1260 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_9307
timestamp 1745462530
transform 1 0 2300 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_9308
timestamp 1745462530
transform 1 0 2300 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_9309
timestamp 1745462530
transform 1 0 2084 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_9310
timestamp 1745462530
transform 1 0 1916 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_9311
timestamp 1745462530
transform 1 0 1668 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_9312
timestamp 1745462530
transform 1 0 1508 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_9313
timestamp 1745462530
transform 1 0 1308 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_9314
timestamp 1745462530
transform 1 0 1300 0 1 1295
box -2 -2 2 2
use M2_M1  M2_M1_9315
timestamp 1745462530
transform 1 0 660 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_9316
timestamp 1745462530
transform 1 0 636 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_9317
timestamp 1745462530
transform 1 0 692 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_9318
timestamp 1745462530
transform 1 0 676 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_9319
timestamp 1745462530
transform 1 0 684 0 1 1035
box -2 -2 2 2
use M2_M1  M2_M1_9320
timestamp 1745462530
transform 1 0 428 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_9321
timestamp 1745462530
transform 1 0 412 0 1 945
box -2 -2 2 2
use M2_M1  M2_M1_9322
timestamp 1745462530
transform 1 0 332 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_9323
timestamp 1745462530
transform 1 0 484 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_9324
timestamp 1745462530
transform 1 0 452 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_9325
timestamp 1745462530
transform 1 0 836 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_9326
timestamp 1745462530
transform 1 0 508 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_9327
timestamp 1745462530
transform 1 0 500 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_9328
timestamp 1745462530
transform 1 0 452 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_9329
timestamp 1745462530
transform 1 0 356 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_9330
timestamp 1745462530
transform 1 0 356 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_9331
timestamp 1745462530
transform 1 0 316 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_9332
timestamp 1745462530
transform 1 0 300 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_9333
timestamp 1745462530
transform 1 0 916 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_9334
timestamp 1745462530
transform 1 0 540 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_9335
timestamp 1745462530
transform 1 0 500 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_9336
timestamp 1745462530
transform 1 0 412 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_9337
timestamp 1745462530
transform 1 0 412 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_9338
timestamp 1745462530
transform 1 0 388 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_9339
timestamp 1745462530
transform 1 0 348 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_9340
timestamp 1745462530
transform 1 0 348 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_9341
timestamp 1745462530
transform 1 0 836 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_9342
timestamp 1745462530
transform 1 0 468 0 1 845
box -2 -2 2 2
use M2_M1  M2_M1_9343
timestamp 1745462530
transform 1 0 468 0 1 785
box -2 -2 2 2
use M2_M1  M2_M1_9344
timestamp 1745462530
transform 1 0 460 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_9345
timestamp 1745462530
transform 1 0 420 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_9346
timestamp 1745462530
transform 1 0 404 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_9347
timestamp 1745462530
transform 1 0 308 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_9348
timestamp 1745462530
transform 1 0 300 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_9349
timestamp 1745462530
transform 1 0 276 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_9350
timestamp 1745462530
transform 1 0 900 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_9351
timestamp 1745462530
transform 1 0 516 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_9352
timestamp 1745462530
transform 1 0 516 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_9353
timestamp 1745462530
transform 1 0 436 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_9354
timestamp 1745462530
transform 1 0 436 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_9355
timestamp 1745462530
transform 1 0 356 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_9356
timestamp 1745462530
transform 1 0 348 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_9357
timestamp 1745462530
transform 1 0 324 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_9358
timestamp 1745462530
transform 1 0 972 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_9359
timestamp 1745462530
transform 1 0 916 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_9360
timestamp 1745462530
transform 1 0 892 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_9361
timestamp 1745462530
transform 1 0 892 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_9362
timestamp 1745462530
transform 1 0 764 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_9363
timestamp 1745462530
transform 1 0 748 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_9364
timestamp 1745462530
transform 1 0 708 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_9365
timestamp 1745462530
transform 1 0 684 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_9366
timestamp 1745462530
transform 1 0 684 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_9367
timestamp 1745462530
transform 1 0 1020 0 1 1085
box -2 -2 2 2
use M2_M1  M2_M1_9368
timestamp 1745462530
transform 1 0 964 0 1 1115
box -2 -2 2 2
use M2_M1  M2_M1_9369
timestamp 1745462530
transform 1 0 940 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_9370
timestamp 1745462530
transform 1 0 908 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_9371
timestamp 1745462530
transform 1 0 812 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_9372
timestamp 1745462530
transform 1 0 796 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_9373
timestamp 1745462530
transform 1 0 764 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_9374
timestamp 1745462530
transform 1 0 716 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_9375
timestamp 1745462530
transform 1 0 700 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_9376
timestamp 1745462530
transform 1 0 1124 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_9377
timestamp 1745462530
transform 1 0 1044 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_9378
timestamp 1745462530
transform 1 0 988 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_9379
timestamp 1745462530
transform 1 0 804 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_9380
timestamp 1745462530
transform 1 0 804 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_9381
timestamp 1745462530
transform 1 0 748 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_9382
timestamp 1745462530
transform 1 0 676 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_9383
timestamp 1745462530
transform 1 0 628 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_9384
timestamp 1745462530
transform 1 0 1164 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_9385
timestamp 1745462530
transform 1 0 1092 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_9386
timestamp 1745462530
transform 1 0 1028 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_9387
timestamp 1745462530
transform 1 0 836 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_9388
timestamp 1745462530
transform 1 0 836 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_9389
timestamp 1745462530
transform 1 0 764 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_9390
timestamp 1745462530
transform 1 0 700 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_9391
timestamp 1745462530
transform 1 0 668 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_9392
timestamp 1745462530
transform 1 0 2564 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_9393
timestamp 1745462530
transform 1 0 1652 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_9394
timestamp 1745462530
transform 1 0 1620 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_9395
timestamp 1745462530
transform 1 0 1516 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_9396
timestamp 1745462530
transform 1 0 1492 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_9397
timestamp 1745462530
transform 1 0 1500 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_9398
timestamp 1745462530
transform 1 0 1404 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_9399
timestamp 1745462530
transform 1 0 3044 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_9400
timestamp 1745462530
transform 1 0 1484 0 1 1585
box -2 -2 2 2
use M2_M1  M2_M1_9401
timestamp 1745462530
transform 1 0 3020 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_9402
timestamp 1745462530
transform 1 0 3004 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_9403
timestamp 1745462530
transform 1 0 3156 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_9404
timestamp 1745462530
transform 1 0 3156 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_9405
timestamp 1745462530
transform 1 0 3148 0 1 985
box -2 -2 2 2
use M2_M1  M2_M1_9406
timestamp 1745462530
transform 1 0 3012 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_9407
timestamp 1745462530
transform 1 0 3140 0 1 795
box -2 -2 2 2
use M2_M1  M2_M1_9408
timestamp 1745462530
transform 1 0 3028 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_9409
timestamp 1745462530
transform 1 0 3308 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_9410
timestamp 1745462530
transform 1 0 3164 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_9411
timestamp 1745462530
transform 1 0 3332 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_9412
timestamp 1745462530
transform 1 0 3268 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_9413
timestamp 1745462530
transform 1 0 3340 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_9414
timestamp 1745462530
transform 1 0 3276 0 1 835
box -2 -2 2 2
use M2_M1  M2_M1_9415
timestamp 1745462530
transform 1 0 3332 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_9416
timestamp 1745462530
transform 1 0 3292 0 1 835
box -2 -2 2 2
use M2_M1  M2_M1_9417
timestamp 1745462530
transform 1 0 3308 0 1 545
box -2 -2 2 2
use M2_M1  M2_M1_9418
timestamp 1745462530
transform 1 0 3284 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_9419
timestamp 1745462530
transform 1 0 3380 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_9420
timestamp 1745462530
transform 1 0 3356 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_9421
timestamp 1745462530
transform 1 0 3012 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_9422
timestamp 1745462530
transform 1 0 3004 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_9423
timestamp 1745462530
transform 1 0 3060 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_9424
timestamp 1745462530
transform 1 0 3012 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_9425
timestamp 1745462530
transform 1 0 2996 0 1 785
box -2 -2 2 2
use M2_M1  M2_M1_9426
timestamp 1745462530
transform 1 0 2996 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_9427
timestamp 1745462530
transform 1 0 2964 0 1 745
box -2 -2 2 2
use M2_M1  M2_M1_9428
timestamp 1745462530
transform 1 0 2940 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_9429
timestamp 1745462530
transform 1 0 2996 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_9430
timestamp 1745462530
transform 1 0 2844 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_9431
timestamp 1745462530
transform 1 0 3108 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_9432
timestamp 1745462530
transform 1 0 3044 0 1 1745
box -2 -2 2 2
use M2_M1  M2_M1_9433
timestamp 1745462530
transform 1 0 3164 0 1 2625
box -2 -2 2 2
use M2_M1  M2_M1_9434
timestamp 1745462530
transform 1 0 3068 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_9435
timestamp 1745462530
transform 1 0 3132 0 1 2625
box -2 -2 2 2
use M2_M1  M2_M1_9436
timestamp 1745462530
transform 1 0 3020 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_9437
timestamp 1745462530
transform 1 0 3148 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_9438
timestamp 1745462530
transform 1 0 3108 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_9439
timestamp 1745462530
transform 1 0 3188 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_9440
timestamp 1745462530
transform 1 0 3156 0 1 2635
box -2 -2 2 2
use M2_M1  M2_M1_9441
timestamp 1745462530
transform 1 0 3212 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_9442
timestamp 1745462530
transform 1 0 3204 0 1 2545
box -2 -2 2 2
use M2_M1  M2_M1_9443
timestamp 1745462530
transform 1 0 3068 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_9444
timestamp 1745462530
transform 1 0 2932 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_9445
timestamp 1745462530
transform 1 0 3212 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_9446
timestamp 1745462530
transform 1 0 3084 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_9447
timestamp 1745462530
transform 1 0 3356 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_9448
timestamp 1745462530
transform 1 0 3092 0 1 1705
box -2 -2 2 2
use M2_M1  M2_M1_9449
timestamp 1745462530
transform 1 0 3420 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_9450
timestamp 1745462530
transform 1 0 3372 0 1 1595
box -2 -2 2 2
use M2_M1  M2_M1_9451
timestamp 1745462530
transform 1 0 3484 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_9452
timestamp 1745462530
transform 1 0 3388 0 1 1595
box -2 -2 2 2
use M2_M1  M2_M1_9453
timestamp 1745462530
transform 1 0 1452 0 1 2395
box -2 -2 2 2
use M2_M1  M2_M1_9454
timestamp 1745462530
transform 1 0 1412 0 1 2145
box -2 -2 2 2
use M2_M1  M2_M1_9455
timestamp 1745462530
transform 1 0 1436 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_9456
timestamp 1745462530
transform 1 0 772 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_9457
timestamp 1745462530
transform 1 0 796 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_9458
timestamp 1745462530
transform 1 0 724 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_9459
timestamp 1745462530
transform 1 0 740 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_9460
timestamp 1745462530
transform 1 0 652 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_9461
timestamp 1745462530
transform 1 0 748 0 1 2105
box -2 -2 2 2
use M2_M1  M2_M1_9462
timestamp 1745462530
transform 1 0 708 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_9463
timestamp 1745462530
transform 1 0 692 0 1 2795
box -2 -2 2 2
use M2_M1  M2_M1_9464
timestamp 1745462530
transform 1 0 668 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_9465
timestamp 1745462530
transform 1 0 748 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_9466
timestamp 1745462530
transform 1 0 732 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_9467
timestamp 1745462530
transform 1 0 1388 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_9468
timestamp 1745462530
transform 1 0 1364 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_9469
timestamp 1745462530
transform 1 0 1436 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_9470
timestamp 1745462530
transform 1 0 1428 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_9471
timestamp 1745462530
transform 1 0 1420 0 1 2435
box -2 -2 2 2
use M2_M1  M2_M1_9472
timestamp 1745462530
transform 1 0 1316 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_9473
timestamp 1745462530
transform 1 0 1292 0 1 2345
box -2 -2 2 2
use M2_M1  M2_M1_9474
timestamp 1745462530
transform 1 0 1268 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_9475
timestamp 1745462530
transform 1 0 1324 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_9476
timestamp 1745462530
transform 1 0 1204 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_9477
timestamp 1745462530
transform 1 0 1524 0 1 945
box -2 -2 2 2
use M2_M1  M2_M1_9478
timestamp 1745462530
transform 1 0 708 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_9479
timestamp 1745462530
transform 1 0 1540 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_9480
timestamp 1745462530
transform 1 0 1524 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_9481
timestamp 1745462530
transform 1 0 1500 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_9482
timestamp 1745462530
transform 1 0 1476 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_9483
timestamp 1745462530
transform 1 0 1484 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_9484
timestamp 1745462530
transform 1 0 1484 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_9485
timestamp 1745462530
transform 1 0 1460 0 1 905
box -2 -2 2 2
use M2_M1  M2_M1_9486
timestamp 1745462530
transform 1 0 1460 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_9487
timestamp 1745462530
transform 1 0 1460 0 1 595
box -2 -2 2 2
use M2_M1  M2_M1_9488
timestamp 1745462530
transform 1 0 1364 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_9489
timestamp 1745462530
transform 1 0 1492 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_9490
timestamp 1745462530
transform 1 0 1436 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_9491
timestamp 1745462530
transform 1 0 692 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_9492
timestamp 1745462530
transform 1 0 676 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_9493
timestamp 1745462530
transform 1 0 692 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_9494
timestamp 1745462530
transform 1 0 692 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_9495
timestamp 1745462530
transform 1 0 668 0 1 835
box -2 -2 2 2
use M2_M1  M2_M1_9496
timestamp 1745462530
transform 1 0 556 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_9497
timestamp 1745462530
transform 1 0 524 0 1 795
box -2 -2 2 2
use M2_M1  M2_M1_9498
timestamp 1745462530
transform 1 0 500 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_9499
timestamp 1745462530
transform 1 0 540 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_9500
timestamp 1745462530
transform 1 0 388 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_9501
timestamp 1745462530
transform 1 0 2164 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_9502
timestamp 1745462530
transform 1 0 1772 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_9503
timestamp 1745462530
transform 1 0 1644 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_9504
timestamp 1745462530
transform 1 0 1684 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_9505
timestamp 1745462530
transform 1 0 1684 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_9506
timestamp 1745462530
transform 1 0 1684 0 1 1635
box -2 -2 2 2
use M2_M1  M2_M1_9507
timestamp 1745462530
transform 1 0 1596 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_9508
timestamp 1745462530
transform 1 0 1596 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_9509
timestamp 1745462530
transform 1 0 1580 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_9510
timestamp 1745462530
transform 1 0 3084 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_9511
timestamp 1745462530
transform 1 0 1732 0 1 1635
box -2 -2 2 2
use M2_M1  M2_M1_9512
timestamp 1745462530
transform 1 0 3452 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_9513
timestamp 1745462530
transform 1 0 3060 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_9514
timestamp 1745462530
transform 1 0 3188 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_9515
timestamp 1745462530
transform 1 0 3068 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_9516
timestamp 1745462530
transform 1 0 3148 0 1 955
box -2 -2 2 2
use M2_M1  M2_M1_9517
timestamp 1745462530
transform 1 0 2444 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_9518
timestamp 1745462530
transform 1 0 3884 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_9519
timestamp 1745462530
transform 1 0 3188 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_9520
timestamp 1745462530
transform 1 0 3884 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_9521
timestamp 1745462530
transform 1 0 3860 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_9522
timestamp 1745462530
transform 1 0 3932 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_9523
timestamp 1745462530
transform 1 0 3868 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_9524
timestamp 1745462530
transform 1 0 3892 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_9525
timestamp 1745462530
transform 1 0 3876 0 1 905
box -2 -2 2 2
use M2_M1  M2_M1_9526
timestamp 1745462530
transform 1 0 3844 0 1 395
box -2 -2 2 2
use M2_M1  M2_M1_9527
timestamp 1745462530
transform 1 0 3820 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_9528
timestamp 1745462530
transform 1 0 3924 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_9529
timestamp 1745462530
transform 1 0 3908 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9530
timestamp 1745462530
transform 1 0 2451 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_9531
timestamp 1745462530
transform 1 0 2420 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_9532
timestamp 1745462530
transform 1 0 2484 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_9533
timestamp 1745462530
transform 1 0 2428 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_9534
timestamp 1745462530
transform 1 0 2436 0 1 905
box -2 -2 2 2
use M2_M1  M2_M1_9535
timestamp 1745462530
transform 1 0 2428 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_9536
timestamp 1745462530
transform 1 0 2420 0 1 595
box -2 -2 2 2
use M2_M1  M2_M1_9537
timestamp 1745462530
transform 1 0 2268 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_9538
timestamp 1745462530
transform 1 0 2452 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_9539
timestamp 1745462530
transform 1 0 2404 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_9540
timestamp 1745462530
transform 1 0 4060 0 1 2625
box -2 -2 2 2
use M2_M1  M2_M1_9541
timestamp 1745462530
transform 1 0 3468 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_9542
timestamp 1745462530
transform 1 0 4044 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_9543
timestamp 1745462530
transform 1 0 4036 0 1 2625
box -2 -2 2 2
use M2_M1  M2_M1_9544
timestamp 1745462530
transform 1 0 4020 0 1 2635
box -2 -2 2 2
use M2_M1  M2_M1_9545
timestamp 1745462530
transform 1 0 3996 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_9546
timestamp 1745462530
transform 1 0 4076 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_9547
timestamp 1745462530
transform 1 0 4052 0 1 2635
box -2 -2 2 2
use M2_M1  M2_M1_9548
timestamp 1745462530
transform 1 0 4156 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_9549
timestamp 1745462530
transform 1 0 4084 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_9550
timestamp 1745462530
transform 1 0 3380 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_9551
timestamp 1745462530
transform 1 0 2868 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_9552
timestamp 1745462530
transform 1 0 3420 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_9553
timestamp 1745462530
transform 1 0 3356 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_9554
timestamp 1745462530
transform 1 0 3516 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_9555
timestamp 1745462530
transform 1 0 3428 0 1 1705
box -2 -2 2 2
use M2_M1  M2_M1_9556
timestamp 1745462530
transform 1 0 3588 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_9557
timestamp 1745462530
transform 1 0 3548 0 1 1545
box -2 -2 2 2
use M2_M1  M2_M1_9558
timestamp 1745462530
transform 1 0 3636 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_9559
timestamp 1745462530
transform 1 0 3612 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_9560
timestamp 1745462530
transform 1 0 1620 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_9561
timestamp 1745462530
transform 1 0 1604 0 1 2195
box -2 -2 2 2
use M2_M1  M2_M1_9562
timestamp 1745462530
transform 1 0 1628 0 1 2195
box -2 -2 2 2
use M2_M1  M2_M1_9563
timestamp 1745462530
transform 1 0 724 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_9564
timestamp 1745462530
transform 1 0 676 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_9565
timestamp 1745462530
transform 1 0 660 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_9566
timestamp 1745462530
transform 1 0 692 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_9567
timestamp 1745462530
transform 1 0 596 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_9568
timestamp 1745462530
transform 1 0 700 0 1 2105
box -2 -2 2 2
use M2_M1  M2_M1_9569
timestamp 1745462530
transform 1 0 684 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_9570
timestamp 1745462530
transform 1 0 668 0 1 2595
box -2 -2 2 2
use M2_M1  M2_M1_9571
timestamp 1745462530
transform 1 0 644 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_9572
timestamp 1745462530
transform 1 0 732 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_9573
timestamp 1745462530
transform 1 0 700 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_9574
timestamp 1745462530
transform 1 0 1668 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_9575
timestamp 1745462530
transform 1 0 1596 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_9576
timestamp 1745462530
transform 1 0 1668 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_9577
timestamp 1745462530
transform 1 0 1604 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_9578
timestamp 1745462530
transform 1 0 1612 0 1 2435
box -2 -2 2 2
use M2_M1  M2_M1_9579
timestamp 1745462530
transform 1 0 1596 0 1 2345
box -2 -2 2 2
use M2_M1  M2_M1_9580
timestamp 1745462530
transform 1 0 1668 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_9581
timestamp 1745462530
transform 1 0 1612 0 1 2345
box -2 -2 2 2
use M2_M1  M2_M1_9582
timestamp 1745462530
transform 1 0 1628 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_9583
timestamp 1745462530
transform 1 0 1572 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_9584
timestamp 1745462530
transform 1 0 1708 0 1 945
box -2 -2 2 2
use M2_M1  M2_M1_9585
timestamp 1745462530
transform 1 0 772 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_9586
timestamp 1745462530
transform 1 0 1876 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_9587
timestamp 1745462530
transform 1 0 1732 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_9588
timestamp 1745462530
transform 1 0 1908 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_9589
timestamp 1745462530
transform 1 0 1836 0 1 905
box -2 -2 2 2
use M2_M1  M2_M1_9590
timestamp 1745462530
transform 1 0 1908 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_9591
timestamp 1745462530
transform 1 0 1852 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_9592
timestamp 1745462530
transform 1 0 1860 0 1 905
box -2 -2 2 2
use M2_M1  M2_M1_9593
timestamp 1745462530
transform 1 0 1860 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_9594
timestamp 1745462530
transform 1 0 1868 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_9595
timestamp 1745462530
transform 1 0 1852 0 1 595
box -2 -2 2 2
use M2_M1  M2_M1_9596
timestamp 1745462530
transform 1 0 1876 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_9597
timestamp 1745462530
transform 1 0 1812 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_9598
timestamp 1745462530
transform 1 0 756 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_9599
timestamp 1745462530
transform 1 0 732 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_9600
timestamp 1745462530
transform 1 0 756 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_9601
timestamp 1745462530
transform 1 0 740 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_9602
timestamp 1745462530
transform 1 0 716 0 1 835
box -2 -2 2 2
use M2_M1  M2_M1_9603
timestamp 1745462530
transform 1 0 492 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_9604
timestamp 1745462530
transform 1 0 444 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_9605
timestamp 1745462530
transform 1 0 420 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_9606
timestamp 1745462530
transform 1 0 476 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_9607
timestamp 1745462530
transform 1 0 372 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_9608
timestamp 1745462530
transform 1 0 2140 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_9609
timestamp 1745462530
transform 1 0 1844 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_9610
timestamp 1745462530
transform 1 0 1844 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_9611
timestamp 1745462530
transform 1 0 1908 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_9612
timestamp 1745462530
transform 1 0 1884 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_9613
timestamp 1745462530
transform 1 0 1908 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_9614
timestamp 1745462530
transform 1 0 1876 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_9615
timestamp 1745462530
transform 1 0 3588 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_9616
timestamp 1745462530
transform 1 0 3372 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_9617
timestamp 1745462530
transform 1 0 3348 0 1 1585
box -2 -2 2 2
use M2_M1  M2_M1_9618
timestamp 1745462530
transform 1 0 1884 0 1 1705
box -2 -2 2 2
use M2_M1  M2_M1_9619
timestamp 1745462530
transform 1 0 3748 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_9620
timestamp 1745462530
transform 1 0 3556 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_9621
timestamp 1745462530
transform 1 0 3564 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_9622
timestamp 1745462530
transform 1 0 3556 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_9623
timestamp 1745462530
transform 1 0 3548 0 1 795
box -2 -2 2 2
use M2_M1  M2_M1_9624
timestamp 1745462530
transform 1 0 2580 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_9625
timestamp 1745462530
transform 1 0 3772 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_9626
timestamp 1745462530
transform 1 0 3572 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_9627
timestamp 1745462530
transform 1 0 3748 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_9628
timestamp 1745462530
transform 1 0 3684 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_9629
timestamp 1745462530
transform 1 0 3876 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_9630
timestamp 1745462530
transform 1 0 3740 0 1 835
box -2 -2 2 2
use M2_M1  M2_M1_9631
timestamp 1745462530
transform 1 0 3764 0 1 835
box -2 -2 2 2
use M2_M1  M2_M1_9632
timestamp 1745462530
transform 1 0 3668 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_9633
timestamp 1745462530
transform 1 0 3660 0 1 595
box -2 -2 2 2
use M2_M1  M2_M1_9634
timestamp 1745462530
transform 1 0 3620 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_9635
timestamp 1745462530
transform 1 0 3724 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_9636
timestamp 1745462530
transform 1 0 3692 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_9637
timestamp 1745462530
transform 1 0 2548 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_9638
timestamp 1745462530
transform 1 0 2540 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_9639
timestamp 1745462530
transform 1 0 2540 0 1 835
box -2 -2 2 2
use M2_M1  M2_M1_9640
timestamp 1745462530
transform 1 0 2516 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_9641
timestamp 1745462530
transform 1 0 2572 0 1 835
box -2 -2 2 2
use M2_M1  M2_M1_9642
timestamp 1745462530
transform 1 0 2572 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_9643
timestamp 1745462530
transform 1 0 2556 0 1 745
box -2 -2 2 2
use M2_M1  M2_M1_9644
timestamp 1745462530
transform 1 0 2476 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_9645
timestamp 1745462530
transform 1 0 2588 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_9646
timestamp 1745462530
transform 1 0 2524 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_9647
timestamp 1745462530
transform 1 0 3780 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_9648
timestamp 1745462530
transform 1 0 3772 0 1 1745
box -2 -2 2 2
use M2_M1  M2_M1_9649
timestamp 1745462530
transform 1 0 3812 0 1 2625
box -2 -2 2 2
use M2_M1  M2_M1_9650
timestamp 1745462530
transform 1 0 3788 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_9651
timestamp 1745462530
transform 1 0 3804 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_9652
timestamp 1745462530
transform 1 0 3788 0 1 2625
box -2 -2 2 2
use M2_M1  M2_M1_9653
timestamp 1745462530
transform 1 0 3796 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_9654
timestamp 1745462530
transform 1 0 3756 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_9655
timestamp 1745462530
transform 1 0 3852 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_9656
timestamp 1745462530
transform 1 0 3804 0 1 2635
box -2 -2 2 2
use M2_M1  M2_M1_9657
timestamp 1745462530
transform 1 0 3900 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_9658
timestamp 1745462530
transform 1 0 3852 0 1 2595
box -2 -2 2 2
use M2_M1  M2_M1_9659
timestamp 1745462530
transform 1 0 3748 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_9660
timestamp 1745462530
transform 1 0 2996 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_9661
timestamp 1745462530
transform 1 0 3812 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_9662
timestamp 1745462530
transform 1 0 3748 0 1 1635
box -2 -2 2 2
use M2_M1  M2_M1_9663
timestamp 1745462530
transform 1 0 3812 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_9664
timestamp 1745462530
transform 1 0 3772 0 1 1635
box -2 -2 2 2
use M2_M1  M2_M1_9665
timestamp 1745462530
transform 1 0 3892 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_9666
timestamp 1745462530
transform 1 0 3820 0 1 1545
box -2 -2 2 2
use M2_M1  M2_M1_9667
timestamp 1745462530
transform 1 0 3884 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_9668
timestamp 1745462530
transform 1 0 3868 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_9669
timestamp 1745462530
transform 1 0 1884 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_9670
timestamp 1745462530
transform 1 0 1868 0 1 2145
box -2 -2 2 2
use M2_M1  M2_M1_9671
timestamp 1745462530
transform 1 0 1884 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_9672
timestamp 1745462530
transform 1 0 860 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_9673
timestamp 1745462530
transform 1 0 852 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_9674
timestamp 1745462530
transform 1 0 836 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_9675
timestamp 1745462530
transform 1 0 844 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_9676
timestamp 1745462530
transform 1 0 796 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_9677
timestamp 1745462530
transform 1 0 852 0 1 2795
box -2 -2 2 2
use M2_M1  M2_M1_9678
timestamp 1745462530
transform 1 0 852 0 1 2105
box -2 -2 2 2
use M2_M1  M2_M1_9679
timestamp 1745462530
transform 1 0 820 0 1 2795
box -2 -2 2 2
use M2_M1  M2_M1_9680
timestamp 1745462530
transform 1 0 796 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_9681
timestamp 1745462530
transform 1 0 876 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_9682
timestamp 1745462530
transform 1 0 860 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_9683
timestamp 1745462530
transform 1 0 1916 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_9684
timestamp 1745462530
transform 1 0 1852 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_9685
timestamp 1745462530
transform 1 0 1940 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_9686
timestamp 1745462530
transform 1 0 1860 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_9687
timestamp 1745462530
transform 1 0 1836 0 1 2435
box -2 -2 2 2
use M2_M1  M2_M1_9688
timestamp 1745462530
transform 1 0 1836 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_9689
timestamp 1745462530
transform 1 0 1876 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_9690
timestamp 1745462530
transform 1 0 1828 0 1 2345
box -2 -2 2 2
use M2_M1  M2_M1_9691
timestamp 1745462530
transform 1 0 1844 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_9692
timestamp 1745462530
transform 1 0 1788 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_9693
timestamp 1745462530
transform 1 0 1908 0 1 795
box -2 -2 2 2
use M2_M1  M2_M1_9694
timestamp 1745462530
transform 1 0 908 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_9695
timestamp 1745462530
transform 1 0 2028 0 1 845
box -2 -2 2 2
use M2_M1  M2_M1_9696
timestamp 1745462530
transform 1 0 1940 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_9697
timestamp 1745462530
transform 1 0 2076 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_9698
timestamp 1745462530
transform 1 0 1996 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_9699
timestamp 1745462530
transform 1 0 1988 0 1 835
box -2 -2 2 2
use M2_M1  M2_M1_9700
timestamp 1745462530
transform 1 0 1964 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_9701
timestamp 1745462530
transform 1 0 2044 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_9702
timestamp 1745462530
transform 1 0 2012 0 1 835
box -2 -2 2 2
use M2_M1  M2_M1_9703
timestamp 1745462530
transform 1 0 2020 0 1 545
box -2 -2 2 2
use M2_M1  M2_M1_9704
timestamp 1745462530
transform 1 0 1940 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_9705
timestamp 1745462530
transform 1 0 2060 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_9706
timestamp 1745462530
transform 1 0 1956 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_9707
timestamp 1745462530
transform 1 0 828 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_9708
timestamp 1745462530
transform 1 0 828 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_9709
timestamp 1745462530
transform 1 0 932 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_9710
timestamp 1745462530
transform 1 0 860 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_9711
timestamp 1745462530
transform 1 0 836 0 1 835
box -2 -2 2 2
use M2_M1  M2_M1_9712
timestamp 1745462530
transform 1 0 396 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_9713
timestamp 1745462530
transform 1 0 340 0 1 745
box -2 -2 2 2
use M2_M1  M2_M1_9714
timestamp 1745462530
transform 1 0 316 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_9715
timestamp 1745462530
transform 1 0 372 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_9716
timestamp 1745462530
transform 1 0 316 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_9717
timestamp 1745462530
transform 1 0 2364 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_9718
timestamp 1745462530
transform 1 0 1244 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_9719
timestamp 1745462530
transform 1 0 1148 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_9720
timestamp 1745462530
transform 1 0 1220 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_9721
timestamp 1745462530
transform 1 0 1108 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_9722
timestamp 1745462530
transform 1 0 3252 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_9723
timestamp 1745462530
transform 1 0 1100 0 1 2245
box -2 -2 2 2
use M2_M1  M2_M1_9724
timestamp 1745462530
transform 1 0 3260 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_9725
timestamp 1745462530
transform 1 0 3204 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_9726
timestamp 1745462530
transform 1 0 3228 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_9727
timestamp 1745462530
transform 1 0 3212 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_9728
timestamp 1745462530
transform 1 0 3244 0 1 795
box -2 -2 2 2
use M2_M1  M2_M1_9729
timestamp 1745462530
transform 1 0 2620 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_9730
timestamp 1745462530
transform 1 0 3460 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_9731
timestamp 1745462530
transform 1 0 3268 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_9732
timestamp 1745462530
transform 1 0 3548 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_9733
timestamp 1745462530
transform 1 0 3420 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_9734
timestamp 1745462530
transform 1 0 3500 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_9735
timestamp 1745462530
transform 1 0 3444 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_9736
timestamp 1745462530
transform 1 0 3460 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_9737
timestamp 1745462530
transform 1 0 3452 0 1 835
box -2 -2 2 2
use M2_M1  M2_M1_9738
timestamp 1745462530
transform 1 0 3460 0 1 595
box -2 -2 2 2
use M2_M1  M2_M1_9739
timestamp 1745462530
transform 1 0 3460 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_9740
timestamp 1745462530
transform 1 0 3580 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_9741
timestamp 1745462530
transform 1 0 3500 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_9742
timestamp 1745462530
transform 1 0 2588 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_9743
timestamp 1745462530
transform 1 0 2516 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_9744
timestamp 1745462530
transform 1 0 2643 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_9745
timestamp 1745462530
transform 1 0 2588 0 1 835
box -2 -2 2 2
use M2_M1  M2_M1_9746
timestamp 1745462530
transform 1 0 2604 0 1 835
box -2 -2 2 2
use M2_M1  M2_M1_9747
timestamp 1745462530
transform 1 0 2500 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_9748
timestamp 1745462530
transform 1 0 2452 0 1 595
box -2 -2 2 2
use M2_M1  M2_M1_9749
timestamp 1745462530
transform 1 0 2332 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_9750
timestamp 1745462530
transform 1 0 2484 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_9751
timestamp 1745462530
transform 1 0 2468 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_9752
timestamp 1745462530
transform 1 0 3324 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_9753
timestamp 1745462530
transform 1 0 3236 0 1 2145
box -2 -2 2 2
use M2_M1  M2_M1_9754
timestamp 1745462530
transform 1 0 3364 0 1 2715
box -2 -2 2 2
use M2_M1  M2_M1_9755
timestamp 1745462530
transform 1 0 3284 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_9756
timestamp 1745462530
transform 1 0 3332 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_9757
timestamp 1745462530
transform 1 0 3324 0 1 2715
box -2 -2 2 2
use M2_M1  M2_M1_9758
timestamp 1745462530
transform 1 0 3388 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_9759
timestamp 1745462530
transform 1 0 3332 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_9760
timestamp 1745462530
transform 1 0 3356 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_9761
timestamp 1745462530
transform 1 0 3340 0 1 2705
box -2 -2 2 2
use M2_M1  M2_M1_9762
timestamp 1745462530
transform 1 0 3388 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_9763
timestamp 1745462530
transform 1 0 3372 0 1 2595
box -2 -2 2 2
use M2_M1  M2_M1_9764
timestamp 1745462530
transform 1 0 3292 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_9765
timestamp 1745462530
transform 1 0 2948 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_9766
timestamp 1745462530
transform 1 0 3452 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_9767
timestamp 1745462530
transform 1 0 3308 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_9768
timestamp 1745462530
transform 1 0 3476 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_9769
timestamp 1745462530
transform 1 0 3316 0 1 2035
box -2 -2 2 2
use M2_M1  M2_M1_9770
timestamp 1745462530
transform 1 0 3532 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_9771
timestamp 1745462530
transform 1 0 3468 0 1 1945
box -2 -2 2 2
use M2_M1  M2_M1_9772
timestamp 1745462530
transform 1 0 3660 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_9773
timestamp 1745462530
transform 1 0 3484 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_9774
timestamp 1745462530
transform 1 0 1116 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_9775
timestamp 1745462530
transform 1 0 1076 0 1 2195
box -2 -2 2 2
use M2_M1  M2_M1_9776
timestamp 1745462530
transform 1 0 1092 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_9777
timestamp 1745462530
transform 1 0 900 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_9778
timestamp 1745462530
transform 1 0 924 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_9779
timestamp 1745462530
transform 1 0 860 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_9780
timestamp 1745462530
transform 1 0 852 0 1 2235
box -2 -2 2 2
use M2_M1  M2_M1_9781
timestamp 1745462530
transform 1 0 828 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_9782
timestamp 1745462530
transform 1 0 884 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_9783
timestamp 1745462530
transform 1 0 876 0 1 2235
box -2 -2 2 2
use M2_M1  M2_M1_9784
timestamp 1745462530
transform 1 0 892 0 1 2595
box -2 -2 2 2
use M2_M1  M2_M1_9785
timestamp 1745462530
transform 1 0 860 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_9786
timestamp 1745462530
transform 1 0 908 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_9787
timestamp 1745462530
transform 1 0 892 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_9788
timestamp 1745462530
transform 1 0 1196 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_9789
timestamp 1745462530
transform 1 0 1092 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_9790
timestamp 1745462530
transform 1 0 1452 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_9791
timestamp 1745462530
transform 1 0 1100 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_9792
timestamp 1745462530
transform 1 0 1124 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_9793
timestamp 1745462530
transform 1 0 1108 0 1 2435
box -2 -2 2 2
use M2_M1  M2_M1_9794
timestamp 1745462530
transform 1 0 1260 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_9795
timestamp 1745462530
transform 1 0 1140 0 1 2395
box -2 -2 2 2
use M2_M1  M2_M1_9796
timestamp 1745462530
transform 1 0 1156 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_9797
timestamp 1745462530
transform 1 0 1140 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_9798
timestamp 1745462530
transform 1 0 1172 0 1 1145
box -2 -2 2 2
use M2_M1  M2_M1_9799
timestamp 1745462530
transform 1 0 852 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_9800
timestamp 1745462530
transform 1 0 1252 0 1 1115
box -2 -2 2 2
use M2_M1  M2_M1_9801
timestamp 1745462530
transform 1 0 1236 0 1 1105
box -2 -2 2 2
use M2_M1  M2_M1_9802
timestamp 1745462530
transform 1 0 1268 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_9803
timestamp 1745462530
transform 1 0 1228 0 1 1115
box -2 -2 2 2
use M2_M1  M2_M1_9804
timestamp 1745462530
transform 1 0 1236 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_9805
timestamp 1745462530
transform 1 0 1236 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_9806
timestamp 1745462530
transform 1 0 1244 0 1 1105
box -2 -2 2 2
use M2_M1  M2_M1_9807
timestamp 1745462530
transform 1 0 1212 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_9808
timestamp 1745462530
transform 1 0 1188 0 1 595
box -2 -2 2 2
use M2_M1  M2_M1_9809
timestamp 1745462530
transform 1 0 1180 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_9810
timestamp 1745462530
transform 1 0 1324 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_9811
timestamp 1745462530
transform 1 0 1244 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_9812
timestamp 1745462530
transform 1 0 996 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_9813
timestamp 1745462530
transform 1 0 820 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_9814
timestamp 1745462530
transform 1 0 900 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_9815
timestamp 1745462530
transform 1 0 820 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_9816
timestamp 1745462530
transform 1 0 812 0 1 1035
box -2 -2 2 2
use M2_M1  M2_M1_9817
timestamp 1745462530
transform 1 0 348 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_9818
timestamp 1745462530
transform 1 0 316 0 1 995
box -2 -2 2 2
use M2_M1  M2_M1_9819
timestamp 1745462530
transform 1 0 292 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_9820
timestamp 1745462530
transform 1 0 340 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_9821
timestamp 1745462530
transform 1 0 332 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_9822
timestamp 1745462530
transform 1 0 2212 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_9823
timestamp 1745462530
transform 1 0 1508 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_9824
timestamp 1745462530
transform 1 0 1476 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_9825
timestamp 1745462530
transform 1 0 1460 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_9826
timestamp 1745462530
transform 1 0 1460 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_9827
timestamp 1745462530
transform 1 0 1484 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_9828
timestamp 1745462530
transform 1 0 1132 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_9829
timestamp 1745462530
transform 1 0 1476 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_9830
timestamp 1745462530
transform 1 0 1476 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_9831
timestamp 1745462530
transform 1 0 3140 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_9832
timestamp 1745462530
transform 1 0 1508 0 1 2105
box -2 -2 2 2
use M2_M1  M2_M1_9833
timestamp 1745462530
transform 1 0 3476 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_9834
timestamp 1745462530
transform 1 0 3116 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_9835
timestamp 1745462530
transform 1 0 3212 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_9836
timestamp 1745462530
transform 1 0 3124 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_9837
timestamp 1745462530
transform 1 0 3196 0 1 945
box -2 -2 2 2
use M2_M1  M2_M1_9838
timestamp 1745462530
transform 1 0 2884 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_9839
timestamp 1745462530
transform 1 0 3604 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_9840
timestamp 1745462530
transform 1 0 3244 0 1 895
box -2 -2 2 2
use M2_M1  M2_M1_9841
timestamp 1745462530
transform 1 0 3620 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_9842
timestamp 1745462530
transform 1 0 3588 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_9843
timestamp 1745462530
transform 1 0 3644 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_9844
timestamp 1745462530
transform 1 0 3588 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_9845
timestamp 1745462530
transform 1 0 3612 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_9846
timestamp 1745462530
transform 1 0 3596 0 1 835
box -2 -2 2 2
use M2_M1  M2_M1_9847
timestamp 1745462530
transform 1 0 3612 0 1 395
box -2 -2 2 2
use M2_M1  M2_M1_9848
timestamp 1745462530
transform 1 0 3580 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9849
timestamp 1745462530
transform 1 0 3684 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_9850
timestamp 1745462530
transform 1 0 3668 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9851
timestamp 1745462530
transform 1 0 3252 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_9852
timestamp 1745462530
transform 1 0 3236 0 1 1145
box -2 -2 2 2
use M2_M1  M2_M1_9853
timestamp 1745462530
transform 1 0 3188 0 1 1195
box -2 -2 2 2
use M2_M1  M2_M1_9854
timestamp 1745462530
transform 1 0 3188 0 1 1145
box -2 -2 2 2
use M2_M1  M2_M1_9855
timestamp 1745462530
transform 1 0 2668 0 1 1345
box -2 -2 2 2
use M2_M1  M2_M1_9856
timestamp 1745462530
transform 1 0 2260 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_9857
timestamp 1745462530
transform 1 0 3228 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_9858
timestamp 1745462530
transform 1 0 3188 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_9859
timestamp 1745462530
transform 1 0 2748 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_9860
timestamp 1745462530
transform 1 0 2300 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_9861
timestamp 1745462530
transform 1 0 2212 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_9862
timestamp 1745462530
transform 1 0 1412 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_9863
timestamp 1745462530
transform 1 0 1052 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_9864
timestamp 1745462530
transform 1 0 996 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_9865
timestamp 1745462530
transform 1 0 3324 0 1 1785
box -2 -2 2 2
use M2_M1  M2_M1_9866
timestamp 1745462530
transform 1 0 3308 0 1 1785
box -2 -2 2 2
use M2_M1  M2_M1_9867
timestamp 1745462530
transform 1 0 3260 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_9868
timestamp 1745462530
transform 1 0 3260 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_9869
timestamp 1745462530
transform 1 0 2700 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_9870
timestamp 1745462530
transform 1 0 2324 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_9871
timestamp 1745462530
transform 1 0 2228 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_9872
timestamp 1745462530
transform 1 0 1604 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_9873
timestamp 1745462530
transform 1 0 980 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_9874
timestamp 1745462530
transform 1 0 980 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_9875
timestamp 1745462530
transform 1 0 3252 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_9876
timestamp 1745462530
transform 1 0 3212 0 1 1345
box -2 -2 2 2
use M2_M1  M2_M1_9877
timestamp 1745462530
transform 1 0 3188 0 1 1795
box -2 -2 2 2
use M2_M1  M2_M1_9878
timestamp 1745462530
transform 1 0 3172 0 1 1795
box -2 -2 2 2
use M2_M1  M2_M1_9879
timestamp 1745462530
transform 1 0 3156 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_9880
timestamp 1745462530
transform 1 0 2956 0 1 1945
box -2 -2 2 2
use M2_M1  M2_M1_9881
timestamp 1745462530
transform 1 0 2308 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_9882
timestamp 1745462530
transform 1 0 3228 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_9883
timestamp 1745462530
transform 1 0 2932 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_9884
timestamp 1745462530
transform 1 0 2684 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_9885
timestamp 1745462530
transform 1 0 2300 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_9886
timestamp 1745462530
transform 1 0 2284 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_9887
timestamp 1745462530
transform 1 0 1220 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_9888
timestamp 1745462530
transform 1 0 1108 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_9889
timestamp 1745462530
transform 1 0 1060 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_9890
timestamp 1745462530
transform 1 0 3204 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_9891
timestamp 1745462530
transform 1 0 2972 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_9892
timestamp 1745462530
transform 1 0 2900 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_9893
timestamp 1745462530
transform 1 0 2444 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_9894
timestamp 1745462530
transform 1 0 2380 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_9895
timestamp 1745462530
transform 1 0 2052 0 1 2345
box -2 -2 2 2
use M2_M1  M2_M1_9896
timestamp 1745462530
transform 1 0 1236 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_9897
timestamp 1745462530
transform 1 0 1148 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_9898
timestamp 1745462530
transform 1 0 956 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_9899
timestamp 1745462530
transform 1 0 2972 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_9900
timestamp 1745462530
transform 1 0 2956 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_9901
timestamp 1745462530
transform 1 0 2828 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_9902
timestamp 1745462530
transform 1 0 2796 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_9903
timestamp 1745462530
transform 1 0 2844 0 1 905
box -2 -2 2 2
use M2_M1  M2_M1_9904
timestamp 1745462530
transform 1 0 2844 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_9905
timestamp 1745462530
transform 1 0 2860 0 1 905
box -2 -2 2 2
use M2_M1  M2_M1_9906
timestamp 1745462530
transform 1 0 2860 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_9907
timestamp 1745462530
transform 1 0 2804 0 1 595
box -2 -2 2 2
use M2_M1  M2_M1_9908
timestamp 1745462530
transform 1 0 2780 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_9909
timestamp 1745462530
transform 1 0 2836 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_9910
timestamp 1745462530
transform 1 0 2708 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_9911
timestamp 1745462530
transform 1 0 2724 0 1 995
box -2 -2 2 2
use M2_M1  M2_M1_9912
timestamp 1745462530
transform 1 0 2684 0 1 995
box -2 -2 2 2
use M2_M1  M2_M1_9913
timestamp 1745462530
transform 1 0 2676 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_9914
timestamp 1745462530
transform 1 0 2668 0 1 995
box -2 -2 2 2
use M2_M1  M2_M1_9915
timestamp 1745462530
transform 1 0 2404 0 1 1345
box -2 -2 2 2
use M2_M1  M2_M1_9916
timestamp 1745462530
transform 1 0 2284 0 1 1195
box -2 -2 2 2
use M2_M1  M2_M1_9917
timestamp 1745462530
transform 1 0 2212 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_9918
timestamp 1745462530
transform 1 0 3532 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_9919
timestamp 1745462530
transform 1 0 3500 0 1 2145
box -2 -2 2 2
use M2_M1  M2_M1_9920
timestamp 1745462530
transform 1 0 3548 0 1 2625
box -2 -2 2 2
use M2_M1  M2_M1_9921
timestamp 1745462530
transform 1 0 3524 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_9922
timestamp 1745462530
transform 1 0 3564 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_9923
timestamp 1745462530
transform 1 0 3524 0 1 2625
box -2 -2 2 2
use M2_M1  M2_M1_9924
timestamp 1745462530
transform 1 0 3588 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_9925
timestamp 1745462530
transform 1 0 3516 0 1 2635
box -2 -2 2 2
use M2_M1  M2_M1_9926
timestamp 1745462530
transform 1 0 3540 0 1 2635
box -2 -2 2 2
use M2_M1  M2_M1_9927
timestamp 1745462530
transform 1 0 3516 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_9928
timestamp 1745462530
transform 1 0 3540 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_9929
timestamp 1745462530
transform 1 0 3516 0 1 2595
box -2 -2 2 2
use M2_M1  M2_M1_9930
timestamp 1745462530
transform 1 0 2908 0 1 2395
box -2 -2 2 2
use M2_M1  M2_M1_9931
timestamp 1745462530
transform 1 0 2876 0 1 2345
box -2 -2 2 2
use M2_M1  M2_M1_9932
timestamp 1745462530
transform 1 0 2692 0 1 2545
box -2 -2 2 2
use M2_M1  M2_M1_9933
timestamp 1745462530
transform 1 0 2676 0 1 2545
box -2 -2 2 2
use M2_M1  M2_M1_9934
timestamp 1745462530
transform 1 0 2660 0 1 2545
box -2 -2 2 2
use M2_M1  M2_M1_9935
timestamp 1745462530
transform 1 0 2652 0 1 2395
box -2 -2 2 2
use M2_M1  M2_M1_9936
timestamp 1745462530
transform 1 0 2628 0 1 2395
box -2 -2 2 2
use M2_M1  M2_M1_9937
timestamp 1745462530
transform 1 0 2612 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_9938
timestamp 1745462530
transform 1 0 2284 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_9939
timestamp 1745462530
transform 1 0 2692 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_9940
timestamp 1745462530
transform 1 0 2284 0 1 2515
box -2 -2 2 2
use M2_M1  M2_M1_9941
timestamp 1745462530
transform 1 0 2212 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_9942
timestamp 1745462530
transform 1 0 2084 0 1 2545
box -2 -2 2 2
use M2_M1  M2_M1_9943
timestamp 1745462530
transform 1 0 2724 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_9944
timestamp 1745462530
transform 1 0 2636 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_9945
timestamp 1745462530
transform 1 0 2332 0 1 2515
box -2 -2 2 2
use M2_M1  M2_M1_9946
timestamp 1745462530
transform 1 0 2212 0 1 2545
box -2 -2 2 2
use M2_M1  M2_M1_9947
timestamp 1745462530
transform 1 0 2692 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_9948
timestamp 1745462530
transform 1 0 2564 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_9949
timestamp 1745462530
transform 1 0 2332 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_9950
timestamp 1745462530
transform 1 0 2188 0 1 2395
box -2 -2 2 2
use M2_M1  M2_M1_9951
timestamp 1745462530
transform 1 0 2652 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_9952
timestamp 1745462530
transform 1 0 2532 0 1 2395
box -2 -2 2 2
use M2_M1  M2_M1_9953
timestamp 1745462530
transform 1 0 2388 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_9954
timestamp 1745462530
transform 1 0 2140 0 1 2395
box -2 -2 2 2
use M2_M1  M2_M1_9955
timestamp 1745462530
transform 1 0 3508 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_9956
timestamp 1745462530
transform 1 0 3012 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_9957
timestamp 1745462530
transform 1 0 3556 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_9958
timestamp 1745462530
transform 1 0 3508 0 1 2035
box -2 -2 2 2
use M2_M1  M2_M1_9959
timestamp 1745462530
transform 1 0 3684 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_9960
timestamp 1745462530
transform 1 0 3524 0 1 2035
box -2 -2 2 2
use M2_M1  M2_M1_9961
timestamp 1745462530
transform 1 0 3772 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_9962
timestamp 1745462530
transform 1 0 3708 0 1 1945
box -2 -2 2 2
use M2_M1  M2_M1_9963
timestamp 1745462530
transform 1 0 3756 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_9964
timestamp 1745462530
transform 1 0 3724 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_9965
timestamp 1745462530
transform 1 0 1500 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_9966
timestamp 1745462530
transform 1 0 1492 0 1 2195
box -2 -2 2 2
use M2_M1  M2_M1_9967
timestamp 1745462530
transform 1 0 1508 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_9968
timestamp 1745462530
transform 1 0 796 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_9969
timestamp 1745462530
transform 1 0 788 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_9970
timestamp 1745462530
transform 1 0 756 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_9971
timestamp 1745462530
transform 1 0 748 0 1 2235
box -2 -2 2 2
use M2_M1  M2_M1_9972
timestamp 1745462530
transform 1 0 724 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_9973
timestamp 1745462530
transform 1 0 772 0 1 2235
box -2 -2 2 2
use M2_M1  M2_M1_9974
timestamp 1745462530
transform 1 0 684 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_9975
timestamp 1745462530
transform 1 0 668 0 1 2745
box -2 -2 2 2
use M2_M1  M2_M1_9976
timestamp 1745462530
transform 1 0 644 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_9977
timestamp 1745462530
transform 1 0 716 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_9978
timestamp 1745462530
transform 1 0 692 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_9979
timestamp 1745462530
transform 1 0 2180 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_9980
timestamp 1745462530
transform 1 0 996 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_9981
timestamp 1745462530
transform 1 0 980 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_9982
timestamp 1745462530
transform 1 0 956 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_9983
timestamp 1745462530
transform 1 0 948 0 1 2185
box -2 -2 2 2
use M2_M1  M2_M1_9984
timestamp 1745462530
transform 1 0 940 0 1 2145
box -2 -2 2 2
use M2_M1  M2_M1_9985
timestamp 1745462530
transform 1 0 2180 0 1 2105
box -2 -2 2 2
use M2_M1  M2_M1_9986
timestamp 1745462530
transform 1 0 1092 0 1 1945
box -2 -2 2 2
use M2_M1  M2_M1_9987
timestamp 1745462530
transform 1 0 1092 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_9988
timestamp 1745462530
transform 1 0 1036 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_9989
timestamp 1745462530
transform 1 0 1028 0 1 1195
box -2 -2 2 2
use M2_M1  M2_M1_9990
timestamp 1745462530
transform 1 0 1028 0 1 1145
box -2 -2 2 2
use M2_M1  M2_M1_9991
timestamp 1745462530
transform 1 0 964 0 1 995
box -2 -2 2 2
use M2_M1  M2_M1_9992
timestamp 1745462530
transform 1 0 964 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_9993
timestamp 1745462530
transform 1 0 1548 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_9994
timestamp 1745462530
transform 1 0 1468 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_9995
timestamp 1745462530
transform 1 0 1508 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_9996
timestamp 1745462530
transform 1 0 1484 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_9997
timestamp 1745462530
transform 1 0 1452 0 1 2435
box -2 -2 2 2
use M2_M1  M2_M1_9998
timestamp 1745462530
transform 1 0 1404 0 1 2355
box -2 -2 2 2
use M2_M1  M2_M1_9999
timestamp 1745462530
transform 1 0 1460 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_10000
timestamp 1745462530
transform 1 0 1412 0 1 2345
box -2 -2 2 2
use M2_M1  M2_M1_10001
timestamp 1745462530
transform 1 0 1428 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_10002
timestamp 1745462530
transform 1 0 1364 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_10003
timestamp 1745462530
transform 1 0 2228 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_10004
timestamp 1745462530
transform 1 0 2212 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_10005
timestamp 1745462530
transform 1 0 2188 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_10006
timestamp 1745462530
transform 1 0 2164 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_10007
timestamp 1745462530
transform 1 0 2100 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_10008
timestamp 1745462530
transform 1 0 2100 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_10009
timestamp 1745462530
transform 1 0 2060 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_10010
timestamp 1745462530
transform 1 0 1116 0 1 945
box -2 -2 2 2
use M2_M1  M2_M1_10011
timestamp 1745462530
transform 1 0 772 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_10012
timestamp 1745462530
transform 1 0 1188 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_10013
timestamp 1745462530
transform 1 0 1172 0 1 905
box -2 -2 2 2
use M2_M1  M2_M1_10014
timestamp 1745462530
transform 1 0 1300 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_10015
timestamp 1745462530
transform 1 0 1164 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_10016
timestamp 1745462530
transform 1 0 1236 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_10017
timestamp 1745462530
transform 1 0 1172 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_10018
timestamp 1745462530
transform 1 0 1180 0 1 905
box -2 -2 2 2
use M2_M1  M2_M1_10019
timestamp 1745462530
transform 1 0 1164 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_10020
timestamp 1745462530
transform 1 0 1156 0 1 595
box -2 -2 2 2
use M2_M1  M2_M1_10021
timestamp 1745462530
transform 1 0 1108 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_10022
timestamp 1745462530
transform 1 0 1260 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_10023
timestamp 1745462530
transform 1 0 1196 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_10024
timestamp 1745462530
transform 1 0 2124 0 1 2095
box -2 -2 2 2
use M2_M1  M2_M1_10025
timestamp 1745462530
transform 1 0 1636 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_10026
timestamp 1745462530
transform 1 0 1620 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_10027
timestamp 1745462530
transform 1 0 1572 0 1 995
box -2 -2 2 2
use M2_M1  M2_M1_10028
timestamp 1745462530
transform 1 0 1556 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_10029
timestamp 1745462530
transform 1 0 1396 0 1 1145
box -2 -2 2 2
use M2_M1  M2_M1_10030
timestamp 1745462530
transform 1 0 1380 0 1 1145
box -2 -2 2 2
use M2_M1  M2_M1_10031
timestamp 1745462530
transform 1 0 1220 0 1 1195
box -2 -2 2 2
use M2_M1  M2_M1_10032
timestamp 1745462530
transform 1 0 1164 0 1 1195
box -2 -2 2 2
use M2_M1  M2_M1_10033
timestamp 1745462530
transform 1 0 820 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_10034
timestamp 1745462530
transform 1 0 740 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_10035
timestamp 1745462530
transform 1 0 804 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_10036
timestamp 1745462530
transform 1 0 748 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_10037
timestamp 1745462530
transform 1 0 716 0 1 905
box -2 -2 2 2
use M2_M1  M2_M1_10038
timestamp 1745462530
transform 1 0 540 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_10039
timestamp 1745462530
transform 1 0 500 0 1 945
box -2 -2 2 2
use M2_M1  M2_M1_10040
timestamp 1745462530
transform 1 0 476 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_10041
timestamp 1745462530
transform 1 0 540 0 1 895
box -2 -2 2 2
use M2_M1  M2_M1_10042
timestamp 1745462530
transform 1 0 524 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_10043
timestamp 1745462530
transform 1 0 2284 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_10044
timestamp 1745462530
transform 1 0 2236 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_10045
timestamp 1745462530
transform 1 0 2228 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_10046
timestamp 1745462530
transform 1 0 2204 0 1 2995
box -2 -2 2 2
use M2_M1  M2_M1_10047
timestamp 1745462530
transform 1 0 2204 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_10048
timestamp 1745462530
transform 1 0 2124 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_10049
timestamp 1745462530
transform 1 0 2108 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_10050
timestamp 1745462530
transform 1 0 2076 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_10051
timestamp 1745462530
transform 1 0 2060 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_10052
timestamp 1745462530
transform 1 0 2028 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_10053
timestamp 1745462530
transform 1 0 2028 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_10054
timestamp 1745462530
transform 1 0 2332 0 1 2825
box -2 -2 2 2
use M2_M1  M2_M1_10055
timestamp 1745462530
transform 1 0 2180 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_10056
timestamp 1745462530
transform 1 0 2148 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_10057
timestamp 1745462530
transform 1 0 2148 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_10058
timestamp 1745462530
transform 1 0 2100 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_10059
timestamp 1745462530
transform 1 0 2100 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_10060
timestamp 1745462530
transform 1 0 2044 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_10061
timestamp 1745462530
transform 1 0 2036 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_10062
timestamp 1745462530
transform 1 0 2252 0 1 2915
box -2 -2 2 2
use M2_M1  M2_M1_10063
timestamp 1745462530
transform 1 0 2180 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_10064
timestamp 1745462530
transform 1 0 2172 0 1 2825
box -2 -2 2 2
use M2_M1  M2_M1_10065
timestamp 1745462530
transform 1 0 2132 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_10066
timestamp 1745462530
transform 1 0 2076 0 1 2825
box -2 -2 2 2
use M2_M1  M2_M1_10067
timestamp 1745462530
transform 1 0 2052 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_10068
timestamp 1745462530
transform 1 0 2244 0 1 3025
box -2 -2 2 2
use M2_M1  M2_M1_10069
timestamp 1745462530
transform 1 0 2076 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_10070
timestamp 1745462530
transform 1 0 2124 0 1 2825
box -2 -2 2 2
use M2_M1  M2_M1_10071
timestamp 1745462530
transform 1 0 2116 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_10072
timestamp 1745462530
transform 1 0 1132 0 1 3145
box -2 -2 2 2
use M2_M1  M2_M1_10073
timestamp 1745462530
transform 1 0 1108 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_10074
timestamp 1745462530
transform 1 0 988 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_10075
timestamp 1745462530
transform 1 0 252 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_10076
timestamp 1745462530
transform 1 0 212 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_10077
timestamp 1745462530
transform 1 0 516 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_10078
timestamp 1745462530
transform 1 0 452 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_10079
timestamp 1745462530
transform 1 0 356 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_10080
timestamp 1745462530
transform 1 0 244 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_10081
timestamp 1745462530
transform 1 0 244 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_10082
timestamp 1745462530
transform 1 0 252 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_10083
timestamp 1745462530
transform 1 0 220 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_10084
timestamp 1745462530
transform 1 0 364 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_10085
timestamp 1745462530
transform 1 0 308 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_10086
timestamp 1745462530
transform 1 0 460 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_10087
timestamp 1745462530
transform 1 0 412 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_10088
timestamp 1745462530
transform 1 0 724 0 1 3225
box -2 -2 2 2
use M2_M1  M2_M1_10089
timestamp 1745462530
transform 1 0 692 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_10090
timestamp 1745462530
transform 1 0 580 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_10091
timestamp 1745462530
transform 1 0 564 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_10092
timestamp 1745462530
transform 1 0 1532 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_10093
timestamp 1745462530
transform 1 0 1268 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_10094
timestamp 1745462530
transform 1 0 1100 0 1 3235
box -2 -2 2 2
use M2_M1  M2_M1_10095
timestamp 1745462530
transform 1 0 1316 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_10096
timestamp 1745462530
transform 1 0 1284 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_10097
timestamp 1745462530
transform 1 0 1060 0 1 3515
box -2 -2 2 2
use M2_M1  M2_M1_10098
timestamp 1745462530
transform 1 0 956 0 1 3395
box -2 -2 2 2
use M2_M1  M2_M1_10099
timestamp 1745462530
transform 1 0 1084 0 1 3425
box -2 -2 2 2
use M2_M1  M2_M1_10100
timestamp 1745462530
transform 1 0 964 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_10101
timestamp 1745462530
transform 1 0 1060 0 1 3425
box -2 -2 2 2
use M2_M1  M2_M1_10102
timestamp 1745462530
transform 1 0 1052 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_10103
timestamp 1745462530
transform 1 0 1092 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_10104
timestamp 1745462530
transform 1 0 1068 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_10105
timestamp 1745462530
transform 1 0 1132 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_10106
timestamp 1745462530
transform 1 0 1076 0 1 3435
box -2 -2 2 2
use M2_M1  M2_M1_10107
timestamp 1745462530
transform 1 0 1220 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_10108
timestamp 1745462530
transform 1 0 1044 0 1 3515
box -2 -2 2 2
use M2_M1  M2_M1_10109
timestamp 1745462530
transform 1 0 1100 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_10110
timestamp 1745462530
transform 1 0 1044 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_10111
timestamp 1745462530
transform 1 0 1452 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_10112
timestamp 1745462530
transform 1 0 1396 0 1 3745
box -2 -2 2 2
use M2_M1  M2_M1_10113
timestamp 1745462530
transform 1 0 1516 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_10114
timestamp 1745462530
transform 1 0 1404 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_10115
timestamp 1745462530
transform 1 0 1556 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_10116
timestamp 1745462530
transform 1 0 1492 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_10117
timestamp 1745462530
transform 1 0 1444 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_10118
timestamp 1745462530
transform 1 0 1340 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_10119
timestamp 1745462530
transform 1 0 1276 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_10120
timestamp 1745462530
transform 1 0 1524 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_10121
timestamp 1745462530
transform 1 0 1316 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_10122
timestamp 1745462530
transform 1 0 1300 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_10123
timestamp 1745462530
transform 1 0 1292 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_10124
timestamp 1745462530
transform 1 0 1428 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_10125
timestamp 1745462530
transform 1 0 1364 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_10126
timestamp 1745462530
transform 1 0 1308 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_10127
timestamp 1745462530
transform 1 0 1228 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_10128
timestamp 1745462530
transform 1 0 1492 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_10129
timestamp 1745462530
transform 1 0 1492 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_10130
timestamp 1745462530
transform 1 0 1468 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_10131
timestamp 1745462530
transform 1 0 1412 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_10132
timestamp 1745462530
transform 1 0 1580 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_10133
timestamp 1745462530
transform 1 0 1492 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_10134
timestamp 1745462530
transform 1 0 1436 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_10135
timestamp 1745462530
transform 1 0 1396 0 1 3515
box -2 -2 2 2
use M2_M1  M2_M1_10136
timestamp 1745462530
transform 1 0 1356 0 1 3715
box -2 -2 2 2
use M2_M1  M2_M1_10137
timestamp 1745462530
transform 1 0 1356 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_10138
timestamp 1745462530
transform 1 0 1260 0 1 3745
box -2 -2 2 2
use M2_M1  M2_M1_10139
timestamp 1745462530
transform 1 0 1292 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_10140
timestamp 1745462530
transform 1 0 1268 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_10141
timestamp 1745462530
transform 1 0 1612 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_10142
timestamp 1745462530
transform 1 0 1316 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_10143
timestamp 1745462530
transform 1 0 1292 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_10144
timestamp 1745462530
transform 1 0 1468 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_10145
timestamp 1745462530
transform 1 0 1412 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_10146
timestamp 1745462530
transform 1 0 1516 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_10147
timestamp 1745462530
transform 1 0 1492 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_10148
timestamp 1745462530
transform 1 0 1492 0 1 3345
box -2 -2 2 2
use M2_M1  M2_M1_10149
timestamp 1745462530
transform 1 0 1476 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_10150
timestamp 1745462530
transform 1 0 1204 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_10151
timestamp 1745462530
transform 1 0 1516 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_10152
timestamp 1745462530
transform 1 0 1380 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_10153
timestamp 1745462530
transform 1 0 1364 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_10154
timestamp 1745462530
transform 1 0 1364 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_10155
timestamp 1745462530
transform 1 0 1316 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_10156
timestamp 1745462530
transform 1 0 1436 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_10157
timestamp 1745462530
transform 1 0 1428 0 1 3425
box -2 -2 2 2
use M2_M1  M2_M1_10158
timestamp 1745462530
transform 1 0 1508 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_10159
timestamp 1745462530
transform 1 0 1476 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_10160
timestamp 1745462530
transform 1 0 1484 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_10161
timestamp 1745462530
transform 1 0 1420 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_10162
timestamp 1745462530
transform 1 0 1500 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_10163
timestamp 1745462530
transform 1 0 1396 0 1 3345
box -2 -2 2 2
use M2_M1  M2_M1_10164
timestamp 1745462530
transform 1 0 1332 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_10165
timestamp 1745462530
transform 1 0 1564 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_10166
timestamp 1745462530
transform 1 0 1420 0 1 3425
box -2 -2 2 2
use M2_M1  M2_M1_10167
timestamp 1745462530
transform 1 0 1628 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_10168
timestamp 1745462530
transform 1 0 1580 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_10169
timestamp 1745462530
transform 1 0 996 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_10170
timestamp 1745462530
transform 1 0 916 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_10171
timestamp 1745462530
transform 1 0 1156 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_10172
timestamp 1745462530
transform 1 0 1044 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_10173
timestamp 1745462530
transform 1 0 836 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_10174
timestamp 1745462530
transform 1 0 780 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_10175
timestamp 1745462530
transform 1 0 3132 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_10176
timestamp 1745462530
transform 1 0 3068 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_10177
timestamp 1745462530
transform 1 0 3380 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_10178
timestamp 1745462530
transform 1 0 3380 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_10179
timestamp 1745462530
transform 1 0 3308 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_10180
timestamp 1745462530
transform 1 0 3292 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_10181
timestamp 1745462530
transform 1 0 3364 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_10182
timestamp 1745462530
transform 1 0 3300 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_10183
timestamp 1745462530
transform 1 0 3172 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_10184
timestamp 1745462530
transform 1 0 3172 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_10185
timestamp 1745462530
transform 1 0 2484 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_10186
timestamp 1745462530
transform 1 0 2396 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_10187
timestamp 1745462530
transform 1 0 2092 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_10188
timestamp 1745462530
transform 1 0 2084 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_10189
timestamp 1745462530
transform 1 0 2852 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_10190
timestamp 1745462530
transform 1 0 2772 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_10191
timestamp 1745462530
transform 1 0 3108 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_10192
timestamp 1745462530
transform 1 0 3100 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_10193
timestamp 1745462530
transform 1 0 3868 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_10194
timestamp 1745462530
transform 1 0 3644 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_10195
timestamp 1745462530
transform 1 0 3684 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_10196
timestamp 1745462530
transform 1 0 3612 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_10197
timestamp 1745462530
transform 1 0 3756 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_10198
timestamp 1745462530
transform 1 0 3604 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_10199
timestamp 1745462530
transform 1 0 3316 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_10200
timestamp 1745462530
transform 1 0 3244 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_10201
timestamp 1745462530
transform 1 0 2484 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_10202
timestamp 1745462530
transform 1 0 2388 0 1 4005
box -2 -2 2 2
use M2_M1  M2_M1_10203
timestamp 1745462530
transform 1 0 2276 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_10204
timestamp 1745462530
transform 1 0 2228 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_10205
timestamp 1745462530
transform 1 0 2836 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_10206
timestamp 1745462530
transform 1 0 2756 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_10207
timestamp 1745462530
transform 1 0 3124 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_10208
timestamp 1745462530
transform 1 0 3028 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_10209
timestamp 1745462530
transform 1 0 3564 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_10210
timestamp 1745462530
transform 1 0 3500 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_10211
timestamp 1745462530
transform 1 0 3412 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_10212
timestamp 1745462530
transform 1 0 3396 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_10213
timestamp 1745462530
transform 1 0 3660 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_10214
timestamp 1745462530
transform 1 0 3516 0 1 4005
box -2 -2 2 2
use M2_M1  M2_M1_10215
timestamp 1745462530
transform 1 0 3220 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_10216
timestamp 1745462530
transform 1 0 3188 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_10217
timestamp 1745462530
transform 1 0 2420 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_10218
timestamp 1745462530
transform 1 0 2396 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_10219
timestamp 1745462530
transform 1 0 2188 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_10220
timestamp 1745462530
transform 1 0 2084 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_10221
timestamp 1745462530
transform 1 0 2756 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_10222
timestamp 1745462530
transform 1 0 2660 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_10223
timestamp 1745462530
transform 1 0 2996 0 1 4005
box -2 -2 2 2
use M2_M1  M2_M1_10224
timestamp 1745462530
transform 1 0 2956 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_10225
timestamp 1745462530
transform 1 0 3868 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_10226
timestamp 1745462530
transform 1 0 3772 0 1 4005
box -2 -2 2 2
use M2_M1  M2_M1_10227
timestamp 1745462530
transform 1 0 3948 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_10228
timestamp 1745462530
transform 1 0 3868 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_10229
timestamp 1745462530
transform 1 0 3788 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_10230
timestamp 1745462530
transform 1 0 3700 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_10231
timestamp 1745462530
transform 1 0 3756 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_10232
timestamp 1745462530
transform 1 0 3724 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_10233
timestamp 1745462530
transform 1 0 2500 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_10234
timestamp 1745462530
transform 1 0 2492 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_10235
timestamp 1745462530
transform 1 0 2300 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_10236
timestamp 1745462530
transform 1 0 2260 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_10237
timestamp 1745462530
transform 1 0 2604 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_10238
timestamp 1745462530
transform 1 0 2604 0 1 4005
box -2 -2 2 2
use M2_M1  M2_M1_10239
timestamp 1745462530
transform 1 0 2932 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_10240
timestamp 1745462530
transform 1 0 2916 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_10241
timestamp 1745462530
transform 1 0 4316 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_10242
timestamp 1745462530
transform 1 0 4316 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_10243
timestamp 1745462530
transform 1 0 4308 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_10244
timestamp 1745462530
transform 1 0 4228 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_10245
timestamp 1745462530
transform 1 0 4316 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_10246
timestamp 1745462530
transform 1 0 4244 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_10247
timestamp 1745462530
transform 1 0 3972 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_10248
timestamp 1745462530
transform 1 0 3972 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_10249
timestamp 1745462530
transform 1 0 1996 0 1 3736
box -2 -2 2 2
use M2_M1  M2_M1_10250
timestamp 1745462530
transform 1 0 1948 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_10251
timestamp 1745462530
transform 1 0 2028 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_10252
timestamp 1745462530
transform 1 0 2020 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_10253
timestamp 1745462530
transform 1 0 2692 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_10254
timestamp 1745462530
transform 1 0 2628 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_10255
timestamp 1745462530
transform 1 0 2940 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_10256
timestamp 1745462530
transform 1 0 2868 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_10257
timestamp 1745462530
transform 1 0 4188 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_10258
timestamp 1745462530
transform 1 0 4084 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_10259
timestamp 1745462530
transform 1 0 4140 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_10260
timestamp 1745462530
transform 1 0 4060 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_10261
timestamp 1745462530
transform 1 0 4308 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_10262
timestamp 1745462530
transform 1 0 4148 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_10263
timestamp 1745462530
transform 1 0 4076 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_10264
timestamp 1745462530
transform 1 0 3980 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_10265
timestamp 1745462530
transform 1 0 2028 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_10266
timestamp 1745462530
transform 1 0 1964 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_10267
timestamp 1745462530
transform 1 0 1980 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_10268
timestamp 1745462530
transform 1 0 1940 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_10269
timestamp 1745462530
transform 1 0 1876 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_10270
timestamp 1745462530
transform 1 0 1876 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_10271
timestamp 1745462530
transform 1 0 1796 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_10272
timestamp 1745462530
transform 1 0 1796 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_10273
timestamp 1745462530
transform 1 0 4316 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_10274
timestamp 1745462530
transform 1 0 4236 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_10275
timestamp 1745462530
transform 1 0 4316 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_10276
timestamp 1745462530
transform 1 0 4228 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_10277
timestamp 1745462530
transform 1 0 4124 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_10278
timestamp 1745462530
transform 1 0 4044 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_10279
timestamp 1745462530
transform 1 0 3964 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_10280
timestamp 1745462530
transform 1 0 3964 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_10281
timestamp 1745462530
transform 1 0 1676 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_10282
timestamp 1745462530
transform 1 0 1564 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_10283
timestamp 1745462530
transform 1 0 1660 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_10284
timestamp 1745462530
transform 1 0 1436 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_10285
timestamp 1745462530
transform 1 0 1724 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_10286
timestamp 1745462530
transform 1 0 1668 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_10287
timestamp 1745462530
transform 1 0 1700 0 1 4005
box -2 -2 2 2
use M2_M1  M2_M1_10288
timestamp 1745462530
transform 1 0 1548 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_10289
timestamp 1745462530
transform 1 0 4308 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_10290
timestamp 1745462530
transform 1 0 4220 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_10291
timestamp 1745462530
transform 1 0 4308 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_10292
timestamp 1745462530
transform 1 0 4228 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_10293
timestamp 1745462530
transform 1 0 4140 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_10294
timestamp 1745462530
transform 1 0 4044 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_10295
timestamp 1745462530
transform 1 0 3932 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_10296
timestamp 1745462530
transform 1 0 3836 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_10297
timestamp 1745462530
transform 1 0 1572 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_10298
timestamp 1745462530
transform 1 0 1508 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_10299
timestamp 1745462530
transform 1 0 2812 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_10300
timestamp 1745462530
transform 1 0 2796 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_10301
timestamp 1745462530
transform 1 0 1604 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_10302
timestamp 1745462530
transform 1 0 1396 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_10303
timestamp 1745462530
transform 1 0 836 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_10304
timestamp 1745462530
transform 1 0 740 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_10305
timestamp 1745462530
transform 1 0 876 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_10306
timestamp 1745462530
transform 1 0 812 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_10307
timestamp 1745462530
transform 1 0 1020 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_10308
timestamp 1745462530
transform 1 0 948 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_10309
timestamp 1745462530
transform 1 0 860 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_10310
timestamp 1745462530
transform 1 0 764 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_10311
timestamp 1745462530
transform 1 0 1276 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_10312
timestamp 1745462530
transform 1 0 1196 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_10313
timestamp 1745462530
transform 1 0 1452 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_10314
timestamp 1745462530
transform 1 0 1452 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_10315
timestamp 1745462530
transform 1 0 1580 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_10316
timestamp 1745462530
transform 1 0 1516 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_10317
timestamp 1745462530
transform 1 0 1428 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_10318
timestamp 1745462530
transform 1 0 1380 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_10319
timestamp 1745462530
transform 1 0 1940 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_10320
timestamp 1745462530
transform 1 0 1628 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_10321
timestamp 1745462530
transform 1 0 1068 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_10322
timestamp 1745462530
transform 1 0 1060 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_10323
timestamp 1745462530
transform 1 0 1964 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_10324
timestamp 1745462530
transform 1 0 1892 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_10325
timestamp 1745462530
transform 1 0 2076 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_10326
timestamp 1745462530
transform 1 0 1988 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_10327
timestamp 1745462530
transform 1 0 2052 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_10328
timestamp 1745462530
transform 1 0 1908 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_10329
timestamp 1745462530
transform 1 0 2108 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_10330
timestamp 1745462530
transform 1 0 1804 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_10331
timestamp 1745462530
transform 1 0 1788 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_10332
timestamp 1745462530
transform 1 0 1772 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_10333
timestamp 1745462530
transform 1 0 1772 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_10334
timestamp 1745462530
transform 1 0 1732 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_10335
timestamp 1745462530
transform 1 0 380 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_10336
timestamp 1745462530
transform 1 0 308 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_10337
timestamp 1745462530
transform 1 0 588 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_10338
timestamp 1745462530
transform 1 0 548 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_10339
timestamp 1745462530
transform 1 0 220 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_10340
timestamp 1745462530
transform 1 0 140 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_10341
timestamp 1745462530
transform 1 0 972 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_10342
timestamp 1745462530
transform 1 0 956 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_10343
timestamp 1745462530
transform 1 0 308 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_10344
timestamp 1745462530
transform 1 0 284 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_10345
timestamp 1745462530
transform 1 0 292 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_10346
timestamp 1745462530
transform 1 0 260 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_10347
timestamp 1745462530
transform 1 0 284 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_10348
timestamp 1745462530
transform 1 0 268 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_10349
timestamp 1745462530
transform 1 0 620 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_10350
timestamp 1745462530
transform 1 0 580 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_10351
timestamp 1745462530
transform 1 0 356 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_10352
timestamp 1745462530
transform 1 0 252 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_10353
timestamp 1745462530
transform 1 0 252 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_10354
timestamp 1745462530
transform 1 0 148 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_10355
timestamp 1745462530
transform 1 0 260 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_10356
timestamp 1745462530
transform 1 0 188 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_10357
timestamp 1745462530
transform 1 0 596 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_10358
timestamp 1745462530
transform 1 0 476 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_10359
timestamp 1745462530
transform 1 0 716 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_10360
timestamp 1745462530
transform 1 0 620 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_10361
timestamp 1745462530
transform 1 0 852 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_10362
timestamp 1745462530
transform 1 0 780 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_10363
timestamp 1745462530
transform 1 0 580 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_10364
timestamp 1745462530
transform 1 0 492 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_10365
timestamp 1745462530
transform 1 0 724 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_10366
timestamp 1745462530
transform 1 0 692 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_10367
timestamp 1745462530
transform 1 0 1500 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_10368
timestamp 1745462530
transform 1 0 1404 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_10369
timestamp 1745462530
transform 1 0 1772 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_10370
timestamp 1745462530
transform 1 0 1684 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_10371
timestamp 1745462530
transform 1 0 1668 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_10372
timestamp 1745462530
transform 1 0 1572 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_10373
timestamp 1745462530
transform 1 0 1740 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_10374
timestamp 1745462530
transform 1 0 1716 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_10375
timestamp 1745462530
transform 1 0 1740 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_10376
timestamp 1745462530
transform 1 0 1732 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_10377
timestamp 1745462530
transform 1 0 1796 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_10378
timestamp 1745462530
transform 1 0 1796 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_10379
timestamp 1745462530
transform 1 0 1844 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_10380
timestamp 1745462530
transform 1 0 1756 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_10381
timestamp 1745462530
transform 1 0 1844 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_10382
timestamp 1745462530
transform 1 0 1764 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_10383
timestamp 1745462530
transform 1 0 2932 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_10384
timestamp 1745462530
transform 1 0 2908 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_10385
timestamp 1745462530
transform 1 0 3124 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_10386
timestamp 1745462530
transform 1 0 3036 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_10387
timestamp 1745462530
transform 1 0 2820 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_10388
timestamp 1745462530
transform 1 0 2820 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_10389
timestamp 1745462530
transform 1 0 3028 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_10390
timestamp 1745462530
transform 1 0 2940 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_10391
timestamp 1745462530
transform 1 0 3148 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_10392
timestamp 1745462530
transform 1 0 3116 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_10393
timestamp 1745462530
transform 1 0 2988 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_10394
timestamp 1745462530
transform 1 0 2916 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_10395
timestamp 1745462530
transform 1 0 3028 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_10396
timestamp 1745462530
transform 1 0 2860 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_10397
timestamp 1745462530
transform 1 0 2916 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_10398
timestamp 1745462530
transform 1 0 2812 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_10399
timestamp 1745462530
transform 1 0 3372 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_10400
timestamp 1745462530
transform 1 0 3316 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_10401
timestamp 1745462530
transform 1 0 3940 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_10402
timestamp 1745462530
transform 1 0 3892 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_10403
timestamp 1745462530
transform 1 0 4164 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_10404
timestamp 1745462530
transform 1 0 4156 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_10405
timestamp 1745462530
transform 1 0 4060 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_10406
timestamp 1745462530
transform 1 0 3996 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_10407
timestamp 1745462530
transform 1 0 4188 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_10408
timestamp 1745462530
transform 1 0 4164 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_10409
timestamp 1745462530
transform 1 0 4316 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_10410
timestamp 1745462530
transform 1 0 4316 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_10411
timestamp 1745462530
transform 1 0 4220 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_10412
timestamp 1745462530
transform 1 0 4140 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_10413
timestamp 1745462530
transform 1 0 4116 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_10414
timestamp 1745462530
transform 1 0 3884 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_10415
timestamp 1745462530
transform 1 0 4188 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_10416
timestamp 1745462530
transform 1 0 4116 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_10417
timestamp 1745462530
transform 1 0 3988 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_10418
timestamp 1745462530
transform 1 0 3836 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_10419
timestamp 1745462530
transform 1 0 4324 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_10420
timestamp 1745462530
transform 1 0 4188 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_10421
timestamp 1745462530
transform 1 0 4036 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_10422
timestamp 1745462530
transform 1 0 3860 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_10423
timestamp 1745462530
transform 1 0 4228 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_10424
timestamp 1745462530
transform 1 0 4228 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_10425
timestamp 1745462530
transform 1 0 3980 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_10426
timestamp 1745462530
transform 1 0 3860 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_10427
timestamp 1745462530
transform 1 0 3220 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_10428
timestamp 1745462530
transform 1 0 3124 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_10429
timestamp 1745462530
transform 1 0 3028 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_10430
timestamp 1745462530
transform 1 0 2940 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_10431
timestamp 1745462530
transform 1 0 4268 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_10432
timestamp 1745462530
transform 1 0 4196 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_10433
timestamp 1745462530
transform 1 0 4020 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_10434
timestamp 1745462530
transform 1 0 3924 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_10435
timestamp 1745462530
transform 1 0 4212 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_10436
timestamp 1745462530
transform 1 0 4092 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_10437
timestamp 1745462530
transform 1 0 4276 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_10438
timestamp 1745462530
transform 1 0 4180 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_10439
timestamp 1745462530
transform 1 0 4308 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_10440
timestamp 1745462530
transform 1 0 4220 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_10441
timestamp 1745462530
transform 1 0 4316 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_10442
timestamp 1745462530
transform 1 0 4236 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_10443
timestamp 1745462530
transform 1 0 4108 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_10444
timestamp 1745462530
transform 1 0 4108 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_10445
timestamp 1745462530
transform 1 0 2916 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_10446
timestamp 1745462530
transform 1 0 2884 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_10447
timestamp 1745462530
transform 1 0 2812 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_10448
timestamp 1745462530
transform 1 0 2780 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_10449
timestamp 1745462530
transform 1 0 1372 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_10450
timestamp 1745462530
transform 1 0 1308 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_10451
timestamp 1745462530
transform 1 0 1308 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_10452
timestamp 1745462530
transform 1 0 1300 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_10453
timestamp 1745462530
transform 1 0 1284 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_10454
timestamp 1745462530
transform 1 0 1260 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_10455
timestamp 1745462530
transform 1 0 1340 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_10456
timestamp 1745462530
transform 1 0 1236 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_10457
timestamp 1745462530
transform 1 0 1252 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_10458
timestamp 1745462530
transform 1 0 1244 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_10459
timestamp 1745462530
transform 1 0 1260 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_10460
timestamp 1745462530
transform 1 0 1244 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_10461
timestamp 1745462530
transform 1 0 396 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_10462
timestamp 1745462530
transform 1 0 380 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_10463
timestamp 1745462530
transform 1 0 588 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_10464
timestamp 1745462530
transform 1 0 540 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_10465
timestamp 1745462530
transform 1 0 300 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_10466
timestamp 1745462530
transform 1 0 236 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_10467
timestamp 1745462530
transform 1 0 1148 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_10468
timestamp 1745462530
transform 1 0 964 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_10469
timestamp 1745462530
transform 1 0 444 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_10470
timestamp 1745462530
transform 1 0 404 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_10471
timestamp 1745462530
transform 1 0 500 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_10472
timestamp 1745462530
transform 1 0 428 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_10473
timestamp 1745462530
transform 1 0 428 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_10474
timestamp 1745462530
transform 1 0 396 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_10475
timestamp 1745462530
transform 1 0 828 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_10476
timestamp 1745462530
transform 1 0 724 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_10477
timestamp 1745462530
transform 1 0 492 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_10478
timestamp 1745462530
transform 1 0 484 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_10479
timestamp 1745462530
transform 1 0 500 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_10480
timestamp 1745462530
transform 1 0 388 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_10481
timestamp 1745462530
transform 1 0 332 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_10482
timestamp 1745462530
transform 1 0 332 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_10483
timestamp 1745462530
transform 1 0 412 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_10484
timestamp 1745462530
transform 1 0 412 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_10485
timestamp 1745462530
transform 1 0 716 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_10486
timestamp 1745462530
transform 1 0 644 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_10487
timestamp 1745462530
transform 1 0 948 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_10488
timestamp 1745462530
transform 1 0 908 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_10489
timestamp 1745462530
transform 1 0 476 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_10490
timestamp 1745462530
transform 1 0 388 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_10491
timestamp 1745462530
transform 1 0 708 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_10492
timestamp 1745462530
transform 1 0 620 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_10493
timestamp 1745462530
transform 1 0 1172 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_10494
timestamp 1745462530
transform 1 0 1084 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_10495
timestamp 1745462530
transform 1 0 1532 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_10496
timestamp 1745462530
transform 1 0 1436 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_10497
timestamp 1745462530
transform 1 0 1460 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_10498
timestamp 1745462530
transform 1 0 1420 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_10499
timestamp 1745462530
transform 1 0 1428 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_10500
timestamp 1745462530
transform 1 0 1332 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_10501
timestamp 1745462530
transform 1 0 1596 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_10502
timestamp 1745462530
transform 1 0 1500 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_10503
timestamp 1745462530
transform 1 0 1604 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_10504
timestamp 1745462530
transform 1 0 1572 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_10505
timestamp 1745462530
transform 1 0 1596 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_10506
timestamp 1745462530
transform 1 0 1596 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_10507
timestamp 1745462530
transform 1 0 1668 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_10508
timestamp 1745462530
transform 1 0 1604 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_10509
timestamp 1745462530
transform 1 0 2876 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_10510
timestamp 1745462530
transform 1 0 2852 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_10511
timestamp 1745462530
transform 1 0 3188 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_10512
timestamp 1745462530
transform 1 0 3084 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_10513
timestamp 1745462530
transform 1 0 2748 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_10514
timestamp 1745462530
transform 1 0 2676 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_10515
timestamp 1745462530
transform 1 0 3108 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_10516
timestamp 1745462530
transform 1 0 3012 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_10517
timestamp 1745462530
transform 1 0 3060 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_10518
timestamp 1745462530
transform 1 0 2972 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_10519
timestamp 1745462530
transform 1 0 2940 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_10520
timestamp 1745462530
transform 1 0 2908 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_10521
timestamp 1745462530
transform 1 0 2916 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_10522
timestamp 1745462530
transform 1 0 2844 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_10523
timestamp 1745462530
transform 1 0 2948 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_10524
timestamp 1745462530
transform 1 0 2852 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_10525
timestamp 1745462530
transform 1 0 3276 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_10526
timestamp 1745462530
transform 1 0 3188 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_10527
timestamp 1745462530
transform 1 0 3364 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_10528
timestamp 1745462530
transform 1 0 3164 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_10529
timestamp 1745462530
transform 1 0 4140 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_10530
timestamp 1745462530
transform 1 0 4084 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_10531
timestamp 1745462530
transform 1 0 3380 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_10532
timestamp 1745462530
transform 1 0 3380 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_10533
timestamp 1745462530
transform 1 0 4228 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_10534
timestamp 1745462530
transform 1 0 4156 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_10535
timestamp 1745462530
transform 1 0 4068 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_10536
timestamp 1745462530
transform 1 0 4036 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_10537
timestamp 1745462530
transform 1 0 3396 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_10538
timestamp 1745462530
transform 1 0 3308 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_10539
timestamp 1745462530
transform 1 0 3380 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_10540
timestamp 1745462530
transform 1 0 3276 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_10541
timestamp 1745462530
transform 1 0 4100 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_10542
timestamp 1745462530
transform 1 0 4092 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_10543
timestamp 1745462530
transform 1 0 3540 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_10544
timestamp 1745462530
transform 1 0 3516 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_10545
timestamp 1745462530
transform 1 0 4140 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_10546
timestamp 1745462530
transform 1 0 4076 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_10547
timestamp 1745462530
transform 1 0 3580 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_10548
timestamp 1745462530
transform 1 0 3500 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_10549
timestamp 1745462530
transform 1 0 4252 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_10550
timestamp 1745462530
transform 1 0 4172 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_10551
timestamp 1745462530
transform 1 0 3292 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_10552
timestamp 1745462530
transform 1 0 3292 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_10553
timestamp 1745462530
transform 1 0 2828 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_10554
timestamp 1745462530
transform 1 0 2780 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_10555
timestamp 1745462530
transform 1 0 2780 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_10556
timestamp 1745462530
transform 1 0 2780 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_10557
timestamp 1745462530
transform 1 0 3284 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_10558
timestamp 1745462530
transform 1 0 3212 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_10559
timestamp 1745462530
transform 1 0 3012 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_10560
timestamp 1745462530
transform 1 0 2932 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_10561
timestamp 1745462530
transform 1 0 3260 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_10562
timestamp 1745462530
transform 1 0 3116 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_10563
timestamp 1745462530
transform 1 0 3212 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_10564
timestamp 1745462530
transform 1 0 3132 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_10565
timestamp 1745462530
transform 1 0 3292 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_10566
timestamp 1745462530
transform 1 0 3292 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_10567
timestamp 1745462530
transform 1 0 3252 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_10568
timestamp 1745462530
transform 1 0 3180 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_10569
timestamp 1745462530
transform 1 0 3188 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_10570
timestamp 1745462530
transform 1 0 3108 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_10571
timestamp 1745462530
transform 1 0 2764 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_10572
timestamp 1745462530
transform 1 0 2732 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_10573
timestamp 1745462530
transform 1 0 2804 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_10574
timestamp 1745462530
transform 1 0 2732 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_10575
timestamp 1745462530
transform 1 0 1756 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_10576
timestamp 1745462530
transform 1 0 1756 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_10577
timestamp 1745462530
transform 1 0 1708 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_10578
timestamp 1745462530
transform 1 0 1692 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_10579
timestamp 1745462530
transform 1 0 1748 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_10580
timestamp 1745462530
transform 1 0 1692 0 1 2737
box -2 -2 2 2
use M2_M1  M2_M1_10581
timestamp 1745462530
transform 1 0 1700 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_10582
timestamp 1745462530
transform 1 0 1596 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_10583
timestamp 1745462530
transform 1 0 1644 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_10584
timestamp 1745462530
transform 1 0 1532 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_10585
timestamp 1745462530
transform 1 0 1572 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_10586
timestamp 1745462530
transform 1 0 1572 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_10587
timestamp 1745462530
transform 1 0 436 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_10588
timestamp 1745462530
transform 1 0 356 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_10589
timestamp 1745462530
transform 1 0 524 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_10590
timestamp 1745462530
transform 1 0 452 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_10591
timestamp 1745462530
transform 1 0 348 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_10592
timestamp 1745462530
transform 1 0 260 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_10593
timestamp 1745462530
transform 1 0 1060 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_10594
timestamp 1745462530
transform 1 0 964 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_10595
timestamp 1745462530
transform 1 0 452 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_10596
timestamp 1745462530
transform 1 0 364 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_10597
timestamp 1745462530
transform 1 0 476 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_10598
timestamp 1745462530
transform 1 0 444 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_10599
timestamp 1745462530
transform 1 0 460 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_10600
timestamp 1745462530
transform 1 0 436 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_10601
timestamp 1745462530
transform 1 0 580 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_10602
timestamp 1745462530
transform 1 0 580 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_10603
timestamp 1745462530
transform 1 0 428 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_10604
timestamp 1745462530
transform 1 0 380 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_10605
timestamp 1745462530
transform 1 0 380 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_10606
timestamp 1745462530
transform 1 0 316 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_10607
timestamp 1745462530
transform 1 0 260 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_10608
timestamp 1745462530
transform 1 0 220 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_10609
timestamp 1745462530
transform 1 0 332 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_10610
timestamp 1745462530
transform 1 0 316 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_10611
timestamp 1745462530
transform 1 0 548 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_10612
timestamp 1745462530
transform 1 0 476 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_10613
timestamp 1745462530
transform 1 0 844 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_10614
timestamp 1745462530
transform 1 0 844 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_10615
timestamp 1745462530
transform 1 0 324 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_10616
timestamp 1745462530
transform 1 0 308 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_10617
timestamp 1745462530
transform 1 0 772 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_10618
timestamp 1745462530
transform 1 0 708 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_10619
timestamp 1745462530
transform 1 0 1700 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_10620
timestamp 1745462530
transform 1 0 1700 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_10621
timestamp 1745462530
transform 1 0 1844 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_10622
timestamp 1745462530
transform 1 0 1828 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_10623
timestamp 1745462530
transform 1 0 1812 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_10624
timestamp 1745462530
transform 1 0 1804 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_10625
timestamp 1745462530
transform 1 0 1852 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_10626
timestamp 1745462530
transform 1 0 1836 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_10627
timestamp 1745462530
transform 1 0 2004 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_10628
timestamp 1745462530
transform 1 0 1908 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_10629
timestamp 1745462530
transform 1 0 2036 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_10630
timestamp 1745462530
transform 1 0 1948 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_10631
timestamp 1745462530
transform 1 0 2004 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_10632
timestamp 1745462530
transform 1 0 1940 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_10633
timestamp 1745462530
transform 1 0 1940 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_10634
timestamp 1745462530
transform 1 0 1916 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_10635
timestamp 1745462530
transform 1 0 2244 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_10636
timestamp 1745462530
transform 1 0 2132 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_10637
timestamp 1745462530
transform 1 0 2204 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_10638
timestamp 1745462530
transform 1 0 2116 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_10639
timestamp 1745462530
transform 1 0 2252 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_10640
timestamp 1745462530
transform 1 0 2236 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_10641
timestamp 1745462530
transform 1 0 2244 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_10642
timestamp 1745462530
transform 1 0 2148 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_10643
timestamp 1745462530
transform 1 0 2508 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_10644
timestamp 1745462530
transform 1 0 2404 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_10645
timestamp 1745462530
transform 1 0 2356 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_10646
timestamp 1745462530
transform 1 0 2220 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_10647
timestamp 1745462530
transform 1 0 2308 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_10648
timestamp 1745462530
transform 1 0 2236 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_10649
timestamp 1745462530
transform 1 0 2380 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_10650
timestamp 1745462530
transform 1 0 2268 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_10651
timestamp 1745462530
transform 1 0 3484 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_10652
timestamp 1745462530
transform 1 0 3444 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_10653
timestamp 1745462530
transform 1 0 3828 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_10654
timestamp 1745462530
transform 1 0 3820 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_10655
timestamp 1745462530
transform 1 0 4300 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_10656
timestamp 1745462530
transform 1 0 4228 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_10657
timestamp 1745462530
transform 1 0 4076 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_10658
timestamp 1745462530
transform 1 0 3996 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_10659
timestamp 1745462530
transform 1 0 4316 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_10660
timestamp 1745462530
transform 1 0 4316 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_10661
timestamp 1745462530
transform 1 0 4316 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_10662
timestamp 1745462530
transform 1 0 4252 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_10663
timestamp 1745462530
transform 1 0 4316 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_10664
timestamp 1745462530
transform 1 0 4228 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_10665
timestamp 1745462530
transform 1 0 4028 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_10666
timestamp 1745462530
transform 1 0 3932 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_10667
timestamp 1745462530
transform 1 0 4308 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_10668
timestamp 1745462530
transform 1 0 4220 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_10669
timestamp 1745462530
transform 1 0 3684 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_10670
timestamp 1745462530
transform 1 0 3676 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_10671
timestamp 1745462530
transform 1 0 4316 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_10672
timestamp 1745462530
transform 1 0 4228 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_10673
timestamp 1745462530
transform 1 0 3660 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_10674
timestamp 1745462530
transform 1 0 3636 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_10675
timestamp 1745462530
transform 1 0 4324 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_10676
timestamp 1745462530
transform 1 0 4316 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_10677
timestamp 1745462530
transform 1 0 3316 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_10678
timestamp 1745462530
transform 1 0 3284 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_10679
timestamp 1745462530
transform 1 0 2876 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_10680
timestamp 1745462530
transform 1 0 2876 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_10681
timestamp 1745462530
transform 1 0 2676 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_10682
timestamp 1745462530
transform 1 0 2596 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_10683
timestamp 1745462530
transform 1 0 4276 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_10684
timestamp 1745462530
transform 1 0 4204 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_10685
timestamp 1745462530
transform 1 0 3988 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_10686
timestamp 1745462530
transform 1 0 3908 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_10687
timestamp 1745462530
transform 1 0 4316 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_10688
timestamp 1745462530
transform 1 0 4156 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_10689
timestamp 1745462530
transform 1 0 4316 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_10690
timestamp 1745462530
transform 1 0 4236 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_10691
timestamp 1745462530
transform 1 0 4300 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_10692
timestamp 1745462530
transform 1 0 4228 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_10693
timestamp 1745462530
transform 1 0 4188 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_10694
timestamp 1745462530
transform 1 0 4188 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_10695
timestamp 1745462530
transform 1 0 4140 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_10696
timestamp 1745462530
transform 1 0 4068 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_10697
timestamp 1745462530
transform 1 0 2836 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_10698
timestamp 1745462530
transform 1 0 2828 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_10699
timestamp 1745462530
transform 1 0 2620 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_10700
timestamp 1745462530
transform 1 0 2556 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_10701
timestamp 1745462530
transform 1 0 1844 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_10702
timestamp 1745462530
transform 1 0 1820 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_10703
timestamp 1745462530
transform 1 0 1940 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_10704
timestamp 1745462530
transform 1 0 1908 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_10705
timestamp 1745462530
transform 1 0 1900 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_10706
timestamp 1745462530
transform 1 0 1836 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_10707
timestamp 1745462530
transform 1 0 2012 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_10708
timestamp 1745462530
transform 1 0 1844 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_10709
timestamp 1745462530
transform 1 0 1740 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_10710
timestamp 1745462530
transform 1 0 1724 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_10711
timestamp 1745462530
transform 1 0 1908 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_10712
timestamp 1745462530
transform 1 0 1804 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_10713
timestamp 1745462530
transform 1 0 780 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_10714
timestamp 1745462530
transform 1 0 764 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_10715
timestamp 1745462530
transform 1 0 692 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_10716
timestamp 1745462530
transform 1 0 692 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_10717
timestamp 1745462530
transform 1 0 468 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_10718
timestamp 1745462530
transform 1 0 452 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_10719
timestamp 1745462530
transform 1 0 1036 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_10720
timestamp 1745462530
transform 1 0 916 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_10721
timestamp 1745462530
transform 1 0 380 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_10722
timestamp 1745462530
transform 1 0 332 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_10723
timestamp 1745462530
transform 1 0 364 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_10724
timestamp 1745462530
transform 1 0 300 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_10725
timestamp 1745462530
transform 1 0 348 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_10726
timestamp 1745462530
transform 1 0 348 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_10727
timestamp 1745462530
transform 1 0 788 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_10728
timestamp 1745462530
transform 1 0 668 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_10729
timestamp 1745462530
transform 1 0 364 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_10730
timestamp 1745462530
transform 1 0 260 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_10731
timestamp 1745462530
transform 1 0 212 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_10732
timestamp 1745462530
transform 1 0 140 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_10733
timestamp 1745462530
transform 1 0 212 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_10734
timestamp 1745462530
transform 1 0 148 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_10735
timestamp 1745462530
transform 1 0 220 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_10736
timestamp 1745462530
transform 1 0 148 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_10737
timestamp 1745462530
transform 1 0 812 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_10738
timestamp 1745462530
transform 1 0 716 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_10739
timestamp 1745462530
transform 1 0 916 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_10740
timestamp 1745462530
transform 1 0 908 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_10741
timestamp 1745462530
transform 1 0 204 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_10742
timestamp 1745462530
transform 1 0 164 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_10743
timestamp 1745462530
transform 1 0 852 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_10744
timestamp 1745462530
transform 1 0 852 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_10745
timestamp 1745462530
transform 1 0 1636 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_10746
timestamp 1745462530
transform 1 0 1620 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_10747
timestamp 1745462530
transform 1 0 2020 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_10748
timestamp 1745462530
transform 1 0 1932 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_10749
timestamp 1745462530
transform 1 0 2004 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_10750
timestamp 1745462530
transform 1 0 1900 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_10751
timestamp 1745462530
transform 1 0 2020 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_10752
timestamp 1745462530
transform 1 0 1900 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_10753
timestamp 1745462530
transform 1 0 2012 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_10754
timestamp 1745462530
transform 1 0 1908 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_10755
timestamp 1745462530
transform 1 0 2084 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_10756
timestamp 1745462530
transform 1 0 2012 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_10757
timestamp 1745462530
transform 1 0 2180 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_10758
timestamp 1745462530
transform 1 0 2012 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_10759
timestamp 1745462530
transform 1 0 2116 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_10760
timestamp 1745462530
transform 1 0 2004 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_10761
timestamp 1745462530
transform 1 0 2380 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_10762
timestamp 1745462530
transform 1 0 2372 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_10763
timestamp 1745462530
transform 1 0 2364 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_10764
timestamp 1745462530
transform 1 0 2292 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_10765
timestamp 1745462530
transform 1 0 2524 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_10766
timestamp 1745462530
transform 1 0 2516 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_10767
timestamp 1745462530
transform 1 0 2380 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_10768
timestamp 1745462530
transform 1 0 2308 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_10769
timestamp 1745462530
transform 1 0 2484 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_10770
timestamp 1745462530
transform 1 0 2460 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_10771
timestamp 1745462530
transform 1 0 2292 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_10772
timestamp 1745462530
transform 1 0 2204 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_10773
timestamp 1745462530
transform 1 0 2612 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_10774
timestamp 1745462530
transform 1 0 2612 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_10775
timestamp 1745462530
transform 1 0 2612 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_10776
timestamp 1745462530
transform 1 0 2612 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_10777
timestamp 1745462530
transform 1 0 3460 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_10778
timestamp 1745462530
transform 1 0 3388 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_10779
timestamp 1745462530
transform 1 0 3748 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_10780
timestamp 1745462530
transform 1 0 3740 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_10781
timestamp 1745462530
transform 1 0 4308 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_10782
timestamp 1745462530
transform 1 0 4228 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_10783
timestamp 1745462530
transform 1 0 3868 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_10784
timestamp 1745462530
transform 1 0 3788 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_10785
timestamp 1745462530
transform 1 0 4316 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_10786
timestamp 1745462530
transform 1 0 4228 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_10787
timestamp 1745462530
transform 1 0 4156 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_10788
timestamp 1745462530
transform 1 0 4156 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_10789
timestamp 1745462530
transform 1 0 3812 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_10790
timestamp 1745462530
transform 1 0 3804 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_10791
timestamp 1745462530
transform 1 0 3788 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_10792
timestamp 1745462530
transform 1 0 3748 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_10793
timestamp 1745462530
transform 1 0 4220 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_10794
timestamp 1745462530
transform 1 0 4156 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_10795
timestamp 1745462530
transform 1 0 3812 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_10796
timestamp 1745462530
transform 1 0 3804 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_10797
timestamp 1745462530
transform 1 0 4308 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_10798
timestamp 1745462530
transform 1 0 4220 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_10799
timestamp 1745462530
transform 1 0 3900 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_10800
timestamp 1745462530
transform 1 0 3820 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_10801
timestamp 1745462530
transform 1 0 4012 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_10802
timestamp 1745462530
transform 1 0 3996 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_10803
timestamp 1745462530
transform 1 0 3972 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_10804
timestamp 1745462530
transform 1 0 3884 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_10805
timestamp 1745462530
transform 1 0 3084 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_10806
timestamp 1745462530
transform 1 0 2980 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_10807
timestamp 1745462530
transform 1 0 2708 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_10808
timestamp 1745462530
transform 1 0 2588 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_10809
timestamp 1745462530
transform 1 0 3900 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_10810
timestamp 1745462530
transform 1 0 3876 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_10811
timestamp 1745462530
transform 1 0 3772 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_10812
timestamp 1745462530
transform 1 0 3684 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_10813
timestamp 1745462530
transform 1 0 3932 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_10814
timestamp 1745462530
transform 1 0 3868 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_10815
timestamp 1745462530
transform 1 0 3820 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_10816
timestamp 1745462530
transform 1 0 3740 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_10817
timestamp 1745462530
transform 1 0 3916 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_10818
timestamp 1745462530
transform 1 0 3844 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_10819
timestamp 1745462530
transform 1 0 4004 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_10820
timestamp 1745462530
transform 1 0 3940 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_10821
timestamp 1745462530
transform 1 0 3852 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_10822
timestamp 1745462530
transform 1 0 3852 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_10823
timestamp 1745462530
transform 1 0 3092 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_10824
timestamp 1745462530
transform 1 0 2980 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_10825
timestamp 1745462530
transform 1 0 2508 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_10826
timestamp 1745462530
transform 1 0 2444 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_10827
timestamp 1745462530
transform 1 0 1252 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_10828
timestamp 1745462530
transform 1 0 1100 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_10829
timestamp 1745462530
transform 1 0 1236 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_10830
timestamp 1745462530
transform 1 0 1060 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_10831
timestamp 1745462530
transform 1 0 1236 0 1 2737
box -2 -2 2 2
use M2_M1  M2_M1_10832
timestamp 1745462530
transform 1 0 1132 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_10833
timestamp 1745462530
transform 1 0 1212 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_10834
timestamp 1745462530
transform 1 0 1020 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_10835
timestamp 1745462530
transform 1 0 1196 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_10836
timestamp 1745462530
transform 1 0 1100 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_10837
timestamp 1745462530
transform 1 0 1172 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_10838
timestamp 1745462530
transform 1 0 1156 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_10839
timestamp 1745462530
transform 1 0 892 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_10840
timestamp 1745462530
transform 1 0 844 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_10841
timestamp 1745462530
transform 1 0 836 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_10842
timestamp 1745462530
transform 1 0 788 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_10843
timestamp 1745462530
transform 1 0 228 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_10844
timestamp 1745462530
transform 1 0 124 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_10845
timestamp 1745462530
transform 1 0 1004 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_10846
timestamp 1745462530
transform 1 0 964 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_10847
timestamp 1745462530
transform 1 0 212 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_10848
timestamp 1745462530
transform 1 0 140 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_10849
timestamp 1745462530
transform 1 0 220 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_10850
timestamp 1745462530
transform 1 0 140 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_10851
timestamp 1745462530
transform 1 0 220 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_10852
timestamp 1745462530
transform 1 0 140 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_10853
timestamp 1745462530
transform 1 0 820 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_10854
timestamp 1745462530
transform 1 0 692 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_10855
timestamp 1745462530
transform 1 0 228 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_10856
timestamp 1745462530
transform 1 0 132 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_10857
timestamp 1745462530
transform 1 0 212 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_10858
timestamp 1745462530
transform 1 0 116 0 1 1014
box -2 -2 2 2
use M2_M1  M2_M1_10859
timestamp 1745462530
transform 1 0 244 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_10860
timestamp 1745462530
transform 1 0 148 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_10861
timestamp 1745462530
transform 1 0 212 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_10862
timestamp 1745462530
transform 1 0 140 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_10863
timestamp 1745462530
transform 1 0 692 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_10864
timestamp 1745462530
transform 1 0 692 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_10865
timestamp 1745462530
transform 1 0 924 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_10866
timestamp 1745462530
transform 1 0 908 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_10867
timestamp 1745462530
transform 1 0 220 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_10868
timestamp 1745462530
transform 1 0 124 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_10869
timestamp 1745462530
transform 1 0 1044 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_10870
timestamp 1745462530
transform 1 0 956 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_10871
timestamp 1745462530
transform 1 0 1132 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_10872
timestamp 1745462530
transform 1 0 1028 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_10873
timestamp 1745462530
transform 1 0 1164 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_10874
timestamp 1745462530
transform 1 0 1060 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_10875
timestamp 1745462530
transform 1 0 1332 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_10876
timestamp 1745462530
transform 1 0 1244 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_10877
timestamp 1745462530
transform 1 0 1356 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_10878
timestamp 1745462530
transform 1 0 1220 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_10879
timestamp 1745462530
transform 1 0 1428 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_10880
timestamp 1745462530
transform 1 0 1292 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_10881
timestamp 1745462530
transform 1 0 1428 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_10882
timestamp 1745462530
transform 1 0 1332 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_10883
timestamp 1745462530
transform 1 0 1476 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_10884
timestamp 1745462530
transform 1 0 1348 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_10885
timestamp 1745462530
transform 1 0 1532 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_10886
timestamp 1745462530
transform 1 0 1428 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_10887
timestamp 1745462530
transform 1 0 2308 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_10888
timestamp 1745462530
transform 1 0 2148 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_10889
timestamp 1745462530
transform 1 0 2204 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_10890
timestamp 1745462530
transform 1 0 2124 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_10891
timestamp 1745462530
transform 1 0 2308 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_10892
timestamp 1745462530
transform 1 0 2140 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_10893
timestamp 1745462530
transform 1 0 2300 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_10894
timestamp 1745462530
transform 1 0 2156 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_10895
timestamp 1745462530
transform 1 0 2620 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_10896
timestamp 1745462530
transform 1 0 2612 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_10897
timestamp 1745462530
transform 1 0 2636 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_10898
timestamp 1745462530
transform 1 0 2564 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_10899
timestamp 1745462530
transform 1 0 2372 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_10900
timestamp 1745462530
transform 1 0 2372 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_10901
timestamp 1745462530
transform 1 0 2404 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_10902
timestamp 1745462530
transform 1 0 2388 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_10903
timestamp 1745462530
transform 1 0 3332 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_10904
timestamp 1745462530
transform 1 0 3276 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_10905
timestamp 1745462530
transform 1 0 3532 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_10906
timestamp 1745462530
transform 1 0 3460 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_10907
timestamp 1745462530
transform 1 0 4020 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_10908
timestamp 1745462530
transform 1 0 4020 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_10909
timestamp 1745462530
transform 1 0 3524 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_10910
timestamp 1745462530
transform 1 0 3516 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_10911
timestamp 1745462530
transform 1 0 4100 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_10912
timestamp 1745462530
transform 1 0 4004 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_10913
timestamp 1745462530
transform 1 0 3964 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_10914
timestamp 1745462530
transform 1 0 3908 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_10915
timestamp 1745462530
transform 1 0 3460 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_10916
timestamp 1745462530
transform 1 0 3460 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_10917
timestamp 1745462530
transform 1 0 3516 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_10918
timestamp 1745462530
transform 1 0 3460 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_10919
timestamp 1745462530
transform 1 0 4100 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_10920
timestamp 1745462530
transform 1 0 3972 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_10921
timestamp 1745462530
transform 1 0 3484 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_10922
timestamp 1745462530
transform 1 0 3412 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_10923
timestamp 1745462530
transform 1 0 4124 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_10924
timestamp 1745462530
transform 1 0 4124 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_10925
timestamp 1745462530
transform 1 0 3691 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_10926
timestamp 1745462530
transform 1 0 3660 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_10927
timestamp 1745462530
transform 1 0 4148 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_10928
timestamp 1745462530
transform 1 0 4124 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_10929
timestamp 1745462530
transform 1 0 3460 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_10930
timestamp 1745462530
transform 1 0 3388 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_10931
timestamp 1745462530
transform 1 0 2796 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_10932
timestamp 1745462530
transform 1 0 2724 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_10933
timestamp 1745462530
transform 1 0 2636 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_10934
timestamp 1745462530
transform 1 0 2540 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_10935
timestamp 1745462530
transform 1 0 3484 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_10936
timestamp 1745462530
transform 1 0 3452 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_10937
timestamp 1745462530
transform 1 0 3276 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_10938
timestamp 1745462530
transform 1 0 3236 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_10939
timestamp 1745462530
transform 1 0 3404 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_10940
timestamp 1745462530
transform 1 0 3404 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_10941
timestamp 1745462530
transform 1 0 3388 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_10942
timestamp 1745462530
transform 1 0 3300 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_10943
timestamp 1745462530
transform 1 0 3468 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_10944
timestamp 1745462530
transform 1 0 3436 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_10945
timestamp 1745462530
transform 1 0 3444 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_10946
timestamp 1745462530
transform 1 0 3380 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_10947
timestamp 1745462530
transform 1 0 3204 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_10948
timestamp 1745462530
transform 1 0 2892 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_10949
timestamp 1745462530
transform 1 0 2780 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_10950
timestamp 1745462530
transform 1 0 2780 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_10951
timestamp 1745462530
transform 1 0 2700 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_10952
timestamp 1745462530
transform 1 0 2700 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_10953
timestamp 1745462530
transform 1 0 1604 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_10954
timestamp 1745462530
transform 1 0 1596 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_10955
timestamp 1745462530
transform 1 0 1572 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_10956
timestamp 1745462530
transform 1 0 1564 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_10957
timestamp 1745462530
transform 1 0 1556 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_10958
timestamp 1745462530
transform 1 0 1548 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_10959
timestamp 1745462530
transform 1 0 1436 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_10960
timestamp 1745462530
transform 1 0 1420 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_10961
timestamp 1745462530
transform 1 0 1404 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_10962
timestamp 1745462530
transform 1 0 1332 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_10963
timestamp 1745462530
transform 1 0 1372 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_10964
timestamp 1745462530
transform 1 0 1364 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_10965
timestamp 1745462530
transform 1 0 276 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_10966
timestamp 1745462530
transform 1 0 124 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_10967
timestamp 1745462530
transform 1 0 588 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_10968
timestamp 1745462530
transform 1 0 524 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_10969
timestamp 1745462530
transform 1 0 228 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_10970
timestamp 1745462530
transform 1 0 140 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_10971
timestamp 1745462530
transform 1 0 1004 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_10972
timestamp 1745462530
transform 1 0 932 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_10973
timestamp 1745462530
transform 1 0 220 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_10974
timestamp 1745462530
transform 1 0 140 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_10975
timestamp 1745462530
transform 1 0 212 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_10976
timestamp 1745462530
transform 1 0 108 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_10977
timestamp 1745462530
transform 1 0 187 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_10978
timestamp 1745462530
transform 1 0 140 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_10979
timestamp 1745462530
transform 1 0 524 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_10980
timestamp 1745462530
transform 1 0 524 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_10981
timestamp 1745462530
transform 1 0 300 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_10982
timestamp 1745462530
transform 1 0 132 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_10983
timestamp 1745462530
transform 1 0 380 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_10984
timestamp 1745462530
transform 1 0 300 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_10985
timestamp 1745462530
transform 1 0 484 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_10986
timestamp 1745462530
transform 1 0 404 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_10987
timestamp 1745462530
transform 1 0 540 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_10988
timestamp 1745462530
transform 1 0 492 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_10989
timestamp 1745462530
transform 1 0 644 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_10990
timestamp 1745462530
transform 1 0 636 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_10991
timestamp 1745462530
transform 1 0 828 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_10992
timestamp 1745462530
transform 1 0 764 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_10993
timestamp 1745462530
transform 1 0 420 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_10994
timestamp 1745462530
transform 1 0 420 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_10995
timestamp 1745462530
transform 1 0 868 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_10996
timestamp 1745462530
transform 1 0 788 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_10997
timestamp 1745462530
transform 1 0 1116 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_10998
timestamp 1745462530
transform 1 0 1028 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_10999
timestamp 1745462530
transform 1 0 1036 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_11000
timestamp 1745462530
transform 1 0 1004 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_11001
timestamp 1745462530
transform 1 0 1372 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_11002
timestamp 1745462530
transform 1 0 1300 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_11003
timestamp 1745462530
transform 1 0 1268 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_11004
timestamp 1745462530
transform 1 0 1156 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_11005
timestamp 1745462530
transform 1 0 1324 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_11006
timestamp 1745462530
transform 1 0 1220 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_11007
timestamp 1745462530
transform 1 0 1428 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_11008
timestamp 1745462530
transform 1 0 1332 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_11009
timestamp 1745462530
transform 1 0 1420 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_11010
timestamp 1745462530
transform 1 0 1340 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_11011
timestamp 1745462530
transform 1 0 2044 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_11012
timestamp 1745462530
transform 1 0 2036 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_11013
timestamp 1745462530
transform 1 0 2748 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_11014
timestamp 1745462530
transform 1 0 2740 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_11015
timestamp 1745462530
transform 1 0 2852 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_11016
timestamp 1745462530
transform 1 0 2756 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_11017
timestamp 1745462530
transform 1 0 2620 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_11018
timestamp 1745462530
transform 1 0 2604 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_11019
timestamp 1745462530
transform 1 0 2780 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_11020
timestamp 1745462530
transform 1 0 2772 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_11021
timestamp 1745462530
transform 1 0 3044 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_11022
timestamp 1745462530
transform 1 0 3044 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_11023
timestamp 1745462530
transform 1 0 2732 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_11024
timestamp 1745462530
transform 1 0 2732 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_11025
timestamp 1745462530
transform 1 0 2692 0 1 1214
box -2 -2 2 2
use M2_M1  M2_M1_11026
timestamp 1745462530
transform 1 0 2684 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_11027
timestamp 1745462530
transform 1 0 2700 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_11028
timestamp 1745462530
transform 1 0 2644 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_11029
timestamp 1745462530
transform 1 0 3260 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_11030
timestamp 1745462530
transform 1 0 3220 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_11031
timestamp 1745462530
transform 1 0 3596 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_11032
timestamp 1745462530
transform 1 0 3548 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_11033
timestamp 1745462530
transform 1 0 3756 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_11034
timestamp 1745462530
transform 1 0 3732 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_11035
timestamp 1745462530
transform 1 0 3652 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_11036
timestamp 1745462530
transform 1 0 3652 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_11037
timestamp 1745462530
transform 1 0 4332 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_11038
timestamp 1745462530
transform 1 0 4332 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_11039
timestamp 1745462530
transform 1 0 4308 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_11040
timestamp 1745462530
transform 1 0 4236 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_11041
timestamp 1745462530
transform 1 0 4164 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_11042
timestamp 1745462530
transform 1 0 4140 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_11043
timestamp 1745462530
transform 1 0 3620 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_11044
timestamp 1745462530
transform 1 0 3620 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_11045
timestamp 1745462530
transform 1 0 4308 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_11046
timestamp 1745462530
transform 1 0 4228 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_11047
timestamp 1745462530
transform 1 0 3692 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_11048
timestamp 1745462530
transform 1 0 3596 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_11049
timestamp 1745462530
transform 1 0 4316 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_11050
timestamp 1745462530
transform 1 0 4228 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_11051
timestamp 1745462530
transform 1 0 3788 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_11052
timestamp 1745462530
transform 1 0 3748 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_11053
timestamp 1745462530
transform 1 0 4316 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_11054
timestamp 1745462530
transform 1 0 4300 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_11055
timestamp 1745462530
transform 1 0 3668 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_11056
timestamp 1745462530
transform 1 0 3588 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_11057
timestamp 1745462530
transform 1 0 2844 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_11058
timestamp 1745462530
transform 1 0 2844 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_11059
timestamp 1745462530
transform 1 0 2652 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_11060
timestamp 1745462530
transform 1 0 2644 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_11061
timestamp 1745462530
transform 1 0 3684 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_11062
timestamp 1745462530
transform 1 0 3684 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_11063
timestamp 1745462530
transform 1 0 3708 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_11064
timestamp 1745462530
transform 1 0 3620 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_11065
timestamp 1745462530
transform 1 0 3708 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_11066
timestamp 1745462530
transform 1 0 3636 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_11067
timestamp 1745462530
transform 1 0 3628 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_11068
timestamp 1745462530
transform 1 0 3540 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_11069
timestamp 1745462530
transform 1 0 3740 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_11070
timestamp 1745462530
transform 1 0 3668 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_11071
timestamp 1745462530
transform 1 0 3700 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_11072
timestamp 1745462530
transform 1 0 3628 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_11073
timestamp 1745462530
transform 1 0 3492 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_11074
timestamp 1745462530
transform 1 0 3476 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_11075
timestamp 1745462530
transform 1 0 2988 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_11076
timestamp 1745462530
transform 1 0 2876 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_11077
timestamp 1745462530
transform 1 0 2636 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_11078
timestamp 1745462530
transform 1 0 2572 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_11079
timestamp 1745462530
transform 1 0 2404 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_11080
timestamp 1745462530
transform 1 0 2340 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_11081
timestamp 1745462530
transform 1 0 2308 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_11082
timestamp 1745462530
transform 1 0 2252 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_11083
timestamp 1745462530
transform 1 0 2228 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_11084
timestamp 1745462530
transform 1 0 2172 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_11085
timestamp 1745462530
transform 1 0 2076 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_11086
timestamp 1745462530
transform 1 0 2028 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_11087
timestamp 1745462530
transform 1 0 2292 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_11088
timestamp 1745462530
transform 1 0 2252 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_11089
timestamp 1745462530
transform 1 0 2124 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_11090
timestamp 1745462530
transform 1 0 2124 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_11091
timestamp 1745462530
transform 1 0 724 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_11092
timestamp 1745462530
transform 1 0 724 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_11093
timestamp 1745462530
transform 1 0 1324 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_11094
timestamp 1745462530
transform 1 0 1228 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_11095
timestamp 1745462530
transform 1 0 412 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_11096
timestamp 1745462530
transform 1 0 412 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_11097
timestamp 1745462530
transform 1 0 1132 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_11098
timestamp 1745462530
transform 1 0 1076 0 1 4105
box -2 -2 2 2
use M2_M1  M2_M1_11099
timestamp 1745462530
transform 1 0 1076 0 1 4035
box -2 -2 2 2
use M2_M1  M2_M1_11100
timestamp 1745462530
transform 1 0 1068 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_11101
timestamp 1745462530
transform 1 0 1060 0 1 4005
box -2 -2 2 2
use M2_M1  M2_M1_11102
timestamp 1745462530
transform 1 0 1004 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_11103
timestamp 1745462530
transform 1 0 1148 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_11104
timestamp 1745462530
transform 1 0 1116 0 1 4145
box -2 -2 2 2
use M2_M1  M2_M1_11105
timestamp 1745462530
transform 1 0 1084 0 1 4115
box -2 -2 2 2
use M2_M1  M2_M1_11106
timestamp 1745462530
transform 1 0 1084 0 1 4025
box -2 -2 2 2
use M2_M1  M2_M1_11107
timestamp 1745462530
transform 1 0 1020 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_11108
timestamp 1745462530
transform 1 0 908 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_11109
timestamp 1745462530
transform 1 0 4068 0 1 4225
box -2 -2 2 2
use M2_M1  M2_M1_11110
timestamp 1745462530
transform 1 0 4036 0 1 4225
box -2 -2 2 2
use M2_M1  M2_M1_11111
timestamp 1745462530
transform 1 0 4036 0 1 4025
box -2 -2 2 2
use M2_M1  M2_M1_11112
timestamp 1745462530
transform 1 0 4036 0 1 3915
box -2 -2 2 2
use M2_M1  M2_M1_11113
timestamp 1745462530
transform 1 0 2987 0 1 4225
box -2 -2 2 2
use M2_M1  M2_M1_11114
timestamp 1745462530
transform 1 0 2612 0 1 4225
box -2 -2 2 2
use M2_M1  M2_M1_11115
timestamp 1745462530
transform 1 0 2020 0 1 4225
box -2 -2 2 2
use M2_M1  M2_M1_11116
timestamp 1745462530
transform 1 0 1852 0 1 4225
box -2 -2 2 2
use M2_M1  M2_M1_11117
timestamp 1745462530
transform 1 0 1308 0 1 4005
box -2 -2 2 2
use M2_M1  M2_M1_11118
timestamp 1745462530
transform 1 0 1212 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_11119
timestamp 1745462530
transform 1 0 1084 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_11120
timestamp 1745462530
transform 1 0 1036 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_11121
timestamp 1745462530
transform 1 0 948 0 1 4105
box -2 -2 2 2
use M2_M1  M2_M1_11122
timestamp 1745462530
transform 1 0 940 0 1 4005
box -2 -2 2 2
use M2_M1  M2_M1_11123
timestamp 1745462530
transform 1 0 852 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_11124
timestamp 1745462530
transform 1 0 732 0 1 4105
box -2 -2 2 2
use M2_M1  M2_M1_11125
timestamp 1745462530
transform 1 0 628 0 1 4195
box -2 -2 2 2
use M2_M1  M2_M1_11126
timestamp 1745462530
transform 1 0 564 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_11127
timestamp 1745462530
transform 1 0 844 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_11128
timestamp 1745462530
transform 1 0 788 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_11129
timestamp 1745462530
transform 1 0 732 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_11130
timestamp 1745462530
transform 1 0 468 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_11131
timestamp 1745462530
transform 1 0 772 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_11132
timestamp 1745462530
transform 1 0 492 0 1 4005
box -2 -2 2 2
use M2_M1  M2_M1_11133
timestamp 1745462530
transform 1 0 1284 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_11134
timestamp 1745462530
transform 1 0 1236 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_11135
timestamp 1745462530
transform 1 0 1164 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_11136
timestamp 1745462530
transform 1 0 1164 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_11137
timestamp 1745462530
transform 1 0 1236 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_11138
timestamp 1745462530
transform 1 0 1220 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_11139
timestamp 1745462530
transform 1 0 1140 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_11140
timestamp 1745462530
transform 1 0 1068 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_11141
timestamp 1745462530
transform 1 0 1284 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_11142
timestamp 1745462530
transform 1 0 1268 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_11143
timestamp 1745462530
transform 1 0 1156 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_11144
timestamp 1745462530
transform 1 0 1156 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_11145
timestamp 1745462530
transform 1 0 1028 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_11146
timestamp 1745462530
transform 1 0 988 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_11147
timestamp 1745462530
transform 1 0 780 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_11148
timestamp 1745462530
transform 1 0 772 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_11149
timestamp 1745462530
transform 1 0 1748 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_11150
timestamp 1745462530
transform 1 0 1676 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_11151
timestamp 1745462530
transform 1 0 1588 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_11152
timestamp 1745462530
transform 1 0 1588 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_11153
timestamp 1745462530
transform 1 0 4316 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_11154
timestamp 1745462530
transform 1 0 4268 0 1 4005
box -2 -2 2 2
use M2_M1  M2_M1_11155
timestamp 1745462530
transform 1 0 4308 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_11156
timestamp 1745462530
transform 1 0 4268 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_11157
timestamp 1745462530
transform 1 0 4308 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_11158
timestamp 1745462530
transform 1 0 4268 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_11159
timestamp 1745462530
transform 1 0 4204 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_11160
timestamp 1745462530
transform 1 0 4172 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_11161
timestamp 1745462530
transform 1 0 1492 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_11162
timestamp 1745462530
transform 1 0 1444 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_11163
timestamp 1745462530
transform 1 0 1396 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_11164
timestamp 1745462530
transform 1 0 1356 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_11165
timestamp 1745462530
transform 1 0 780 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_11166
timestamp 1745462530
transform 1 0 644 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_11167
timestamp 1745462530
transform 1 0 612 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_11168
timestamp 1745462530
transform 1 0 588 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_11169
timestamp 1745462530
transform 1 0 740 0 1 4115
box -2 -2 2 2
use M2_M1  M2_M1_11170
timestamp 1745462530
transform 1 0 684 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_11171
timestamp 1745462530
transform 1 0 668 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_11172
timestamp 1745462530
transform 1 0 684 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_11173
timestamp 1745462530
transform 1 0 612 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_11174
timestamp 1745462530
transform 1 0 684 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_11175
timestamp 1745462530
transform 1 0 660 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_11176
timestamp 1745462530
transform 1 0 908 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_11177
timestamp 1745462530
transform 1 0 868 0 1 4025
box -2 -2 2 2
use M2_M1  M2_M1_11178
timestamp 1745462530
transform 1 0 860 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_11179
timestamp 1745462530
transform 1 0 836 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_11180
timestamp 1745462530
transform 1 0 748 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_11181
timestamp 1745462530
transform 1 0 716 0 1 4025
box -2 -2 2 2
use M2_M1  M2_M1_11182
timestamp 1745462530
transform 1 0 692 0 1 4145
box -2 -2 2 2
use M2_M1  M2_M1_11183
timestamp 1745462530
transform 1 0 660 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_11184
timestamp 1745462530
transform 1 0 4212 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_11185
timestamp 1745462530
transform 1 0 4212 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_11186
timestamp 1745462530
transform 1 0 4212 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_11187
timestamp 1745462530
transform 1 0 4124 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_11188
timestamp 1745462530
transform 1 0 1716 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_11189
timestamp 1745462530
transform 1 0 1556 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_11190
timestamp 1745462530
transform 1 0 1500 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_11191
timestamp 1745462530
transform 1 0 1436 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_11192
timestamp 1745462530
transform 1 0 1108 0 1 4035
box -2 -2 2 2
use M2_M1  M2_M1_11193
timestamp 1745462530
transform 1 0 812 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_11194
timestamp 1745462530
transform 1 0 764 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_11195
timestamp 1745462530
transform 1 0 1372 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_11196
timestamp 1745462530
transform 1 0 1028 0 1 4115
box -2 -2 2 2
use M2_M1  M2_M1_11197
timestamp 1745462530
transform 1 0 876 0 1 4115
box -2 -2 2 2
use M2_M1  M2_M1_11198
timestamp 1745462530
transform 1 0 876 0 1 4025
box -2 -2 2 2
use M2_M1  M2_M1_11199
timestamp 1745462530
transform 1 0 956 0 1 4115
box -2 -2 2 2
use M2_M1  M2_M1_11200
timestamp 1745462530
transform 1 0 924 0 1 4115
box -2 -2 2 2
use M2_M1  M2_M1_11201
timestamp 1745462530
transform 1 0 452 0 1 4005
box -2 -2 2 2
use M2_M1  M2_M1_11202
timestamp 1745462530
transform 1 0 388 0 1 4005
box -2 -2 2 2
use M2_M1  M2_M1_11203
timestamp 1745462530
transform 1 0 332 0 1 4025
box -2 -2 2 2
use M2_M1  M2_M1_11204
timestamp 1745462530
transform 1 0 324 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_11205
timestamp 1745462530
transform 1 0 364 0 1 4005
box -2 -2 2 2
use M2_M1  M2_M1_11206
timestamp 1745462530
transform 1 0 324 0 1 4035
box -2 -2 2 2
use M2_M1  M2_M1_11207
timestamp 1745462530
transform 1 0 372 0 1 4025
box -2 -2 2 2
use M2_M1  M2_M1_11208
timestamp 1745462530
transform 1 0 300 0 1 4005
box -2 -2 2 2
use M2_M1  M2_M1_11209
timestamp 1745462530
transform 1 0 268 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_11210
timestamp 1745462530
transform 1 0 228 0 1 4225
box -2 -2 2 2
use M2_M1  M2_M1_11211
timestamp 1745462530
transform 1 0 84 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_11212
timestamp 1745462530
transform 1 0 588 0 1 4005
box -2 -2 2 2
use M2_M1  M2_M1_11213
timestamp 1745462530
transform 1 0 508 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_11214
timestamp 1745462530
transform 1 0 532 0 1 4005
box -2 -2 2 2
use M2_M1  M2_M1_11215
timestamp 1745462530
transform 1 0 516 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_11216
timestamp 1745462530
transform 1 0 508 0 1 4005
box -2 -2 2 2
use M2_M1  M2_M1_11217
timestamp 1745462530
transform 1 0 476 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_11218
timestamp 1745462530
transform 1 0 636 0 1 4115
box -2 -2 2 2
use M2_M1  M2_M1_11219
timestamp 1745462530
transform 1 0 612 0 1 4005
box -2 -2 2 2
use M2_M1  M2_M1_11220
timestamp 1745462530
transform 1 0 572 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_11221
timestamp 1745462530
transform 1 0 684 0 1 4025
box -2 -2 2 2
use M2_M1  M2_M1_11222
timestamp 1745462530
transform 1 0 628 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_11223
timestamp 1745462530
transform 1 0 612 0 1 3915
box -2 -2 2 2
use M2_M1  M2_M1_11224
timestamp 1745462530
transform 1 0 580 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_11225
timestamp 1745462530
transform 1 0 220 0 1 4025
box -2 -2 2 2
use M2_M1  M2_M1_11226
timestamp 1745462530
transform 1 0 188 0 1 3915
box -2 -2 2 2
use M2_M1  M2_M1_11227
timestamp 1745462530
transform 1 0 148 0 1 4115
box -2 -2 2 2
use M2_M1  M2_M1_11228
timestamp 1745462530
transform 1 0 212 0 1 4035
box -2 -2 2 2
use M2_M1  M2_M1_11229
timestamp 1745462530
transform 1 0 188 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_11230
timestamp 1745462530
transform 1 0 220 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_11231
timestamp 1745462530
transform 1 0 172 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_11232
timestamp 1745462530
transform 1 0 180 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_11233
timestamp 1745462530
transform 1 0 148 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_11234
timestamp 1745462530
transform 1 0 220 0 1 3825
box -2 -2 2 2
use M2_M1  M2_M1_11235
timestamp 1745462530
transform 1 0 196 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_11236
timestamp 1745462530
transform 1 0 148 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_11237
timestamp 1745462530
transform 1 0 140 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_11238
timestamp 1745462530
transform 1 0 140 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_11239
timestamp 1745462530
transform 1 0 116 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_11240
timestamp 1745462530
transform 1 0 156 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_11241
timestamp 1745462530
transform 1 0 124 0 1 4105
box -2 -2 2 2
use M2_M1  M2_M1_11242
timestamp 1745462530
transform 1 0 116 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_11243
timestamp 1745462530
transform 1 0 84 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_11244
timestamp 1745462530
transform 1 0 100 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_11245
timestamp 1745462530
transform 1 0 68 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_11246
timestamp 1745462530
transform 1 0 108 0 1 4025
box -2 -2 2 2
use M2_M1  M2_M1_11247
timestamp 1745462530
transform 1 0 108 0 1 3915
box -2 -2 2 2
use M2_M1  M2_M1_11248
timestamp 1745462530
transform 1 0 84 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_11249
timestamp 1745462530
transform 1 0 68 0 1 4105
box -2 -2 2 2
use M2_M1  M2_M1_11250
timestamp 1745462530
transform 1 0 68 0 1 4035
box -2 -2 2 2
use M2_M1  M2_M1_11251
timestamp 1745462530
transform 1 0 1484 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_11252
timestamp 1745462530
transform 1 0 1404 0 1 4145
box -2 -2 2 2
use M2_M1  M2_M1_11253
timestamp 1745462530
transform 1 0 1460 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_11254
timestamp 1745462530
transform 1 0 1428 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_11255
timestamp 1745462530
transform 1 0 4244 0 1 4115
box -2 -2 2 2
use M2_M1  M2_M1_11256
timestamp 1745462530
transform 1 0 4228 0 1 4025
box -2 -2 2 2
use M2_M1  M2_M1_11257
timestamp 1745462530
transform 1 0 4228 0 1 3915
box -2 -2 2 2
use M2_M1  M2_M1_11258
timestamp 1745462530
transform 1 0 4140 0 1 4115
box -2 -2 2 2
use M2_M1  M2_M1_11259
timestamp 1745462530
transform 1 0 1732 0 1 4115
box -2 -2 2 2
use M2_M1  M2_M1_11260
timestamp 1745462530
transform 1 0 1572 0 1 4115
box -2 -2 2 2
use M2_M1  M2_M1_11261
timestamp 1745462530
transform 1 0 1516 0 1 4115
box -2 -2 2 2
use M2_M1  M2_M1_11262
timestamp 1745462530
transform 1 0 1452 0 1 4115
box -2 -2 2 2
use M2_M1  M2_M1_11263
timestamp 1745462530
transform 1 0 852 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_11264
timestamp 1745462530
transform 1 0 4172 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_11265
timestamp 1745462530
transform 1 0 4172 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_11266
timestamp 1745462530
transform 1 0 4172 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_11267
timestamp 1745462530
transform 1 0 4084 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_11268
timestamp 1745462530
transform 1 0 1788 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_11269
timestamp 1745462530
transform 1 0 1772 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_11270
timestamp 1745462530
transform 1 0 1524 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_11271
timestamp 1745462530
transform 1 0 1468 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_11272
timestamp 1745462530
transform 1 0 1100 0 1 4115
box -2 -2 2 2
use M2_M1  M2_M1_11273
timestamp 1745462530
transform 1 0 1068 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_11274
timestamp 1745462530
transform 1 0 1860 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_11275
timestamp 1745462530
transform 1 0 1484 0 1 4115
box -2 -2 2 2
use M2_M1  M2_M1_11276
timestamp 1745462530
transform 1 0 1852 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_11277
timestamp 1745462530
transform 1 0 1836 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_11278
timestamp 1745462530
transform 1 0 1892 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_11279
timestamp 1745462530
transform 1 0 1844 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_11280
timestamp 1745462530
transform 1 0 1908 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_11281
timestamp 1745462530
transform 1 0 1868 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_11282
timestamp 1745462530
transform 1 0 2036 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_11283
timestamp 1745462530
transform 1 0 1868 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_11284
timestamp 1745462530
transform 1 0 1868 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_11285
timestamp 1745462530
transform 1 0 1828 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_11286
timestamp 1745462530
transform 1 0 2140 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_11287
timestamp 1745462530
transform 1 0 1820 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_11288
timestamp 1745462530
transform 1 0 1540 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_11289
timestamp 1745462530
transform 1 0 1492 0 1 4195
box -2 -2 2 2
use M2_M1  M2_M1_11290
timestamp 1745462530
transform 1 0 1516 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_11291
timestamp 1745462530
transform 1 0 1508 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_11292
timestamp 1745462530
transform 1 0 1908 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_11293
timestamp 1745462530
transform 1 0 1540 0 1 4225
box -2 -2 2 2
use M2_M1  M2_M1_11294
timestamp 1745462530
transform 1 0 2020 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_11295
timestamp 1745462530
transform 1 0 1884 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_11296
timestamp 1745462530
transform 1 0 1940 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_11297
timestamp 1745462530
transform 1 0 1892 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_11298
timestamp 1745462530
transform 1 0 1940 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_11299
timestamp 1745462530
transform 1 0 1916 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_11300
timestamp 1745462530
transform 1 0 2180 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_11301
timestamp 1745462530
transform 1 0 1924 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_11302
timestamp 1745462530
transform 1 0 2316 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_11303
timestamp 1745462530
transform 1 0 1996 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_11304
timestamp 1745462530
transform 1 0 4148 0 1 4145
box -2 -2 2 2
use M2_M1  M2_M1_11305
timestamp 1745462530
transform 1 0 4108 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_11306
timestamp 1745462530
transform 1 0 4164 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_11307
timestamp 1745462530
transform 1 0 4148 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_11308
timestamp 1745462530
transform 1 0 4100 0 1 4115
box -2 -2 2 2
use M2_M1  M2_M1_11309
timestamp 1745462530
transform 1 0 4044 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_11310
timestamp 1745462530
transform 1 0 4036 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_11311
timestamp 1745462530
transform 1 0 4012 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_11312
timestamp 1745462530
transform 1 0 4020 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_11313
timestamp 1745462530
transform 1 0 3988 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_11314
timestamp 1745462530
transform 1 0 3948 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_11315
timestamp 1745462530
transform 1 0 3340 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_11316
timestamp 1745462530
transform 1 0 4012 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_11317
timestamp 1745462530
transform 1 0 4004 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_11318
timestamp 1745462530
transform 1 0 4012 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_11319
timestamp 1745462530
transform 1 0 3836 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_11320
timestamp 1745462530
transform 1 0 4236 0 1 3945
box -2 -2 2 2
use M2_M1  M2_M1_11321
timestamp 1745462530
transform 1 0 4196 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_11322
timestamp 1745462530
transform 1 0 4252 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_11323
timestamp 1745462530
transform 1 0 4236 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_11324
timestamp 1745462530
transform 1 0 4196 0 1 3915
box -2 -2 2 2
use M2_M1  M2_M1_11325
timestamp 1745462530
transform 1 0 4076 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_11326
timestamp 1745462530
transform 1 0 4044 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_11327
timestamp 1745462530
transform 1 0 4004 0 1 4005
box -2 -2 2 2
use M2_M1  M2_M1_11328
timestamp 1745462530
transform 1 0 4092 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_11329
timestamp 1745462530
transform 1 0 3956 0 1 4005
box -2 -2 2 2
use M2_M1  M2_M1_11330
timestamp 1745462530
transform 1 0 3932 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_11331
timestamp 1745462530
transform 1 0 3660 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_11332
timestamp 1745462530
transform 1 0 4068 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_11333
timestamp 1745462530
transform 1 0 3996 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_11334
timestamp 1745462530
transform 1 0 4004 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_11335
timestamp 1745462530
transform 1 0 3788 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_11336
timestamp 1745462530
transform 1 0 4252 0 1 4145
box -2 -2 2 2
use M2_M1  M2_M1_11337
timestamp 1745462530
transform 1 0 4212 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_11338
timestamp 1745462530
transform 1 0 4268 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_11339
timestamp 1745462530
transform 1 0 4252 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_11340
timestamp 1745462530
transform 1 0 4204 0 1 4115
box -2 -2 2 2
use M2_M1  M2_M1_11341
timestamp 1745462530
transform 1 0 4164 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_11342
timestamp 1745462530
transform 1 0 4132 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_11343
timestamp 1745462530
transform 1 0 4068 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_11344
timestamp 1745462530
transform 1 0 4140 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_11345
timestamp 1745462530
transform 1 0 4100 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_11346
timestamp 1745462530
transform 1 0 4100 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_11347
timestamp 1745462530
transform 1 0 4076 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_11348
timestamp 1745462530
transform 1 0 4076 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_11349
timestamp 1745462530
transform 1 0 3508 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_11350
timestamp 1745462530
transform 1 0 4092 0 1 4005
box -2 -2 2 2
use M2_M1  M2_M1_11351
timestamp 1745462530
transform 1 0 4044 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_11352
timestamp 1745462530
transform 1 0 4036 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_11353
timestamp 1745462530
transform 1 0 3876 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_11354
timestamp 1745462530
transform 1 0 4236 0 1 3995
box -2 -2 2 2
use M2_M1  M2_M1_11355
timestamp 1745462530
transform 1 0 4196 0 1 4005
box -2 -2 2 2
use M2_M1  M2_M1_11356
timestamp 1745462530
transform 1 0 4252 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_11357
timestamp 1745462530
transform 1 0 4236 0 1 4005
box -2 -2 2 2
use M2_M1  M2_M1_11358
timestamp 1745462530
transform 1 0 4196 0 1 4025
box -2 -2 2 2
use M2_M1  M2_M1_11359
timestamp 1745462530
transform 1 0 4100 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_11360
timestamp 1745462530
transform 1 0 4068 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_11361
timestamp 1745462530
transform 1 0 4060 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_11362
timestamp 1745462530
transform 1 0 4132 0 1 4005
box -2 -2 2 2
use M2_M1  M2_M1_11363
timestamp 1745462530
transform 1 0 4044 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_11364
timestamp 1745462530
transform 1 0 4052 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_11365
timestamp 1745462530
transform 1 0 3604 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_11366
timestamp 1745462530
transform 1 0 4116 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_11367
timestamp 1745462530
transform 1 0 4012 0 1 4005
box -2 -2 2 2
use M2_M1  M2_M1_11368
timestamp 1745462530
transform 1 0 4004 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_11369
timestamp 1745462530
transform 1 0 3828 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_11370
timestamp 1745462530
transform 1 0 1788 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_11371
timestamp 1745462530
transform 1 0 1580 0 1 4145
box -2 -2 2 2
use M2_M1  M2_M1_11372
timestamp 1745462530
transform 1 0 1596 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_11373
timestamp 1745462530
transform 1 0 1580 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_11374
timestamp 1745462530
transform 1 0 2876 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_11375
timestamp 1745462530
transform 1 0 1788 0 1 4225
box -2 -2 2 2
use M2_M1  M2_M1_11376
timestamp 1745462530
transform 1 0 2996 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_11377
timestamp 1745462530
transform 1 0 2852 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_11378
timestamp 1745462530
transform 1 0 2908 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_11379
timestamp 1745462530
transform 1 0 2860 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_11380
timestamp 1745462530
transform 1 0 2908 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_11381
timestamp 1745462530
transform 1 0 2884 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_11382
timestamp 1745462530
transform 1 0 3052 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_11383
timestamp 1745462530
transform 1 0 2892 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_11384
timestamp 1745462530
transform 1 0 3012 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_11385
timestamp 1745462530
transform 1 0 2972 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_11386
timestamp 1745462530
transform 1 0 1820 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_11387
timestamp 1745462530
transform 1 0 1740 0 1 4195
box -2 -2 2 2
use M2_M1  M2_M1_11388
timestamp 1745462530
transform 1 0 1756 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_11389
timestamp 1745462530
transform 1 0 1732 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_11390
timestamp 1745462530
transform 1 0 2556 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_11391
timestamp 1745462530
transform 1 0 1820 0 1 4225
box -2 -2 2 2
use M2_M1  M2_M1_11392
timestamp 1745462530
transform 1 0 2612 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_11393
timestamp 1745462530
transform 1 0 2532 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_11394
timestamp 1745462530
transform 1 0 2668 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_11395
timestamp 1745462530
transform 1 0 2540 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_11396
timestamp 1745462530
transform 1 0 2828 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_11397
timestamp 1745462530
transform 1 0 2652 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_11398
timestamp 1745462530
transform 1 0 2692 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_11399
timestamp 1745462530
transform 1 0 2588 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_11400
timestamp 1745462530
transform 1 0 1524 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_11401
timestamp 1745462530
transform 1 0 1244 0 1 4115
box -2 -2 2 2
use M2_M1  M2_M1_11402
timestamp 1745462530
transform 1 0 1188 0 1 4115
box -2 -2 2 2
use M2_M1  M2_M1_11403
timestamp 1745462530
transform 1 0 1124 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_11404
timestamp 1745462530
transform 1 0 1380 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_11405
timestamp 1745462530
transform 1 0 1220 0 1 4115
box -2 -2 2 2
use M2_M1  M2_M1_11406
timestamp 1745462530
transform 1 0 1164 0 1 4115
box -2 -2 2 2
use M2_M1  M2_M1_11407
timestamp 1745462530
transform 1 0 1060 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_11408
timestamp 1745462530
transform 1 0 1364 0 1 4005
box -2 -2 2 2
use M2_M1  M2_M1_11409
timestamp 1745462530
transform 1 0 1308 0 1 4025
box -2 -2 2 2
use M2_M1  M2_M1_11410
timestamp 1745462530
transform 1 0 1180 0 1 4025
box -2 -2 2 2
use M2_M1  M2_M1_11411
timestamp 1745462530
transform 1 0 1140 0 1 4005
box -2 -2 2 2
use M2_M1  M2_M1_11412
timestamp 1745462530
transform 1 0 1236 0 1 4005
box -2 -2 2 2
use M2_M1  M2_M1_11413
timestamp 1745462530
transform 1 0 1180 0 1 4005
box -2 -2 2 2
use M2_M1  M2_M1_11414
timestamp 1745462530
transform 1 0 1028 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_11415
timestamp 1745462530
transform 1 0 788 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_11416
timestamp 1745462530
transform 1 0 780 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_11417
timestamp 1745462530
transform 1 0 1228 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_11418
timestamp 1745462530
transform 1 0 1172 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_11419
timestamp 1745462530
transform 1 0 1164 0 1 4005
box -2 -2 2 2
use M2_M1  M2_M1_11420
timestamp 1745462530
transform 1 0 1148 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_11421
timestamp 1745462530
transform 1 0 1284 0 1 3995
box -2 -2 2 2
use M2_M1  M2_M1_11422
timestamp 1745462530
transform 1 0 1276 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_11423
timestamp 1745462530
transform 1 0 1228 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_11424
timestamp 1745462530
transform 1 0 1204 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_11425
timestamp 1745462530
transform 1 0 500 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_11426
timestamp 1745462530
transform 1 0 500 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_11427
timestamp 1745462530
transform 1 0 660 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_11428
timestamp 1745462530
transform 1 0 548 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_11429
timestamp 1745462530
transform 1 0 604 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_11430
timestamp 1745462530
transform 1 0 516 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_11431
timestamp 1745462530
transform 1 0 996 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_11432
timestamp 1745462530
transform 1 0 972 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_11433
timestamp 1745462530
transform 1 0 980 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_11434
timestamp 1745462530
transform 1 0 900 0 1 4005
box -2 -2 2 2
use M2_M1  M2_M1_11435
timestamp 1745462530
transform 1 0 924 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_11436
timestamp 1745462530
transform 1 0 876 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_11437
timestamp 1745462530
transform 1 0 812 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_11438
timestamp 1745462530
transform 1 0 772 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_11439
timestamp 1745462530
transform 1 0 404 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_11440
timestamp 1745462530
transform 1 0 524 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_11441
timestamp 1745462530
transform 1 0 276 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_11442
timestamp 1745462530
transform 1 0 228 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_11443
timestamp 1745462530
transform 1 0 652 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_11444
timestamp 1745462530
transform 1 0 340 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_11445
timestamp 1745462530
transform 1 0 236 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_11446
timestamp 1745462530
transform 1 0 172 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_11447
timestamp 1745462530
transform 1 0 84 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_11448
timestamp 1745462530
transform 1 0 524 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_11449
timestamp 1745462530
transform 1 0 220 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_11450
timestamp 1745462530
transform 1 0 172 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_11451
timestamp 1745462530
transform 1 0 604 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_11452
timestamp 1745462530
transform 1 0 236 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_11453
timestamp 1745462530
transform 1 0 220 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_11454
timestamp 1745462530
transform 1 0 180 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_11455
timestamp 1745462530
transform 1 0 660 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_11456
timestamp 1745462530
transform 1 0 372 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_11457
timestamp 1745462530
transform 1 0 348 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_11458
timestamp 1745462530
transform 1 0 244 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_11459
timestamp 1745462530
transform 1 0 484 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_11460
timestamp 1745462530
transform 1 0 484 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_11461
timestamp 1745462530
transform 1 0 404 0 1 3505
box -2 -2 2 2
use M2_M1  M2_M1_11462
timestamp 1745462530
transform 1 0 324 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_11463
timestamp 1745462530
transform 1 0 2868 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_11464
timestamp 1745462530
transform 1 0 2844 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_11465
timestamp 1745462530
transform 1 0 2812 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_11466
timestamp 1745462530
transform 1 0 3100 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_11467
timestamp 1745462530
transform 1 0 3068 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_11468
timestamp 1745462530
transform 1 0 3020 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_11469
timestamp 1745462530
transform 1 0 3620 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_11470
timestamp 1745462530
transform 1 0 3436 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_11471
timestamp 1745462530
transform 1 0 3420 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_11472
timestamp 1745462530
transform 1 0 3524 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_11473
timestamp 1745462530
transform 1 0 3452 0 1 4005
box -2 -2 2 2
use M2_M1  M2_M1_11474
timestamp 1745462530
transform 1 0 3324 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_11475
timestamp 1745462530
transform 1 0 3676 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_11476
timestamp 1745462530
transform 1 0 3420 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_11477
timestamp 1745462530
transform 1 0 3332 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_11478
timestamp 1745462530
transform 1 0 3356 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_11479
timestamp 1745462530
transform 1 0 3212 0 1 4005
box -2 -2 2 2
use M2_M1  M2_M1_11480
timestamp 1745462530
transform 1 0 3212 0 1 3955
box -2 -2 2 2
use M2_M1  M2_M1_11481
timestamp 1745462530
transform 1 0 2548 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_11482
timestamp 1745462530
transform 1 0 2364 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_11483
timestamp 1745462530
transform 1 0 2196 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_11484
timestamp 1745462530
transform 1 0 2156 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_11485
timestamp 1745462530
transform 1 0 2068 0 1 4005
box -2 -2 2 2
use M2_M1  M2_M1_11486
timestamp 1745462530
transform 1 0 2052 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_11487
timestamp 1745462530
transform 1 0 2828 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_11488
timestamp 1745462530
transform 1 0 2716 0 1 4005
box -2 -2 2 2
use M2_M1  M2_M1_11489
timestamp 1745462530
transform 1 0 2708 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_11490
timestamp 1745462530
transform 1 0 3164 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_11491
timestamp 1745462530
transform 1 0 3084 0 1 4005
box -2 -2 2 2
use M2_M1  M2_M1_11492
timestamp 1745462530
transform 1 0 3028 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_11493
timestamp 1745462530
transform 1 0 3916 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_11494
timestamp 1745462530
transform 1 0 3844 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_11495
timestamp 1745462530
transform 1 0 3676 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_11496
timestamp 1745462530
transform 1 0 3892 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_11497
timestamp 1745462530
transform 1 0 3716 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_11498
timestamp 1745462530
transform 1 0 3628 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_11499
timestamp 1745462530
transform 1 0 3804 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_11500
timestamp 1745462530
transform 1 0 3804 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_11501
timestamp 1745462530
transform 1 0 3692 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_11502
timestamp 1745462530
transform 1 0 3852 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_11503
timestamp 1745462530
transform 1 0 3372 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_11504
timestamp 1745462530
transform 1 0 3284 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_11505
timestamp 1745462530
transform 1 0 2548 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_11506
timestamp 1745462530
transform 1 0 2340 0 1 4005
box -2 -2 2 2
use M2_M1  M2_M1_11507
timestamp 1745462530
transform 1 0 2332 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_11508
timestamp 1745462530
transform 1 0 2332 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_11509
timestamp 1745462530
transform 1 0 2204 0 1 4005
box -2 -2 2 2
use M2_M1  M2_M1_11510
timestamp 1745462530
transform 1 0 2156 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_11511
timestamp 1745462530
transform 1 0 2892 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_11512
timestamp 1745462530
transform 1 0 2812 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_11513
timestamp 1745462530
transform 1 0 2780 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_11514
timestamp 1745462530
transform 1 0 3180 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_11515
timestamp 1745462530
transform 1 0 3076 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_11516
timestamp 1745462530
transform 1 0 3036 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_11517
timestamp 1745462530
transform 1 0 3620 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_11518
timestamp 1745462530
transform 1 0 3580 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_11519
timestamp 1745462530
transform 1 0 3564 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_11520
timestamp 1745462530
transform 1 0 3492 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_11521
timestamp 1745462530
transform 1 0 3476 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_11522
timestamp 1745462530
transform 1 0 3716 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_11523
timestamp 1745462530
transform 1 0 3644 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_11524
timestamp 1745462530
transform 1 0 3588 0 1 4005
box -2 -2 2 2
use M2_M1  M2_M1_11525
timestamp 1745462530
transform 1 0 3324 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_11526
timestamp 1745462530
transform 1 0 3308 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_11527
timestamp 1745462530
transform 1 0 3276 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_11528
timestamp 1745462530
transform 1 0 2428 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_11529
timestamp 1745462530
transform 1 0 2380 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_11530
timestamp 1745462530
transform 1 0 2164 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_11531
timestamp 1745462530
transform 1 0 2156 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_11532
timestamp 1745462530
transform 1 0 2116 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_11533
timestamp 1745462530
transform 1 0 2020 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_11534
timestamp 1745462530
transform 1 0 2804 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_11535
timestamp 1745462530
transform 1 0 2684 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_11536
timestamp 1745462530
transform 1 0 2676 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_11537
timestamp 1745462530
transform 1 0 2996 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_11538
timestamp 1745462530
transform 1 0 2996 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_11539
timestamp 1745462530
transform 1 0 2996 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_11540
timestamp 1745462530
transform 1 0 3924 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_11541
timestamp 1745462530
transform 1 0 3812 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_11542
timestamp 1745462530
transform 1 0 3804 0 1 4005
box -2 -2 2 2
use M2_M1  M2_M1_11543
timestamp 1745462530
transform 1 0 4004 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_11544
timestamp 1745462530
transform 1 0 3900 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_11545
timestamp 1745462530
transform 1 0 3860 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_11546
timestamp 1745462530
transform 1 0 3844 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_11547
timestamp 1745462530
transform 1 0 3772 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_11548
timestamp 1745462530
transform 1 0 3732 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_11549
timestamp 1745462530
transform 1 0 3820 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_11550
timestamp 1745462530
transform 1 0 3748 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_11551
timestamp 1745462530
transform 1 0 2524 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_11552
timestamp 1745462530
transform 1 0 2468 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_11553
timestamp 1745462530
transform 1 0 2300 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_11554
timestamp 1745462530
transform 1 0 2292 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_11555
timestamp 1745462530
transform 1 0 2268 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_11556
timestamp 1745462530
transform 1 0 2124 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_11557
timestamp 1745462530
transform 1 0 2636 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_11558
timestamp 1745462530
transform 1 0 2620 0 1 4195
box -2 -2 2 2
use M2_M1  M2_M1_11559
timestamp 1745462530
transform 1 0 2564 0 1 4005
box -2 -2 2 2
use M2_M1  M2_M1_11560
timestamp 1745462530
transform 1 0 2948 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_11561
timestamp 1745462530
transform 1 0 2916 0 1 4195
box -2 -2 2 2
use M2_M1  M2_M1_11562
timestamp 1745462530
transform 1 0 2900 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_11563
timestamp 1745462530
transform 1 0 4372 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_11564
timestamp 1745462530
transform 1 0 4356 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_11565
timestamp 1745462530
transform 1 0 4132 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_11566
timestamp 1745462530
transform 1 0 4124 0 1 3995
box -2 -2 2 2
use M2_M1  M2_M1_11567
timestamp 1745462530
transform 1 0 4364 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_11568
timestamp 1745462530
transform 1 0 4252 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_11569
timestamp 1745462530
transform 1 0 4108 0 1 4195
box -2 -2 2 2
use M2_M1  M2_M1_11570
timestamp 1745462530
transform 1 0 4108 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_11571
timestamp 1745462530
transform 1 0 4372 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_11572
timestamp 1745462530
transform 1 0 4268 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_11573
timestamp 1745462530
transform 1 0 4100 0 1 3945
box -2 -2 2 2
use M2_M1  M2_M1_11574
timestamp 1745462530
transform 1 0 4076 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_11575
timestamp 1745462530
transform 1 0 4012 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_11576
timestamp 1745462530
transform 1 0 4004 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_11577
timestamp 1745462530
transform 1 0 3924 0 1 4145
box -2 -2 2 2
use M2_M1  M2_M1_11578
timestamp 1745462530
transform 1 0 3908 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_11579
timestamp 1745462530
transform 1 0 1988 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_11580
timestamp 1745462530
transform 1 0 1948 0 1 4195
box -2 -2 2 2
use M2_M1  M2_M1_11581
timestamp 1745462530
transform 1 0 2076 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_11582
timestamp 1745462530
transform 1 0 2052 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_11583
timestamp 1745462530
transform 1 0 1900 0 1 4145
box -2 -2 2 2
use M2_M1  M2_M1_11584
timestamp 1745462530
transform 1 0 2660 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_11585
timestamp 1745462530
transform 1 0 2564 0 1 4195
box -2 -2 2 2
use M2_M1  M2_M1_11586
timestamp 1745462530
transform 1 0 2556 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_11587
timestamp 1745462530
transform 1 0 2996 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_11588
timestamp 1745462530
transform 1 0 2940 0 1 4195
box -2 -2 2 2
use M2_M1  M2_M1_11589
timestamp 1745462530
transform 1 0 2884 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_11590
timestamp 1745462530
transform 1 0 4244 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_11591
timestamp 1745462530
transform 1 0 4132 0 1 3945
box -2 -2 2 2
use M2_M1  M2_M1_11592
timestamp 1745462530
transform 1 0 4108 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_11593
timestamp 1745462530
transform 1 0 4100 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_11594
timestamp 1745462530
transform 1 0 4196 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_11595
timestamp 1745462530
transform 1 0 4092 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_11596
timestamp 1745462530
transform 1 0 4084 0 1 3995
box -2 -2 2 2
use M2_M1  M2_M1_11597
timestamp 1745462530
transform 1 0 4076 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_11598
timestamp 1745462530
transform 1 0 4068 0 1 3785
box -2 -2 2 2
use M2_M1  M2_M1_11599
timestamp 1745462530
transform 1 0 4364 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_11600
timestamp 1745462530
transform 1 0 4132 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_11601
timestamp 1745462530
transform 1 0 4076 0 1 3945
box -2 -2 2 2
use M2_M1  M2_M1_11602
timestamp 1745462530
transform 1 0 4036 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_11603
timestamp 1745462530
transform 1 0 4124 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_11604
timestamp 1745462530
transform 1 0 4004 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_11605
timestamp 1745462530
transform 1 0 3980 0 1 4145
box -2 -2 2 2
use M2_M1  M2_M1_11606
timestamp 1745462530
transform 1 0 3972 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_11607
timestamp 1745462530
transform 1 0 2020 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_11608
timestamp 1745462530
transform 1 0 1996 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_11609
timestamp 1745462530
transform 1 0 1972 0 1 4195
box -2 -2 2 2
use M2_M1  M2_M1_11610
timestamp 1745462530
transform 1 0 2020 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_11611
timestamp 1745462530
transform 1 0 1940 0 1 4005
box -2 -2 2 2
use M2_M1  M2_M1_11612
timestamp 1745462530
transform 1 0 1860 0 1 4195
box -2 -2 2 2
use M2_M1  M2_M1_11613
timestamp 1745462530
transform 1 0 1908 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_11614
timestamp 1745462530
transform 1 0 1844 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_11615
timestamp 1745462530
transform 1 0 1796 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_11616
timestamp 1745462530
transform 1 0 1828 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_11617
timestamp 1745462530
transform 1 0 1772 0 1 4005
box -2 -2 2 2
use M2_M1  M2_M1_11618
timestamp 1745462530
transform 1 0 1764 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_11619
timestamp 1745462530
transform 1 0 4372 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_11620
timestamp 1745462530
transform 1 0 4268 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_11621
timestamp 1745462530
transform 1 0 4260 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_11622
timestamp 1745462530
transform 1 0 4140 0 1 4005
box -2 -2 2 2
use M2_M1  M2_M1_11623
timestamp 1745462530
transform 1 0 4372 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_11624
timestamp 1745462530
transform 1 0 4260 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_11625
timestamp 1745462530
transform 1 0 4188 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_11626
timestamp 1745462530
transform 1 0 4180 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_11627
timestamp 1745462530
transform 1 0 4180 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_11628
timestamp 1745462530
transform 1 0 4180 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_11629
timestamp 1745462530
transform 1 0 4164 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_11630
timestamp 1745462530
transform 1 0 4076 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_11631
timestamp 1745462530
transform 1 0 4076 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_11632
timestamp 1745462530
transform 1 0 4060 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_11633
timestamp 1745462530
transform 1 0 4012 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_11634
timestamp 1745462530
transform 1 0 4004 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_11635
timestamp 1745462530
transform 1 0 1604 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_11636
timestamp 1745462530
transform 1 0 1516 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_11637
timestamp 1745462530
transform 1 0 1468 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_11638
timestamp 1745462530
transform 1 0 1460 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_11639
timestamp 1745462530
transform 1 0 1756 0 1 4005
box -2 -2 2 2
use M2_M1  M2_M1_11640
timestamp 1745462530
transform 1 0 1708 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_11641
timestamp 1745462530
transform 1 0 1636 0 1 4005
box -2 -2 2 2
use M2_M1  M2_M1_11642
timestamp 1745462530
transform 1 0 1580 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_11643
timestamp 1745462530
transform 1 0 1548 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_11644
timestamp 1745462530
transform 1 0 4364 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_11645
timestamp 1745462530
transform 1 0 4244 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_11646
timestamp 1745462530
transform 1 0 4228 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_11647
timestamp 1745462530
transform 1 0 4204 0 1 4005
box -2 -2 2 2
use M2_M1  M2_M1_11648
timestamp 1745462530
transform 1 0 4364 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_11649
timestamp 1745462530
transform 1 0 4260 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_11650
timestamp 1745462530
transform 1 0 4220 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_11651
timestamp 1745462530
transform 1 0 4132 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_11652
timestamp 1745462530
transform 1 0 4204 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_11653
timestamp 1745462530
transform 1 0 4196 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_11654
timestamp 1745462530
transform 1 0 4148 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_11655
timestamp 1745462530
transform 1 0 4092 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_11656
timestamp 1745462530
transform 1 0 4116 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_11657
timestamp 1745462530
transform 1 0 4020 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_11658
timestamp 1745462530
transform 1 0 3988 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_11659
timestamp 1745462530
transform 1 0 3876 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_11660
timestamp 1745462530
transform 1 0 1540 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_11661
timestamp 1745462530
transform 1 0 1524 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_11662
timestamp 1745462530
transform 1 0 1492 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_11663
timestamp 1745462530
transform 1 0 1548 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_11664
timestamp 1745462530
transform 1 0 1428 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_11665
timestamp 1745462530
transform 1 0 1420 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_11666
timestamp 1745462530
transform 1 0 692 0 1 4025
box -2 -2 2 2
use M2_M1  M2_M1_11667
timestamp 1745462530
transform 1 0 636 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_11668
timestamp 1745462530
transform 1 0 588 0 1 4025
box -2 -2 2 2
use M2_M1  M2_M1_11669
timestamp 1745462530
transform 1 0 564 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_11670
timestamp 1745462530
transform 1 0 540 0 1 4005
box -2 -2 2 2
use M2_M1  M2_M1_11671
timestamp 1745462530
transform 1 0 724 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_11672
timestamp 1745462530
transform 1 0 700 0 1 4035
box -2 -2 2 2
use M2_M1  M2_M1_11673
timestamp 1745462530
transform 1 0 596 0 1 4005
box -2 -2 2 2
use M2_M1  M2_M1_11674
timestamp 1745462530
transform 1 0 516 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_11675
timestamp 1745462530
transform 1 0 1236 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_11676
timestamp 1745462530
transform 1 0 1212 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_11677
timestamp 1745462530
transform 1 0 1164 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_11678
timestamp 1745462530
transform 1 0 460 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_11679
timestamp 1745462530
transform 1 0 108 0 1 4225
box -2 -2 2 2
use M2_M1  M2_M1_11680
timestamp 1745462530
transform 1 0 108 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_11681
timestamp 1745462530
transform 1 0 1300 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_11682
timestamp 1745462530
transform 1 0 1196 0 1 3825
box -2 -2 2 2
use M2_M1  M2_M1_11683
timestamp 1745462530
transform 1 0 476 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_11684
timestamp 1745462530
transform 1 0 468 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_11685
timestamp 1745462530
transform 1 0 428 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_11686
timestamp 1745462530
transform 1 0 212 0 1 3985
box -2 -2 2 2
use M2_M1  M2_M1_11687
timestamp 1745462530
transform 1 0 484 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_11688
timestamp 1745462530
transform 1 0 340 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_11689
timestamp 1745462530
transform 1 0 340 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_11690
timestamp 1745462530
transform 1 0 468 0 1 4145
box -2 -2 2 2
use M2_M1  M2_M1_11691
timestamp 1745462530
transform 1 0 452 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_11692
timestamp 1745462530
transform 1 0 452 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_11693
timestamp 1745462530
transform 1 0 964 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_11694
timestamp 1745462530
transform 1 0 956 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_11695
timestamp 1745462530
transform 1 0 588 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_11696
timestamp 1745462530
transform 1 0 1076 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_11697
timestamp 1745462530
transform 1 0 460 0 1 4005
box -2 -2 2 2
use M2_M1  M2_M1_11698
timestamp 1745462530
transform 1 0 340 0 1 4005
box -2 -2 2 2
use M2_M1  M2_M1_11699
timestamp 1745462530
transform 1 0 900 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_11700
timestamp 1745462530
transform 1 0 900 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_11701
timestamp 1745462530
transform 1 0 828 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_11702
timestamp 1745462530
transform 1 0 788 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_11703
timestamp 1745462530
transform 1 0 1732 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_11704
timestamp 1745462530
transform 1 0 1636 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_11705
timestamp 1745462530
transform 1 0 4380 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_11706
timestamp 1745462530
transform 1 0 4364 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_11707
timestamp 1745462530
transform 1 0 4364 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_11708
timestamp 1745462530
transform 1 0 4260 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_11709
timestamp 1745462530
transform 1 0 1484 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_11710
timestamp 1745462530
transform 1 0 1388 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_11711
timestamp 1745462530
transform 1 0 1340 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_11712
timestamp 1745462530
transform 1 0 1196 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_11713
timestamp 1745462530
transform 1 0 1292 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_11714
timestamp 1745462530
transform 1 0 1100 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_11715
timestamp 1745462530
transform 1 0 1316 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_11716
timestamp 1745462530
transform 1 0 1196 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_11717
timestamp 1745462530
transform 1 0 1020 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_11718
timestamp 1745462530
transform 1 0 812 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_11719
timestamp 1745462530
transform 1 0 252 0 1 4005
box -2 -2 2 2
use M2_M1  M2_M1_11720
timestamp 1745462530
transform 1 0 196 0 1 4145
box -2 -2 2 2
use M2_M1  M2_M1_11721
timestamp 1745462530
transform 1 0 116 0 1 4005
box -2 -2 2 2
use M2_M1  M2_M1_11722
timestamp 1745462530
transform 1 0 172 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_11723
timestamp 1745462530
transform 1 0 172 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_11724
timestamp 1745462530
transform 1 0 156 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_11725
timestamp 1745462530
transform 1 0 84 0 1 4025
box -2 -2 2 2
use M2_M1  M2_M1_11726
timestamp 1745462530
transform 1 0 172 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_11727
timestamp 1745462530
transform 1 0 156 0 1 4145
box -2 -2 2 2
use M2_M1  M2_M1_11728
timestamp 1745462530
transform 1 0 92 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_11729
timestamp 1745462530
transform 1 0 140 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_11730
timestamp 1745462530
transform 1 0 132 0 1 3995
box -2 -2 2 2
use M2_M1  M2_M1_11731
timestamp 1745462530
transform 1 0 124 0 1 4115
box -2 -2 2 2
use M2_M1  M2_M1_11732
timestamp 1745462530
transform 1 0 76 0 1 4145
box -2 -2 2 2
use M2_M1  M2_M1_11733
timestamp 1745462530
transform 1 0 540 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_11734
timestamp 1745462530
transform 1 0 532 0 1 3945
box -2 -2 2 2
use M2_M1  M2_M1_11735
timestamp 1745462530
transform 1 0 452 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_11736
timestamp 1745462530
transform 1 0 292 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_11737
timestamp 1745462530
transform 1 0 188 0 1 3795
box -2 -2 2 2
use M2_M1  M2_M1_11738
timestamp 1745462530
transform 1 0 2108 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_11739
timestamp 1745462530
transform 1 0 2036 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_11740
timestamp 1745462530
transform 1 0 2012 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_11741
timestamp 1745462530
transform 1 0 2012 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_11742
timestamp 1745462530
transform 1 0 1844 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_11743
timestamp 1745462530
transform 1 0 892 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_11744
timestamp 1745462530
transform 1 0 652 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_11745
timestamp 1745462530
transform 1 0 652 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_11746
timestamp 1745462530
transform 1 0 468 0 1 4205
box -2 -2 2 2
use M3_M2  M3_M2_0
timestamp 1745462530
transform 1 0 828 0 1 3145
box -3 -3 3 3
use M3_M2  M3_M2_1
timestamp 1745462530
transform 1 0 604 0 1 3145
box -3 -3 3 3
use M3_M2  M3_M2_2
timestamp 1745462530
transform 1 0 556 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_3
timestamp 1745462530
transform 1 0 452 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_4
timestamp 1745462530
transform 1 0 444 0 1 3005
box -3 -3 3 3
use M3_M2  M3_M2_5
timestamp 1745462530
transform 1 0 340 0 1 3005
box -3 -3 3 3
use M3_M2  M3_M2_6
timestamp 1745462530
transform 1 0 508 0 1 3105
box -3 -3 3 3
use M3_M2  M3_M2_7
timestamp 1745462530
transform 1 0 404 0 1 3105
box -3 -3 3 3
use M3_M2  M3_M2_8
timestamp 1745462530
transform 1 0 420 0 1 3085
box -3 -3 3 3
use M3_M2  M3_M2_9
timestamp 1745462530
transform 1 0 300 0 1 3085
box -3 -3 3 3
use M3_M2  M3_M2_10
timestamp 1745462530
transform 1 0 316 0 1 3025
box -3 -3 3 3
use M3_M2  M3_M2_11
timestamp 1745462530
transform 1 0 164 0 1 3025
box -3 -3 3 3
use M3_M2  M3_M2_12
timestamp 1745462530
transform 1 0 188 0 1 3015
box -3 -3 3 3
use M3_M2  M3_M2_13
timestamp 1745462530
transform 1 0 84 0 1 3015
box -3 -3 3 3
use M3_M2  M3_M2_14
timestamp 1745462530
transform 1 0 1660 0 1 3035
box -3 -3 3 3
use M3_M2  M3_M2_15
timestamp 1745462530
transform 1 0 1540 0 1 3325
box -3 -3 3 3
use M3_M2  M3_M2_16
timestamp 1745462530
transform 1 0 1508 0 1 3035
box -3 -3 3 3
use M3_M2  M3_M2_17
timestamp 1745462530
transform 1 0 1492 0 1 3325
box -3 -3 3 3
use M3_M2  M3_M2_18
timestamp 1745462530
transform 1 0 1444 0 1 3325
box -3 -3 3 3
use M3_M2  M3_M2_19
timestamp 1745462530
transform 1 0 1364 0 1 3325
box -3 -3 3 3
use M3_M2  M3_M2_20
timestamp 1745462530
transform 1 0 1276 0 1 3035
box -3 -3 3 3
use M3_M2  M3_M2_21
timestamp 1745462530
transform 1 0 1580 0 1 3285
box -3 -3 3 3
use M3_M2  M3_M2_22
timestamp 1745462530
transform 1 0 1532 0 1 3285
box -3 -3 3 3
use M3_M2  M3_M2_23
timestamp 1745462530
transform 1 0 1492 0 1 3285
box -3 -3 3 3
use M3_M2  M3_M2_24
timestamp 1745462530
transform 1 0 1492 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_25
timestamp 1745462530
transform 1 0 1436 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_26
timestamp 1745462530
transform 1 0 1996 0 1 3115
box -3 -3 3 3
use M3_M2  M3_M2_27
timestamp 1745462530
transform 1 0 1948 0 1 3115
box -3 -3 3 3
use M3_M2  M3_M2_28
timestamp 1745462530
transform 1 0 1716 0 1 3115
box -3 -3 3 3
use M3_M2  M3_M2_29
timestamp 1745462530
transform 1 0 1700 0 1 3195
box -3 -3 3 3
use M3_M2  M3_M2_30
timestamp 1745462530
transform 1 0 1540 0 1 3185
box -3 -3 3 3
use M3_M2  M3_M2_31
timestamp 1745462530
transform 1 0 1508 0 1 3355
box -3 -3 3 3
use M3_M2  M3_M2_32
timestamp 1745462530
transform 1 0 1428 0 1 3355
box -3 -3 3 3
use M3_M2  M3_M2_33
timestamp 1745462530
transform 1 0 1684 0 1 3575
box -3 -3 3 3
use M3_M2  M3_M2_34
timestamp 1745462530
transform 1 0 1644 0 1 3575
box -3 -3 3 3
use M3_M2  M3_M2_35
timestamp 1745462530
transform 1 0 1644 0 1 2935
box -3 -3 3 3
use M3_M2  M3_M2_36
timestamp 1745462530
transform 1 0 1572 0 1 2935
box -3 -3 3 3
use M3_M2  M3_M2_37
timestamp 1745462530
transform 1 0 1556 0 1 3255
box -3 -3 3 3
use M3_M2  M3_M2_38
timestamp 1745462530
transform 1 0 1556 0 1 3045
box -3 -3 3 3
use M3_M2  M3_M2_39
timestamp 1745462530
transform 1 0 1548 0 1 3575
box -3 -3 3 3
use M3_M2  M3_M2_40
timestamp 1745462530
transform 1 0 1492 0 1 3255
box -3 -3 3 3
use M3_M2  M3_M2_41
timestamp 1745462530
transform 1 0 1492 0 1 3045
box -3 -3 3 3
use M3_M2  M3_M2_42
timestamp 1745462530
transform 1 0 1372 0 1 3575
box -3 -3 3 3
use M3_M2  M3_M2_43
timestamp 1745462530
transform 1 0 1692 0 1 3615
box -3 -3 3 3
use M3_M2  M3_M2_44
timestamp 1745462530
transform 1 0 1628 0 1 3615
box -3 -3 3 3
use M3_M2  M3_M2_45
timestamp 1745462530
transform 1 0 1532 0 1 3615
box -3 -3 3 3
use M3_M2  M3_M2_46
timestamp 1745462530
transform 1 0 1396 0 1 3615
box -3 -3 3 3
use M3_M2  M3_M2_47
timestamp 1745462530
transform 1 0 1388 0 1 3445
box -3 -3 3 3
use M3_M2  M3_M2_48
timestamp 1745462530
transform 1 0 1388 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_49
timestamp 1745462530
transform 1 0 1244 0 1 3445
box -3 -3 3 3
use M3_M2  M3_M2_50
timestamp 1745462530
transform 1 0 1244 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_51
timestamp 1745462530
transform 1 0 1996 0 1 2965
box -3 -3 3 3
use M3_M2  M3_M2_52
timestamp 1745462530
transform 1 0 1988 0 1 3695
box -3 -3 3 3
use M3_M2  M3_M2_53
timestamp 1745462530
transform 1 0 1972 0 1 2965
box -3 -3 3 3
use M3_M2  M3_M2_54
timestamp 1745462530
transform 1 0 1940 0 1 3695
box -3 -3 3 3
use M3_M2  M3_M2_55
timestamp 1745462530
transform 1 0 1900 0 1 3695
box -3 -3 3 3
use M3_M2  M3_M2_56
timestamp 1745462530
transform 1 0 1892 0 1 2965
box -3 -3 3 3
use M3_M2  M3_M2_57
timestamp 1745462530
transform 1 0 1852 0 1 3695
box -3 -3 3 3
use M3_M2  M3_M2_58
timestamp 1745462530
transform 1 0 1804 0 1 3695
box -3 -3 3 3
use M3_M2  M3_M2_59
timestamp 1745462530
transform 1 0 1700 0 1 3695
box -3 -3 3 3
use M3_M2  M3_M2_60
timestamp 1745462530
transform 1 0 1612 0 1 3565
box -3 -3 3 3
use M3_M2  M3_M2_61
timestamp 1745462530
transform 1 0 1156 0 1 3595
box -3 -3 3 3
use M3_M2  M3_M2_62
timestamp 1745462530
transform 1 0 1156 0 1 3565
box -3 -3 3 3
use M3_M2  M3_M2_63
timestamp 1745462530
transform 1 0 940 0 1 3595
box -3 -3 3 3
use M3_M2  M3_M2_64
timestamp 1745462530
transform 1 0 1076 0 1 3625
box -3 -3 3 3
use M3_M2  M3_M2_65
timestamp 1745462530
transform 1 0 836 0 1 3625
box -3 -3 3 3
use M3_M2  M3_M2_66
timestamp 1745462530
transform 1 0 3124 0 1 3335
box -3 -3 3 3
use M3_M2  M3_M2_67
timestamp 1745462530
transform 1 0 3060 0 1 3335
box -3 -3 3 3
use M3_M2  M3_M2_68
timestamp 1745462530
transform 1 0 3044 0 1 3195
box -3 -3 3 3
use M3_M2  M3_M2_69
timestamp 1745462530
transform 1 0 2972 0 1 3235
box -3 -3 3 3
use M3_M2  M3_M2_70
timestamp 1745462530
transform 1 0 2972 0 1 3195
box -3 -3 3 3
use M3_M2  M3_M2_71
timestamp 1745462530
transform 1 0 2324 0 1 3235
box -3 -3 3 3
use M3_M2  M3_M2_72
timestamp 1745462530
transform 1 0 876 0 1 3235
box -3 -3 3 3
use M3_M2  M3_M2_73
timestamp 1745462530
transform 1 0 868 0 1 3385
box -3 -3 3 3
use M3_M2  M3_M2_74
timestamp 1745462530
transform 1 0 596 0 1 3385
box -3 -3 3 3
use M3_M2  M3_M2_75
timestamp 1745462530
transform 1 0 3172 0 1 3145
box -3 -3 3 3
use M3_M2  M3_M2_76
timestamp 1745462530
transform 1 0 3156 0 1 3275
box -3 -3 3 3
use M3_M2  M3_M2_77
timestamp 1745462530
transform 1 0 3156 0 1 3145
box -3 -3 3 3
use M3_M2  M3_M2_78
timestamp 1745462530
transform 1 0 3132 0 1 3275
box -3 -3 3 3
use M3_M2  M3_M2_79
timestamp 1745462530
transform 1 0 3028 0 1 3175
box -3 -3 3 3
use M3_M2  M3_M2_80
timestamp 1745462530
transform 1 0 3028 0 1 3145
box -3 -3 3 3
use M3_M2  M3_M2_81
timestamp 1745462530
transform 1 0 2948 0 1 3175
box -3 -3 3 3
use M3_M2  M3_M2_82
timestamp 1745462530
transform 1 0 2932 0 1 3275
box -3 -3 3 3
use M3_M2  M3_M2_83
timestamp 1745462530
transform 1 0 2316 0 1 3275
box -3 -3 3 3
use M3_M2  M3_M2_84
timestamp 1745462530
transform 1 0 996 0 1 3275
box -3 -3 3 3
use M3_M2  M3_M2_85
timestamp 1745462530
transform 1 0 988 0 1 3335
box -3 -3 3 3
use M3_M2  M3_M2_86
timestamp 1745462530
transform 1 0 700 0 1 3335
box -3 -3 3 3
use M3_M2  M3_M2_87
timestamp 1745462530
transform 1 0 3100 0 1 3275
box -3 -3 3 3
use M3_M2  M3_M2_88
timestamp 1745462530
transform 1 0 3068 0 1 3275
box -3 -3 3 3
use M3_M2  M3_M2_89
timestamp 1745462530
transform 1 0 2948 0 1 3275
box -3 -3 3 3
use M3_M2  M3_M2_90
timestamp 1745462530
transform 1 0 2916 0 1 3155
box -3 -3 3 3
use M3_M2  M3_M2_91
timestamp 1745462530
transform 1 0 2332 0 1 3155
box -3 -3 3 3
use M3_M2  M3_M2_92
timestamp 1745462530
transform 1 0 2268 0 1 3125
box -3 -3 3 3
use M3_M2  M3_M2_93
timestamp 1745462530
transform 1 0 1108 0 1 3295
box -3 -3 3 3
use M3_M2  M3_M2_94
timestamp 1745462530
transform 1 0 1108 0 1 3125
box -3 -3 3 3
use M3_M2  M3_M2_95
timestamp 1745462530
transform 1 0 924 0 1 3405
box -3 -3 3 3
use M3_M2  M3_M2_96
timestamp 1745462530
transform 1 0 924 0 1 3295
box -3 -3 3 3
use M3_M2  M3_M2_97
timestamp 1745462530
transform 1 0 588 0 1 3405
box -3 -3 3 3
use M3_M2  M3_M2_98
timestamp 1745462530
transform 1 0 2116 0 1 3545
box -3 -3 3 3
use M3_M2  M3_M2_99
timestamp 1745462530
transform 1 0 2108 0 1 3355
box -3 -3 3 3
use M3_M2  M3_M2_100
timestamp 1745462530
transform 1 0 2076 0 1 3545
box -3 -3 3 3
use M3_M2  M3_M2_101
timestamp 1745462530
transform 1 0 2076 0 1 3355
box -3 -3 3 3
use M3_M2  M3_M2_102
timestamp 1745462530
transform 1 0 1100 0 1 3545
box -3 -3 3 3
use M3_M2  M3_M2_103
timestamp 1745462530
transform 1 0 1100 0 1 3515
box -3 -3 3 3
use M3_M2  M3_M2_104
timestamp 1745462530
transform 1 0 876 0 1 3515
box -3 -3 3 3
use M3_M2  M3_M2_105
timestamp 1745462530
transform 1 0 676 0 1 3515
box -3 -3 3 3
use M3_M2  M3_M2_106
timestamp 1745462530
transform 1 0 2284 0 1 3265
box -3 -3 3 3
use M3_M2  M3_M2_107
timestamp 1745462530
transform 1 0 2236 0 1 3265
box -3 -3 3 3
use M3_M2  M3_M2_108
timestamp 1745462530
transform 1 0 2140 0 1 3325
box -3 -3 3 3
use M3_M2  M3_M2_109
timestamp 1745462530
transform 1 0 2140 0 1 3265
box -3 -3 3 3
use M3_M2  M3_M2_110
timestamp 1745462530
transform 1 0 2124 0 1 3485
box -3 -3 3 3
use M3_M2  M3_M2_111
timestamp 1745462530
transform 1 0 2084 0 1 3325
box -3 -3 3 3
use M3_M2  M3_M2_112
timestamp 1745462530
transform 1 0 2068 0 1 3475
box -3 -3 3 3
use M3_M2  M3_M2_113
timestamp 1745462530
transform 1 0 2012 0 1 3325
box -3 -3 3 3
use M3_M2  M3_M2_114
timestamp 1745462530
transform 1 0 932 0 1 3545
box -3 -3 3 3
use M3_M2  M3_M2_115
timestamp 1745462530
transform 1 0 932 0 1 3475
box -3 -3 3 3
use M3_M2  M3_M2_116
timestamp 1745462530
transform 1 0 716 0 1 3545
box -3 -3 3 3
use M3_M2  M3_M2_117
timestamp 1745462530
transform 1 0 2276 0 1 3255
box -3 -3 3 3
use M3_M2  M3_M2_118
timestamp 1745462530
transform 1 0 2228 0 1 3255
box -3 -3 3 3
use M3_M2  M3_M2_119
timestamp 1745462530
transform 1 0 2228 0 1 3195
box -3 -3 3 3
use M3_M2  M3_M2_120
timestamp 1745462530
transform 1 0 2220 0 1 3555
box -3 -3 3 3
use M3_M2  M3_M2_121
timestamp 1745462530
transform 1 0 2180 0 1 3195
box -3 -3 3 3
use M3_M2  M3_M2_122
timestamp 1745462530
transform 1 0 2084 0 1 3575
box -3 -3 3 3
use M3_M2  M3_M2_123
timestamp 1745462530
transform 1 0 2084 0 1 3555
box -3 -3 3 3
use M3_M2  M3_M2_124
timestamp 1745462530
transform 1 0 2060 0 1 3455
box -3 -3 3 3
use M3_M2  M3_M2_125
timestamp 1745462530
transform 1 0 2036 0 1 3575
box -3 -3 3 3
use M3_M2  M3_M2_126
timestamp 1745462530
transform 1 0 2036 0 1 3455
box -3 -3 3 3
use M3_M2  M3_M2_127
timestamp 1745462530
transform 1 0 1148 0 1 3525
box -3 -3 3 3
use M3_M2  M3_M2_128
timestamp 1745462530
transform 1 0 1148 0 1 3455
box -3 -3 3 3
use M3_M2  M3_M2_129
timestamp 1745462530
transform 1 0 532 0 1 3525
box -3 -3 3 3
use M3_M2  M3_M2_130
timestamp 1745462530
transform 1 0 1684 0 1 3345
box -3 -3 3 3
use M3_M2  M3_M2_131
timestamp 1745462530
transform 1 0 1644 0 1 3345
box -3 -3 3 3
use M3_M2  M3_M2_132
timestamp 1745462530
transform 1 0 1572 0 1 3345
box -3 -3 3 3
use M3_M2  M3_M2_133
timestamp 1745462530
transform 1 0 1252 0 1 3415
box -3 -3 3 3
use M3_M2  M3_M2_134
timestamp 1745462530
transform 1 0 1252 0 1 3345
box -3 -3 3 3
use M3_M2  M3_M2_135
timestamp 1745462530
transform 1 0 1156 0 1 3415
box -3 -3 3 3
use M3_M2  M3_M2_136
timestamp 1745462530
transform 1 0 1764 0 1 3265
box -3 -3 3 3
use M3_M2  M3_M2_137
timestamp 1745462530
transform 1 0 1708 0 1 3425
box -3 -3 3 3
use M3_M2  M3_M2_138
timestamp 1745462530
transform 1 0 1708 0 1 3265
box -3 -3 3 3
use M3_M2  M3_M2_139
timestamp 1745462530
transform 1 0 1668 0 1 3425
box -3 -3 3 3
use M3_M2  M3_M2_140
timestamp 1745462530
transform 1 0 1636 0 1 3265
box -3 -3 3 3
use M3_M2  M3_M2_141
timestamp 1745462530
transform 1 0 1636 0 1 3215
box -3 -3 3 3
use M3_M2  M3_M2_142
timestamp 1745462530
transform 1 0 1372 0 1 3375
box -3 -3 3 3
use M3_M2  M3_M2_143
timestamp 1745462530
transform 1 0 1300 0 1 3375
box -3 -3 3 3
use M3_M2  M3_M2_144
timestamp 1745462530
transform 1 0 1284 0 1 3215
box -3 -3 3 3
use M3_M2  M3_M2_145
timestamp 1745462530
transform 1 0 1700 0 1 3295
box -3 -3 3 3
use M3_M2  M3_M2_146
timestamp 1745462530
transform 1 0 1668 0 1 3385
box -3 -3 3 3
use M3_M2  M3_M2_147
timestamp 1745462530
transform 1 0 1636 0 1 3305
box -3 -3 3 3
use M3_M2  M3_M2_148
timestamp 1745462530
transform 1 0 1596 0 1 3385
box -3 -3 3 3
use M3_M2  M3_M2_149
timestamp 1745462530
transform 1 0 1596 0 1 3305
box -3 -3 3 3
use M3_M2  M3_M2_150
timestamp 1745462530
transform 1 0 1260 0 1 3405
box -3 -3 3 3
use M3_M2  M3_M2_151
timestamp 1745462530
transform 1 0 1260 0 1 3385
box -3 -3 3 3
use M3_M2  M3_M2_152
timestamp 1745462530
transform 1 0 1060 0 1 3405
box -3 -3 3 3
use M3_M2  M3_M2_153
timestamp 1745462530
transform 1 0 1772 0 1 3385
box -3 -3 3 3
use M3_M2  M3_M2_154
timestamp 1745462530
transform 1 0 1732 0 1 3635
box -3 -3 3 3
use M3_M2  M3_M2_155
timestamp 1745462530
transform 1 0 1732 0 1 3505
box -3 -3 3 3
use M3_M2  M3_M2_156
timestamp 1745462530
transform 1 0 1732 0 1 3385
box -3 -3 3 3
use M3_M2  M3_M2_157
timestamp 1745462530
transform 1 0 1660 0 1 3635
box -3 -3 3 3
use M3_M2  M3_M2_158
timestamp 1745462530
transform 1 0 1652 0 1 3505
box -3 -3 3 3
use M3_M2  M3_M2_159
timestamp 1745462530
transform 1 0 1380 0 1 3535
box -3 -3 3 3
use M3_M2  M3_M2_160
timestamp 1745462530
transform 1 0 1380 0 1 3505
box -3 -3 3 3
use M3_M2  M3_M2_161
timestamp 1745462530
transform 1 0 1356 0 1 3575
box -3 -3 3 3
use M3_M2  M3_M2_162
timestamp 1745462530
transform 1 0 1356 0 1 3535
box -3 -3 3 3
use M3_M2  M3_M2_163
timestamp 1745462530
transform 1 0 1028 0 1 3575
box -3 -3 3 3
use M3_M2  M3_M2_164
timestamp 1745462530
transform 1 0 1612 0 1 3415
box -3 -3 3 3
use M3_M2  M3_M2_165
timestamp 1745462530
transform 1 0 1268 0 1 3415
box -3 -3 3 3
use M3_M2  M3_M2_166
timestamp 1745462530
transform 1 0 1244 0 1 3645
box -3 -3 3 3
use M3_M2  M3_M2_167
timestamp 1745462530
transform 1 0 1124 0 1 3625
box -3 -3 3 3
use M3_M2  M3_M2_168
timestamp 1745462530
transform 1 0 1876 0 1 3085
box -3 -3 3 3
use M3_M2  M3_M2_169
timestamp 1745462530
transform 1 0 1828 0 1 3085
box -3 -3 3 3
use M3_M2  M3_M2_170
timestamp 1745462530
transform 1 0 1820 0 1 3485
box -3 -3 3 3
use M3_M2  M3_M2_171
timestamp 1745462530
transform 1 0 1788 0 1 3485
box -3 -3 3 3
use M3_M2  M3_M2_172
timestamp 1745462530
transform 1 0 1748 0 1 3485
box -3 -3 3 3
use M3_M2  M3_M2_173
timestamp 1745462530
transform 1 0 1636 0 1 3485
box -3 -3 3 3
use M3_M2  M3_M2_174
timestamp 1745462530
transform 1 0 1620 0 1 3645
box -3 -3 3 3
use M3_M2  M3_M2_175
timestamp 1745462530
transform 1 0 1276 0 1 3645
box -3 -3 3 3
use M3_M2  M3_M2_176
timestamp 1745462530
transform 1 0 876 0 1 3155
box -3 -3 3 3
use M3_M2  M3_M2_177
timestamp 1745462530
transform 1 0 772 0 1 3165
box -3 -3 3 3
use M3_M2  M3_M2_178
timestamp 1745462530
transform 1 0 732 0 1 3165
box -3 -3 3 3
use M3_M2  M3_M2_179
timestamp 1745462530
transform 1 0 492 0 1 3165
box -3 -3 3 3
use M3_M2  M3_M2_180
timestamp 1745462530
transform 1 0 660 0 1 3155
box -3 -3 3 3
use M3_M2  M3_M2_181
timestamp 1745462530
transform 1 0 564 0 1 3155
box -3 -3 3 3
use M3_M2  M3_M2_182
timestamp 1745462530
transform 1 0 484 0 1 3155
box -3 -3 3 3
use M3_M2  M3_M2_183
timestamp 1745462530
transform 1 0 620 0 1 3025
box -3 -3 3 3
use M3_M2  M3_M2_184
timestamp 1745462530
transform 1 0 524 0 1 3205
box -3 -3 3 3
use M3_M2  M3_M2_185
timestamp 1745462530
transform 1 0 524 0 1 3025
box -3 -3 3 3
use M3_M2  M3_M2_186
timestamp 1745462530
transform 1 0 476 0 1 3205
box -3 -3 3 3
use M3_M2  M3_M2_187
timestamp 1745462530
transform 1 0 396 0 1 3205
box -3 -3 3 3
use M3_M2  M3_M2_188
timestamp 1745462530
transform 1 0 516 0 1 2985
box -3 -3 3 3
use M3_M2  M3_M2_189
timestamp 1745462530
transform 1 0 420 0 1 2985
box -3 -3 3 3
use M3_M2  M3_M2_190
timestamp 1745462530
transform 1 0 380 0 1 3195
box -3 -3 3 3
use M3_M2  M3_M2_191
timestamp 1745462530
transform 1 0 284 0 1 3195
box -3 -3 3 3
use M3_M2  M3_M2_192
timestamp 1745462530
transform 1 0 412 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_193
timestamp 1745462530
transform 1 0 316 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_194
timestamp 1745462530
transform 1 0 308 0 1 3105
box -3 -3 3 3
use M3_M2  M3_M2_195
timestamp 1745462530
transform 1 0 268 0 1 3105
box -3 -3 3 3
use M3_M2  M3_M2_196
timestamp 1745462530
transform 1 0 180 0 1 3105
box -3 -3 3 3
use M3_M2  M3_M2_197
timestamp 1745462530
transform 1 0 268 0 1 3205
box -3 -3 3 3
use M3_M2  M3_M2_198
timestamp 1745462530
transform 1 0 228 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_199
timestamp 1745462530
transform 1 0 172 0 1 3205
box -3 -3 3 3
use M3_M2  M3_M2_200
timestamp 1745462530
transform 1 0 148 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_201
timestamp 1745462530
transform 1 0 2508 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_202
timestamp 1745462530
transform 1 0 2508 0 1 2385
box -3 -3 3 3
use M3_M2  M3_M2_203
timestamp 1745462530
transform 1 0 2484 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_204
timestamp 1745462530
transform 1 0 2452 0 1 2385
box -3 -3 3 3
use M3_M2  M3_M2_205
timestamp 1745462530
transform 1 0 2444 0 1 2285
box -3 -3 3 3
use M3_M2  M3_M2_206
timestamp 1745462530
transform 1 0 2356 0 1 2285
box -3 -3 3 3
use M3_M2  M3_M2_207
timestamp 1745462530
transform 1 0 2348 0 1 2435
box -3 -3 3 3
use M3_M2  M3_M2_208
timestamp 1745462530
transform 1 0 2324 0 1 2435
box -3 -3 3 3
use M3_M2  M3_M2_209
timestamp 1745462530
transform 1 0 2300 0 1 2285
box -3 -3 3 3
use M3_M2  M3_M2_210
timestamp 1745462530
transform 1 0 2444 0 1 2775
box -3 -3 3 3
use M3_M2  M3_M2_211
timestamp 1745462530
transform 1 0 2380 0 1 2455
box -3 -3 3 3
use M3_M2  M3_M2_212
timestamp 1745462530
transform 1 0 2356 0 1 2455
box -3 -3 3 3
use M3_M2  M3_M2_213
timestamp 1745462530
transform 1 0 2340 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_214
timestamp 1745462530
transform 1 0 2332 0 1 2775
box -3 -3 3 3
use M3_M2  M3_M2_215
timestamp 1745462530
transform 1 0 2316 0 1 2455
box -3 -3 3 3
use M3_M2  M3_M2_216
timestamp 1745462530
transform 1 0 2284 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_217
timestamp 1745462530
transform 1 0 2372 0 1 2275
box -3 -3 3 3
use M3_M2  M3_M2_218
timestamp 1745462530
transform 1 0 2364 0 1 2865
box -3 -3 3 3
use M3_M2  M3_M2_219
timestamp 1745462530
transform 1 0 2348 0 1 2725
box -3 -3 3 3
use M3_M2  M3_M2_220
timestamp 1745462530
transform 1 0 2332 0 1 2725
box -3 -3 3 3
use M3_M2  M3_M2_221
timestamp 1745462530
transform 1 0 2332 0 1 2615
box -3 -3 3 3
use M3_M2  M3_M2_222
timestamp 1745462530
transform 1 0 2316 0 1 2275
box -3 -3 3 3
use M3_M2  M3_M2_223
timestamp 1745462530
transform 1 0 2308 0 1 2615
box -3 -3 3 3
use M3_M2  M3_M2_224
timestamp 1745462530
transform 1 0 2300 0 1 2865
box -3 -3 3 3
use M3_M2  M3_M2_225
timestamp 1745462530
transform 1 0 2300 0 1 2725
box -3 -3 3 3
use M3_M2  M3_M2_226
timestamp 1745462530
transform 1 0 2292 0 1 2275
box -3 -3 3 3
use M3_M2  M3_M2_227
timestamp 1745462530
transform 1 0 2276 0 1 2775
box -3 -3 3 3
use M3_M2  M3_M2_228
timestamp 1745462530
transform 1 0 2244 0 1 2265
box -3 -3 3 3
use M3_M2  M3_M2_229
timestamp 1745462530
transform 1 0 2228 0 1 2775
box -3 -3 3 3
use M3_M2  M3_M2_230
timestamp 1745462530
transform 1 0 2220 0 1 2175
box -3 -3 3 3
use M3_M2  M3_M2_231
timestamp 1745462530
transform 1 0 2212 0 1 2265
box -3 -3 3 3
use M3_M2  M3_M2_232
timestamp 1745462530
transform 1 0 2140 0 1 2175
box -3 -3 3 3
use M3_M2  M3_M2_233
timestamp 1745462530
transform 1 0 2092 0 1 2175
box -3 -3 3 3
use M3_M2  M3_M2_234
timestamp 1745462530
transform 1 0 2276 0 1 2085
box -3 -3 3 3
use M3_M2  M3_M2_235
timestamp 1745462530
transform 1 0 2260 0 1 2365
box -3 -3 3 3
use M3_M2  M3_M2_236
timestamp 1745462530
transform 1 0 2236 0 1 2095
box -3 -3 3 3
use M3_M2  M3_M2_237
timestamp 1745462530
transform 1 0 2236 0 1 2085
box -3 -3 3 3
use M3_M2  M3_M2_238
timestamp 1745462530
transform 1 0 2188 0 1 2725
box -3 -3 3 3
use M3_M2  M3_M2_239
timestamp 1745462530
transform 1 0 2180 0 1 2565
box -3 -3 3 3
use M3_M2  M3_M2_240
timestamp 1745462530
transform 1 0 2180 0 1 2365
box -3 -3 3 3
use M3_M2  M3_M2_241
timestamp 1745462530
transform 1 0 2140 0 1 2095
box -3 -3 3 3
use M3_M2  M3_M2_242
timestamp 1745462530
transform 1 0 2108 0 1 2095
box -3 -3 3 3
use M3_M2  M3_M2_243
timestamp 1745462530
transform 1 0 2100 0 1 2725
box -3 -3 3 3
use M3_M2  M3_M2_244
timestamp 1745462530
transform 1 0 2100 0 1 2565
box -3 -3 3 3
use M3_M2  M3_M2_245
timestamp 1745462530
transform 1 0 2300 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_246
timestamp 1745462530
transform 1 0 2276 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_247
timestamp 1745462530
transform 1 0 2228 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_248
timestamp 1745462530
transform 1 0 2196 0 1 2475
box -3 -3 3 3
use M3_M2  M3_M2_249
timestamp 1745462530
transform 1 0 2196 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_250
timestamp 1745462530
transform 1 0 2180 0 1 2615
box -3 -3 3 3
use M3_M2  M3_M2_251
timestamp 1745462530
transform 1 0 2108 0 1 2615
box -3 -3 3 3
use M3_M2  M3_M2_252
timestamp 1745462530
transform 1 0 2108 0 1 2475
box -3 -3 3 3
use M3_M2  M3_M2_253
timestamp 1745462530
transform 1 0 1164 0 1 3555
box -3 -3 3 3
use M3_M2  M3_M2_254
timestamp 1745462530
transform 1 0 1140 0 1 3555
box -3 -3 3 3
use M3_M2  M3_M2_255
timestamp 1745462530
transform 1 0 372 0 1 3935
box -3 -3 3 3
use M3_M2  M3_M2_256
timestamp 1745462530
transform 1 0 300 0 1 3935
box -3 -3 3 3
use M3_M2  M3_M2_257
timestamp 1745462530
transform 1 0 788 0 1 3795
box -3 -3 3 3
use M3_M2  M3_M2_258
timestamp 1745462530
transform 1 0 732 0 1 3795
box -3 -3 3 3
use M3_M2  M3_M2_259
timestamp 1745462530
transform 1 0 604 0 1 3795
box -3 -3 3 3
use M3_M2  M3_M2_260
timestamp 1745462530
transform 1 0 780 0 1 3905
box -3 -3 3 3
use M3_M2  M3_M2_261
timestamp 1745462530
transform 1 0 764 0 1 3905
box -3 -3 3 3
use M3_M2  M3_M2_262
timestamp 1745462530
transform 1 0 668 0 1 3905
box -3 -3 3 3
use M3_M2  M3_M2_263
timestamp 1745462530
transform 1 0 2228 0 1 2665
box -3 -3 3 3
use M3_M2  M3_M2_264
timestamp 1745462530
transform 1 0 2228 0 1 2565
box -3 -3 3 3
use M3_M2  M3_M2_265
timestamp 1745462530
transform 1 0 2212 0 1 2665
box -3 -3 3 3
use M3_M2  M3_M2_266
timestamp 1745462530
transform 1 0 2204 0 1 2565
box -3 -3 3 3
use M3_M2  M3_M2_267
timestamp 1745462530
transform 1 0 2364 0 1 2565
box -3 -3 3 3
use M3_M2  M3_M2_268
timestamp 1745462530
transform 1 0 2284 0 1 2615
box -3 -3 3 3
use M3_M2  M3_M2_269
timestamp 1745462530
transform 1 0 2284 0 1 2565
box -3 -3 3 3
use M3_M2  M3_M2_270
timestamp 1745462530
transform 1 0 2196 0 1 2615
box -3 -3 3 3
use M3_M2  M3_M2_271
timestamp 1745462530
transform 1 0 2436 0 1 2535
box -3 -3 3 3
use M3_M2  M3_M2_272
timestamp 1745462530
transform 1 0 2380 0 1 2535
box -3 -3 3 3
use M3_M2  M3_M2_273
timestamp 1745462530
transform 1 0 388 0 1 3525
box -3 -3 3 3
use M3_M2  M3_M2_274
timestamp 1745462530
transform 1 0 372 0 1 3525
box -3 -3 3 3
use M3_M2  M3_M2_275
timestamp 1745462530
transform 1 0 300 0 1 3545
box -3 -3 3 3
use M3_M2  M3_M2_276
timestamp 1745462530
transform 1 0 268 0 1 3545
box -3 -3 3 3
use M3_M2  M3_M2_277
timestamp 1745462530
transform 1 0 316 0 1 3585
box -3 -3 3 3
use M3_M2  M3_M2_278
timestamp 1745462530
transform 1 0 236 0 1 3585
box -3 -3 3 3
use M3_M2  M3_M2_279
timestamp 1745462530
transform 1 0 356 0 1 3625
box -3 -3 3 3
use M3_M2  M3_M2_280
timestamp 1745462530
transform 1 0 292 0 1 3625
box -3 -3 3 3
use M3_M2  M3_M2_281
timestamp 1745462530
transform 1 0 188 0 1 3465
box -3 -3 3 3
use M3_M2  M3_M2_282
timestamp 1745462530
transform 1 0 132 0 1 3465
box -3 -3 3 3
use M3_M2  M3_M2_283
timestamp 1745462530
transform 1 0 1588 0 1 3055
box -3 -3 3 3
use M3_M2  M3_M2_284
timestamp 1745462530
transform 1 0 1220 0 1 3055
box -3 -3 3 3
use M3_M2  M3_M2_285
timestamp 1745462530
transform 1 0 1204 0 1 3255
box -3 -3 3 3
use M3_M2  M3_M2_286
timestamp 1745462530
transform 1 0 1196 0 1 3515
box -3 -3 3 3
use M3_M2  M3_M2_287
timestamp 1745462530
transform 1 0 1116 0 1 3515
box -3 -3 3 3
use M3_M2  M3_M2_288
timestamp 1745462530
transform 1 0 1092 0 1 3255
box -3 -3 3 3
use M3_M2  M3_M2_289
timestamp 1745462530
transform 1 0 2188 0 1 2965
box -3 -3 3 3
use M3_M2  M3_M2_290
timestamp 1745462530
transform 1 0 2124 0 1 2965
box -3 -3 3 3
use M3_M2  M3_M2_291
timestamp 1745462530
transform 1 0 2084 0 1 2965
box -3 -3 3 3
use M3_M2  M3_M2_292
timestamp 1745462530
transform 1 0 2068 0 1 3395
box -3 -3 3 3
use M3_M2  M3_M2_293
timestamp 1745462530
transform 1 0 1020 0 1 3355
box -3 -3 3 3
use M3_M2  M3_M2_294
timestamp 1745462530
transform 1 0 972 0 1 3395
box -3 -3 3 3
use M3_M2  M3_M2_295
timestamp 1745462530
transform 1 0 972 0 1 3355
box -3 -3 3 3
use M3_M2  M3_M2_296
timestamp 1745462530
transform 1 0 2340 0 1 3365
box -3 -3 3 3
use M3_M2  M3_M2_297
timestamp 1745462530
transform 1 0 2276 0 1 3355
box -3 -3 3 3
use M3_M2  M3_M2_298
timestamp 1745462530
transform 1 0 2228 0 1 3355
box -3 -3 3 3
use M3_M2  M3_M2_299
timestamp 1745462530
transform 1 0 2204 0 1 3355
box -3 -3 3 3
use M3_M2  M3_M2_300
timestamp 1745462530
transform 1 0 2316 0 1 3395
box -3 -3 3 3
use M3_M2  M3_M2_301
timestamp 1745462530
transform 1 0 2268 0 1 3395
box -3 -3 3 3
use M3_M2  M3_M2_302
timestamp 1745462530
transform 1 0 2204 0 1 3395
box -3 -3 3 3
use M3_M2  M3_M2_303
timestamp 1745462530
transform 1 0 2116 0 1 3395
box -3 -3 3 3
use M3_M2  M3_M2_304
timestamp 1745462530
transform 1 0 2236 0 1 3425
box -3 -3 3 3
use M3_M2  M3_M2_305
timestamp 1745462530
transform 1 0 2132 0 1 3455
box -3 -3 3 3
use M3_M2  M3_M2_306
timestamp 1745462530
transform 1 0 2084 0 1 3455
box -3 -3 3 3
use M3_M2  M3_M2_307
timestamp 1745462530
transform 1 0 2084 0 1 3425
box -3 -3 3 3
use M3_M2  M3_M2_308
timestamp 1745462530
transform 1 0 3140 0 1 3315
box -3 -3 3 3
use M3_M2  M3_M2_309
timestamp 1745462530
transform 1 0 3052 0 1 3315
box -3 -3 3 3
use M3_M2  M3_M2_310
timestamp 1745462530
transform 1 0 3132 0 1 3255
box -3 -3 3 3
use M3_M2  M3_M2_311
timestamp 1745462530
transform 1 0 3108 0 1 3255
box -3 -3 3 3
use M3_M2  M3_M2_312
timestamp 1745462530
transform 1 0 3004 0 1 3255
box -3 -3 3 3
use M3_M2  M3_M2_313
timestamp 1745462530
transform 1 0 1684 0 1 3085
box -3 -3 3 3
use M3_M2  M3_M2_314
timestamp 1745462530
transform 1 0 1596 0 1 3265
box -3 -3 3 3
use M3_M2  M3_M2_315
timestamp 1745462530
transform 1 0 1540 0 1 3305
box -3 -3 3 3
use M3_M2  M3_M2_316
timestamp 1745462530
transform 1 0 1540 0 1 3265
box -3 -3 3 3
use M3_M2  M3_M2_317
timestamp 1745462530
transform 1 0 1516 0 1 3075
box -3 -3 3 3
use M3_M2  M3_M2_318
timestamp 1745462530
transform 1 0 1484 0 1 3075
box -3 -3 3 3
use M3_M2  M3_M2_319
timestamp 1745462530
transform 1 0 1380 0 1 3315
box -3 -3 3 3
use M3_M2  M3_M2_320
timestamp 1745462530
transform 1 0 1380 0 1 3285
box -3 -3 3 3
use M3_M2  M3_M2_321
timestamp 1745462530
transform 1 0 1324 0 1 3285
box -3 -3 3 3
use M3_M2  M3_M2_322
timestamp 1745462530
transform 1 0 1308 0 1 3285
box -3 -3 3 3
use M3_M2  M3_M2_323
timestamp 1745462530
transform 1 0 1300 0 1 3075
box -3 -3 3 3
use M3_M2  M3_M2_324
timestamp 1745462530
transform 1 0 1772 0 1 3255
box -3 -3 3 3
use M3_M2  M3_M2_325
timestamp 1745462530
transform 1 0 1732 0 1 3255
box -3 -3 3 3
use M3_M2  M3_M2_326
timestamp 1745462530
transform 1 0 1684 0 1 3255
box -3 -3 3 3
use M3_M2  M3_M2_327
timestamp 1745462530
transform 1 0 1660 0 1 3255
box -3 -3 3 3
use M3_M2  M3_M2_328
timestamp 1745462530
transform 1 0 1572 0 1 3255
box -3 -3 3 3
use M3_M2  M3_M2_329
timestamp 1745462530
transform 1 0 1572 0 1 3085
box -3 -3 3 3
use M3_M2  M3_M2_330
timestamp 1745462530
transform 1 0 1340 0 1 3085
box -3 -3 3 3
use M3_M2  M3_M2_331
timestamp 1745462530
transform 1 0 1828 0 1 3605
box -3 -3 3 3
use M3_M2  M3_M2_332
timestamp 1745462530
transform 1 0 1748 0 1 3515
box -3 -3 3 3
use M3_M2  M3_M2_333
timestamp 1745462530
transform 1 0 1740 0 1 3605
box -3 -3 3 3
use M3_M2  M3_M2_334
timestamp 1745462530
transform 1 0 1700 0 1 3515
box -3 -3 3 3
use M3_M2  M3_M2_335
timestamp 1745462530
transform 1 0 1676 0 1 3515
box -3 -3 3 3
use M3_M2  M3_M2_336
timestamp 1745462530
transform 1 0 1644 0 1 3535
box -3 -3 3 3
use M3_M2  M3_M2_337
timestamp 1745462530
transform 1 0 1260 0 1 3525
box -3 -3 3 3
use M3_M2  M3_M2_338
timestamp 1745462530
transform 1 0 2164 0 1 2755
box -3 -3 3 3
use M3_M2  M3_M2_339
timestamp 1745462530
transform 1 0 2164 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_340
timestamp 1745462530
transform 1 0 2148 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_341
timestamp 1745462530
transform 1 0 2116 0 1 2755
box -3 -3 3 3
use M3_M2  M3_M2_342
timestamp 1745462530
transform 1 0 2100 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_343
timestamp 1745462530
transform 1 0 2444 0 1 2665
box -3 -3 3 3
use M3_M2  M3_M2_344
timestamp 1745462530
transform 1 0 2404 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_345
timestamp 1745462530
transform 1 0 2372 0 1 2755
box -3 -3 3 3
use M3_M2  M3_M2_346
timestamp 1745462530
transform 1 0 2372 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_347
timestamp 1745462530
transform 1 0 2364 0 1 2665
box -3 -3 3 3
use M3_M2  M3_M2_348
timestamp 1745462530
transform 1 0 2348 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_349
timestamp 1745462530
transform 1 0 2332 0 1 2665
box -3 -3 3 3
use M3_M2  M3_M2_350
timestamp 1745462530
transform 1 0 2332 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_351
timestamp 1745462530
transform 1 0 2300 0 1 2455
box -3 -3 3 3
use M3_M2  M3_M2_352
timestamp 1745462530
transform 1 0 2284 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_353
timestamp 1745462530
transform 1 0 2276 0 1 2455
box -3 -3 3 3
use M3_M2  M3_M2_354
timestamp 1745462530
transform 1 0 2268 0 1 2755
box -3 -3 3 3
use M3_M2  M3_M2_355
timestamp 1745462530
transform 1 0 2244 0 1 2665
box -3 -3 3 3
use M3_M2  M3_M2_356
timestamp 1745462530
transform 1 0 2236 0 1 2755
box -3 -3 3 3
use M3_M2  M3_M2_357
timestamp 1745462530
transform 1 0 2236 0 1 2455
box -3 -3 3 3
use M3_M2  M3_M2_358
timestamp 1745462530
transform 1 0 2212 0 1 3035
box -3 -3 3 3
use M3_M2  M3_M2_359
timestamp 1745462530
transform 1 0 2068 0 1 3035
box -3 -3 3 3
use M3_M2  M3_M2_360
timestamp 1745462530
transform 1 0 2308 0 1 2435
box -3 -3 3 3
use M3_M2  M3_M2_361
timestamp 1745462530
transform 1 0 2284 0 1 2545
box -3 -3 3 3
use M3_M2  M3_M2_362
timestamp 1745462530
transform 1 0 2252 0 1 2545
box -3 -3 3 3
use M3_M2  M3_M2_363
timestamp 1745462530
transform 1 0 2252 0 1 2435
box -3 -3 3 3
use M3_M2  M3_M2_364
timestamp 1745462530
transform 1 0 2484 0 1 2565
box -3 -3 3 3
use M3_M2  M3_M2_365
timestamp 1745462530
transform 1 0 2412 0 1 2565
box -3 -3 3 3
use M3_M2  M3_M2_366
timestamp 1745462530
transform 1 0 2660 0 1 2335
box -3 -3 3 3
use M3_M2  M3_M2_367
timestamp 1745462530
transform 1 0 2252 0 1 2335
box -3 -3 3 3
use M3_M2  M3_M2_368
timestamp 1745462530
transform 1 0 2228 0 1 2285
box -3 -3 3 3
use M3_M2  M3_M2_369
timestamp 1745462530
transform 1 0 2140 0 1 2285
box -3 -3 3 3
use M3_M2  M3_M2_370
timestamp 1745462530
transform 1 0 2596 0 1 2235
box -3 -3 3 3
use M3_M2  M3_M2_371
timestamp 1745462530
transform 1 0 2220 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_372
timestamp 1745462530
transform 1 0 2092 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_373
timestamp 1745462530
transform 1 0 3364 0 1 1435
box -3 -3 3 3
use M3_M2  M3_M2_374
timestamp 1745462530
transform 1 0 3316 0 1 605
box -3 -3 3 3
use M3_M2  M3_M2_375
timestamp 1745462530
transform 1 0 3148 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_376
timestamp 1745462530
transform 1 0 3148 0 1 1435
box -3 -3 3 3
use M3_M2  M3_M2_377
timestamp 1745462530
transform 1 0 3124 0 1 1575
box -3 -3 3 3
use M3_M2  M3_M2_378
timestamp 1745462530
transform 1 0 3124 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_379
timestamp 1745462530
transform 1 0 2580 0 1 1575
box -3 -3 3 3
use M3_M2  M3_M2_380
timestamp 1745462530
transform 1 0 2580 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_381
timestamp 1745462530
transform 1 0 2564 0 1 2425
box -3 -3 3 3
use M3_M2  M3_M2_382
timestamp 1745462530
transform 1 0 2516 0 1 1575
box -3 -3 3 3
use M3_M2  M3_M2_383
timestamp 1745462530
transform 1 0 2516 0 1 1485
box -3 -3 3 3
use M3_M2  M3_M2_384
timestamp 1745462530
transform 1 0 2484 0 1 605
box -3 -3 3 3
use M3_M2  M3_M2_385
timestamp 1745462530
transform 1 0 2484 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_386
timestamp 1745462530
transform 1 0 2308 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_387
timestamp 1745462530
transform 1 0 2300 0 1 1485
box -3 -3 3 3
use M3_M2  M3_M2_388
timestamp 1745462530
transform 1 0 2172 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_389
timestamp 1745462530
transform 1 0 2140 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_390
timestamp 1745462530
transform 1 0 1556 0 1 645
box -3 -3 3 3
use M3_M2  M3_M2_391
timestamp 1745462530
transform 1 0 1556 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_392
timestamp 1745462530
transform 1 0 1532 0 1 645
box -3 -3 3 3
use M3_M2  M3_M2_393
timestamp 1745462530
transform 1 0 852 0 1 2425
box -3 -3 3 3
use M3_M2  M3_M2_394
timestamp 1745462530
transform 1 0 828 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_395
timestamp 1745462530
transform 1 0 2340 0 1 2475
box -3 -3 3 3
use M3_M2  M3_M2_396
timestamp 1745462530
transform 1 0 2324 0 1 2895
box -3 -3 3 3
use M3_M2  M3_M2_397
timestamp 1745462530
transform 1 0 2316 0 1 2475
box -3 -3 3 3
use M3_M2  M3_M2_398
timestamp 1745462530
transform 1 0 2260 0 1 2475
box -3 -3 3 3
use M3_M2  M3_M2_399
timestamp 1745462530
transform 1 0 2228 0 1 2895
box -3 -3 3 3
use M3_M2  M3_M2_400
timestamp 1745462530
transform 1 0 3324 0 1 1415
box -3 -3 3 3
use M3_M2  M3_M2_401
timestamp 1745462530
transform 1 0 3292 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_402
timestamp 1745462530
transform 1 0 3284 0 1 1415
box -3 -3 3 3
use M3_M2  M3_M2_403
timestamp 1745462530
transform 1 0 2628 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_404
timestamp 1745462530
transform 1 0 2532 0 1 2325
box -3 -3 3 3
use M3_M2  M3_M2_405
timestamp 1745462530
transform 1 0 1652 0 1 675
box -3 -3 3 3
use M3_M2  M3_M2_406
timestamp 1745462530
transform 1 0 1652 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_407
timestamp 1745462530
transform 1 0 1596 0 1 675
box -3 -3 3 3
use M3_M2  M3_M2_408
timestamp 1745462530
transform 1 0 1556 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_409
timestamp 1745462530
transform 1 0 1556 0 1 675
box -3 -3 3 3
use M3_M2  M3_M2_410
timestamp 1745462530
transform 1 0 948 0 1 2325
box -3 -3 3 3
use M3_M2  M3_M2_411
timestamp 1745462530
transform 1 0 948 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_412
timestamp 1745462530
transform 1 0 948 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_413
timestamp 1745462530
transform 1 0 932 0 1 2015
box -3 -3 3 3
use M3_M2  M3_M2_414
timestamp 1745462530
transform 1 0 3324 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_415
timestamp 1745462530
transform 1 0 3236 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_416
timestamp 1745462530
transform 1 0 3228 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_417
timestamp 1745462530
transform 1 0 2676 0 1 655
box -3 -3 3 3
use M3_M2  M3_M2_418
timestamp 1745462530
transform 1 0 2676 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_419
timestamp 1745462530
transform 1 0 2220 0 1 2435
box -3 -3 3 3
use M3_M2  M3_M2_420
timestamp 1745462530
transform 1 0 2004 0 1 2435
box -3 -3 3 3
use M3_M2  M3_M2_421
timestamp 1745462530
transform 1 0 2004 0 1 2185
box -3 -3 3 3
use M3_M2  M3_M2_422
timestamp 1745462530
transform 1 0 2004 0 1 685
box -3 -3 3 3
use M3_M2  M3_M2_423
timestamp 1745462530
transform 1 0 1996 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_424
timestamp 1745462530
transform 1 0 1956 0 1 2185
box -3 -3 3 3
use M3_M2  M3_M2_425
timestamp 1745462530
transform 1 0 1956 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_426
timestamp 1745462530
transform 1 0 1596 0 1 685
box -3 -3 3 3
use M3_M2  M3_M2_427
timestamp 1745462530
transform 1 0 892 0 1 2435
box -3 -3 3 3
use M3_M2  M3_M2_428
timestamp 1745462530
transform 1 0 868 0 1 685
box -3 -3 3 3
use M3_M2  M3_M2_429
timestamp 1745462530
transform 1 0 3268 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_430
timestamp 1745462530
transform 1 0 3252 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_431
timestamp 1745462530
transform 1 0 2676 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_432
timestamp 1745462530
transform 1 0 2644 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_433
timestamp 1745462530
transform 1 0 2644 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_434
timestamp 1745462530
transform 1 0 2644 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_435
timestamp 1745462530
transform 1 0 2644 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_436
timestamp 1745462530
transform 1 0 2636 0 1 2475
box -3 -3 3 3
use M3_M2  M3_M2_437
timestamp 1745462530
transform 1 0 2628 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_438
timestamp 1745462530
transform 1 0 2564 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_439
timestamp 1745462530
transform 1 0 2556 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_440
timestamp 1745462530
transform 1 0 2548 0 1 2485
box -3 -3 3 3
use M3_M2  M3_M2_441
timestamp 1745462530
transform 1 0 2532 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_442
timestamp 1745462530
transform 1 0 2468 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_443
timestamp 1745462530
transform 1 0 2444 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_444
timestamp 1745462530
transform 1 0 1564 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_445
timestamp 1745462530
transform 1 0 940 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_446
timestamp 1745462530
transform 1 0 932 0 1 2485
box -3 -3 3 3
use M3_M2  M3_M2_447
timestamp 1745462530
transform 1 0 1308 0 1 2535
box -3 -3 3 3
use M3_M2  M3_M2_448
timestamp 1745462530
transform 1 0 1100 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_449
timestamp 1745462530
transform 1 0 2460 0 1 2985
box -3 -3 3 3
use M3_M2  M3_M2_450
timestamp 1745462530
transform 1 0 2436 0 1 2625
box -3 -3 3 3
use M3_M2  M3_M2_451
timestamp 1745462530
transform 1 0 2396 0 1 2625
box -3 -3 3 3
use M3_M2  M3_M2_452
timestamp 1745462530
transform 1 0 2172 0 1 2985
box -3 -3 3 3
use M3_M2  M3_M2_453
timestamp 1745462530
transform 1 0 2284 0 1 2125
box -3 -3 3 3
use M3_M2  M3_M2_454
timestamp 1745462530
transform 1 0 2204 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_455
timestamp 1745462530
transform 1 0 2204 0 1 2125
box -3 -3 3 3
use M3_M2  M3_M2_456
timestamp 1745462530
transform 1 0 2196 0 1 2665
box -3 -3 3 3
use M3_M2  M3_M2_457
timestamp 1745462530
transform 1 0 2188 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_458
timestamp 1745462530
transform 1 0 2180 0 1 2125
box -3 -3 3 3
use M3_M2  M3_M2_459
timestamp 1745462530
transform 1 0 2148 0 1 2665
box -3 -3 3 3
use M3_M2  M3_M2_460
timestamp 1745462530
transform 1 0 2140 0 1 2125
box -3 -3 3 3
use M3_M2  M3_M2_461
timestamp 1745462530
transform 1 0 2460 0 1 1775
box -3 -3 3 3
use M3_M2  M3_M2_462
timestamp 1745462530
transform 1 0 2388 0 1 1775
box -3 -3 3 3
use M3_M2  M3_M2_463
timestamp 1745462530
transform 1 0 2372 0 1 1775
box -3 -3 3 3
use M3_M2  M3_M2_464
timestamp 1745462530
transform 1 0 2324 0 1 1775
box -3 -3 3 3
use M3_M2  M3_M2_465
timestamp 1745462530
transform 1 0 1004 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_466
timestamp 1745462530
transform 1 0 932 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_467
timestamp 1745462530
transform 1 0 908 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_468
timestamp 1745462530
transform 1 0 852 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_469
timestamp 1745462530
transform 1 0 812 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_470
timestamp 1745462530
transform 1 0 2244 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_471
timestamp 1745462530
transform 1 0 2236 0 1 2295
box -3 -3 3 3
use M3_M2  M3_M2_472
timestamp 1745462530
transform 1 0 2196 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_473
timestamp 1745462530
transform 1 0 2164 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_474
timestamp 1745462530
transform 1 0 2164 0 1 2295
box -3 -3 3 3
use M3_M2  M3_M2_475
timestamp 1745462530
transform 1 0 2092 0 1 2475
box -3 -3 3 3
use M3_M2  M3_M2_476
timestamp 1745462530
transform 1 0 2092 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_477
timestamp 1745462530
transform 1 0 2052 0 1 2475
box -3 -3 3 3
use M3_M2  M3_M2_478
timestamp 1745462530
transform 1 0 3252 0 1 575
box -3 -3 3 3
use M3_M2  M3_M2_479
timestamp 1745462530
transform 1 0 3220 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_480
timestamp 1745462530
transform 1 0 3196 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_481
timestamp 1745462530
transform 1 0 1044 0 1 2475
box -3 -3 3 3
use M3_M2  M3_M2_482
timestamp 1745462530
transform 1 0 996 0 1 2475
box -3 -3 3 3
use M3_M2  M3_M2_483
timestamp 1745462530
transform 1 0 916 0 1 2475
box -3 -3 3 3
use M3_M2  M3_M2_484
timestamp 1745462530
transform 1 0 908 0 1 2405
box -3 -3 3 3
use M3_M2  M3_M2_485
timestamp 1745462530
transform 1 0 852 0 1 2405
box -3 -3 3 3
use M3_M2  M3_M2_486
timestamp 1745462530
transform 1 0 2636 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_487
timestamp 1745462530
transform 1 0 2596 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_488
timestamp 1745462530
transform 1 0 2148 0 1 2295
box -3 -3 3 3
use M3_M2  M3_M2_489
timestamp 1745462530
transform 1 0 2108 0 1 2295
box -3 -3 3 3
use M3_M2  M3_M2_490
timestamp 1745462530
transform 1 0 1340 0 1 2295
box -3 -3 3 3
use M3_M2  M3_M2_491
timestamp 1745462530
transform 1 0 2204 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_492
timestamp 1745462530
transform 1 0 2148 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_493
timestamp 1745462530
transform 1 0 1796 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_494
timestamp 1745462530
transform 1 0 1772 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_495
timestamp 1745462530
transform 1 0 1556 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_496
timestamp 1745462530
transform 1 0 1420 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_497
timestamp 1745462530
transform 1 0 1380 0 1 2055
box -3 -3 3 3
use M3_M2  M3_M2_498
timestamp 1745462530
transform 1 0 1380 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_499
timestamp 1745462530
transform 1 0 1212 0 1 2065
box -3 -3 3 3
use M3_M2  M3_M2_500
timestamp 1745462530
transform 1 0 1180 0 1 2065
box -3 -3 3 3
use M3_M2  M3_M2_501
timestamp 1745462530
transform 1 0 1748 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_502
timestamp 1745462530
transform 1 0 1692 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_503
timestamp 1745462530
transform 1 0 1492 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_504
timestamp 1745462530
transform 1 0 1436 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_505
timestamp 1745462530
transform 1 0 1412 0 1 2555
box -3 -3 3 3
use M3_M2  M3_M2_506
timestamp 1745462530
transform 1 0 1292 0 1 2555
box -3 -3 3 3
use M3_M2  M3_M2_507
timestamp 1745462530
transform 1 0 1228 0 1 2555
box -3 -3 3 3
use M3_M2  M3_M2_508
timestamp 1745462530
transform 1 0 1180 0 1 2555
box -3 -3 3 3
use M3_M2  M3_M2_509
timestamp 1745462530
transform 1 0 1716 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_510
timestamp 1745462530
transform 1 0 1540 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_511
timestamp 1745462530
transform 1 0 1492 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_512
timestamp 1745462530
transform 1 0 1340 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_513
timestamp 1745462530
transform 1 0 1220 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_514
timestamp 1745462530
transform 1 0 1156 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_515
timestamp 1745462530
transform 1 0 804 0 1 2935
box -3 -3 3 3
use M3_M2  M3_M2_516
timestamp 1745462530
transform 1 0 756 0 1 2935
box -3 -3 3 3
use M3_M2  M3_M2_517
timestamp 1745462530
transform 1 0 420 0 1 2935
box -3 -3 3 3
use M3_M2  M3_M2_518
timestamp 1745462530
transform 1 0 420 0 1 2765
box -3 -3 3 3
use M3_M2  M3_M2_519
timestamp 1745462530
transform 1 0 380 0 1 2765
box -3 -3 3 3
use M3_M2  M3_M2_520
timestamp 1745462530
transform 1 0 324 0 1 2765
box -3 -3 3 3
use M3_M2  M3_M2_521
timestamp 1745462530
transform 1 0 260 0 1 2765
box -3 -3 3 3
use M3_M2  M3_M2_522
timestamp 1745462530
transform 1 0 764 0 1 2675
box -3 -3 3 3
use M3_M2  M3_M2_523
timestamp 1745462530
transform 1 0 652 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_524
timestamp 1745462530
transform 1 0 564 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_525
timestamp 1745462530
transform 1 0 564 0 1 2765
box -3 -3 3 3
use M3_M2  M3_M2_526
timestamp 1745462530
transform 1 0 564 0 1 2675
box -3 -3 3 3
use M3_M2  M3_M2_527
timestamp 1745462530
transform 1 0 564 0 1 2565
box -3 -3 3 3
use M3_M2  M3_M2_528
timestamp 1745462530
transform 1 0 516 0 1 2765
box -3 -3 3 3
use M3_M2  M3_M2_529
timestamp 1745462530
transform 1 0 508 0 1 2565
box -3 -3 3 3
use M3_M2  M3_M2_530
timestamp 1745462530
transform 1 0 428 0 1 2785
box -3 -3 3 3
use M3_M2  M3_M2_531
timestamp 1745462530
transform 1 0 324 0 1 2605
box -3 -3 3 3
use M3_M2  M3_M2_532
timestamp 1745462530
transform 1 0 252 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_533
timestamp 1745462530
transform 1 0 212 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_534
timestamp 1745462530
transform 1 0 196 0 1 2605
box -3 -3 3 3
use M3_M2  M3_M2_535
timestamp 1745462530
transform 1 0 940 0 1 2885
box -3 -3 3 3
use M3_M2  M3_M2_536
timestamp 1745462530
transform 1 0 900 0 1 2885
box -3 -3 3 3
use M3_M2  M3_M2_537
timestamp 1745462530
transform 1 0 380 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_538
timestamp 1745462530
transform 1 0 332 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_539
timestamp 1745462530
transform 1 0 244 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_540
timestamp 1745462530
transform 1 0 196 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_541
timestamp 1745462530
transform 1 0 364 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_542
timestamp 1745462530
transform 1 0 204 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_543
timestamp 1745462530
transform 1 0 180 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_544
timestamp 1745462530
transform 1 0 372 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_545
timestamp 1745462530
transform 1 0 284 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_546
timestamp 1745462530
transform 1 0 244 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_547
timestamp 1745462530
transform 1 0 212 0 1 535
box -3 -3 3 3
use M3_M2  M3_M2_548
timestamp 1745462530
transform 1 0 196 0 1 535
box -3 -3 3 3
use M3_M2  M3_M2_549
timestamp 1745462530
transform 1 0 196 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_550
timestamp 1745462530
transform 1 0 460 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_551
timestamp 1745462530
transform 1 0 380 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_552
timestamp 1745462530
transform 1 0 292 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_553
timestamp 1745462530
transform 1 0 244 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_554
timestamp 1745462530
transform 1 0 188 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_555
timestamp 1745462530
transform 1 0 684 0 1 165
box -3 -3 3 3
use M3_M2  M3_M2_556
timestamp 1745462530
transform 1 0 660 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_557
timestamp 1745462530
transform 1 0 628 0 1 165
box -3 -3 3 3
use M3_M2  M3_M2_558
timestamp 1745462530
transform 1 0 620 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_559
timestamp 1745462530
transform 1 0 532 0 1 165
box -3 -3 3 3
use M3_M2  M3_M2_560
timestamp 1745462530
transform 1 0 1884 0 1 415
box -3 -3 3 3
use M3_M2  M3_M2_561
timestamp 1745462530
transform 1 0 1804 0 1 415
box -3 -3 3 3
use M3_M2  M3_M2_562
timestamp 1745462530
transform 1 0 1668 0 1 415
box -3 -3 3 3
use M3_M2  M3_M2_563
timestamp 1745462530
transform 1 0 1468 0 1 405
box -3 -3 3 3
use M3_M2  M3_M2_564
timestamp 1745462530
transform 1 0 1388 0 1 485
box -3 -3 3 3
use M3_M2  M3_M2_565
timestamp 1745462530
transform 1 0 1388 0 1 405
box -3 -3 3 3
use M3_M2  M3_M2_566
timestamp 1745462530
transform 1 0 1124 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_567
timestamp 1745462530
transform 1 0 1124 0 1 485
box -3 -3 3 3
use M3_M2  M3_M2_568
timestamp 1745462530
transform 1 0 1020 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_569
timestamp 1745462530
transform 1 0 1876 0 1 215
box -3 -3 3 3
use M3_M2  M3_M2_570
timestamp 1745462530
transform 1 0 1764 0 1 215
box -3 -3 3 3
use M3_M2  M3_M2_571
timestamp 1745462530
transform 1 0 1660 0 1 215
box -3 -3 3 3
use M3_M2  M3_M2_572
timestamp 1745462530
transform 1 0 1540 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_573
timestamp 1745462530
transform 1 0 1436 0 1 215
box -3 -3 3 3
use M3_M2  M3_M2_574
timestamp 1745462530
transform 1 0 1340 0 1 215
box -3 -3 3 3
use M3_M2  M3_M2_575
timestamp 1745462530
transform 1 0 1868 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_576
timestamp 1745462530
transform 1 0 1812 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_577
timestamp 1745462530
transform 1 0 1708 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_578
timestamp 1745462530
transform 1 0 1604 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_579
timestamp 1745462530
transform 1 0 1380 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_580
timestamp 1745462530
transform 1 0 1324 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_581
timestamp 1745462530
transform 1 0 1244 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_582
timestamp 1745462530
transform 1 0 1876 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_583
timestamp 1745462530
transform 1 0 1692 0 1 295
box -3 -3 3 3
use M3_M2  M3_M2_584
timestamp 1745462530
transform 1 0 1532 0 1 295
box -3 -3 3 3
use M3_M2  M3_M2_585
timestamp 1745462530
transform 1 0 1468 0 1 115
box -3 -3 3 3
use M3_M2  M3_M2_586
timestamp 1745462530
transform 1 0 1404 0 1 295
box -3 -3 3 3
use M3_M2  M3_M2_587
timestamp 1745462530
transform 1 0 1404 0 1 115
box -3 -3 3 3
use M3_M2  M3_M2_588
timestamp 1745462530
transform 1 0 1300 0 1 115
box -3 -3 3 3
use M3_M2  M3_M2_589
timestamp 1745462530
transform 1 0 3068 0 1 685
box -3 -3 3 3
use M3_M2  M3_M2_590
timestamp 1745462530
transform 1 0 3020 0 1 685
box -3 -3 3 3
use M3_M2  M3_M2_591
timestamp 1745462530
transform 1 0 2980 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_592
timestamp 1745462530
transform 1 0 2980 0 1 685
box -3 -3 3 3
use M3_M2  M3_M2_593
timestamp 1745462530
transform 1 0 2716 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_594
timestamp 1745462530
transform 1 0 2268 0 1 725
box -3 -3 3 3
use M3_M2  M3_M2_595
timestamp 1745462530
transform 1 0 2188 0 1 725
box -3 -3 3 3
use M3_M2  M3_M2_596
timestamp 1745462530
transform 1 0 2772 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_597
timestamp 1745462530
transform 1 0 2676 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_598
timestamp 1745462530
transform 1 0 2580 0 1 215
box -3 -3 3 3
use M3_M2  M3_M2_599
timestamp 1745462530
transform 1 0 2508 0 1 215
box -3 -3 3 3
use M3_M2  M3_M2_600
timestamp 1745462530
transform 1 0 2284 0 1 215
box -3 -3 3 3
use M3_M2  M3_M2_601
timestamp 1745462530
transform 1 0 2220 0 1 215
box -3 -3 3 3
use M3_M2  M3_M2_602
timestamp 1745462530
transform 1 0 2972 0 1 445
box -3 -3 3 3
use M3_M2  M3_M2_603
timestamp 1745462530
transform 1 0 2900 0 1 445
box -3 -3 3 3
use M3_M2  M3_M2_604
timestamp 1745462530
transform 1 0 2764 0 1 475
box -3 -3 3 3
use M3_M2  M3_M2_605
timestamp 1745462530
transform 1 0 2700 0 1 475
box -3 -3 3 3
use M3_M2  M3_M2_606
timestamp 1745462530
transform 1 0 2700 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_607
timestamp 1745462530
transform 1 0 2268 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_608
timestamp 1745462530
transform 1 0 2268 0 1 415
box -3 -3 3 3
use M3_M2  M3_M2_609
timestamp 1745462530
transform 1 0 2228 0 1 415
box -3 -3 3 3
use M3_M2  M3_M2_610
timestamp 1745462530
transform 1 0 3068 0 1 215
box -3 -3 3 3
use M3_M2  M3_M2_611
timestamp 1745462530
transform 1 0 2996 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_612
timestamp 1745462530
transform 1 0 2996 0 1 215
box -3 -3 3 3
use M3_M2  M3_M2_613
timestamp 1745462530
transform 1 0 2940 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_614
timestamp 1745462530
transform 1 0 2940 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_615
timestamp 1745462530
transform 1 0 2644 0 1 365
box -3 -3 3 3
use M3_M2  M3_M2_616
timestamp 1745462530
transform 1 0 2596 0 1 365
box -3 -3 3 3
use M3_M2  M3_M2_617
timestamp 1745462530
transform 1 0 2492 0 1 365
box -3 -3 3 3
use M3_M2  M3_M2_618
timestamp 1745462530
transform 1 0 2436 0 1 365
box -3 -3 3 3
use M3_M2  M3_M2_619
timestamp 1745462530
transform 1 0 3844 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_620
timestamp 1745462530
transform 1 0 3796 0 1 415
box -3 -3 3 3
use M3_M2  M3_M2_621
timestamp 1745462530
transform 1 0 3796 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_622
timestamp 1745462530
transform 1 0 3708 0 1 415
box -3 -3 3 3
use M3_M2  M3_M2_623
timestamp 1745462530
transform 1 0 3500 0 1 415
box -3 -3 3 3
use M3_M2  M3_M2_624
timestamp 1745462530
transform 1 0 3348 0 1 415
box -3 -3 3 3
use M3_M2  M3_M2_625
timestamp 1745462530
transform 1 0 4220 0 1 205
box -3 -3 3 3
use M3_M2  M3_M2_626
timestamp 1745462530
transform 1 0 4116 0 1 205
box -3 -3 3 3
use M3_M2  M3_M2_627
timestamp 1745462530
transform 1 0 4068 0 1 205
box -3 -3 3 3
use M3_M2  M3_M2_628
timestamp 1745462530
transform 1 0 4044 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_629
timestamp 1745462530
transform 1 0 3988 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_630
timestamp 1745462530
transform 1 0 3988 0 1 205
box -3 -3 3 3
use M3_M2  M3_M2_631
timestamp 1745462530
transform 1 0 3748 0 1 205
box -3 -3 3 3
use M3_M2  M3_M2_632
timestamp 1745462530
transform 1 0 3948 0 1 325
box -3 -3 3 3
use M3_M2  M3_M2_633
timestamp 1745462530
transform 1 0 3748 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_634
timestamp 1745462530
transform 1 0 3724 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_635
timestamp 1745462530
transform 1 0 3716 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_636
timestamp 1745462530
transform 1 0 3636 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_637
timestamp 1745462530
transform 1 0 3484 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_638
timestamp 1745462530
transform 1 0 3364 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_639
timestamp 1745462530
transform 1 0 4308 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_640
timestamp 1745462530
transform 1 0 4252 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_641
timestamp 1745462530
transform 1 0 4204 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_642
timestamp 1745462530
transform 1 0 4148 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_643
timestamp 1745462530
transform 1 0 4124 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_644
timestamp 1745462530
transform 1 0 3804 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_645
timestamp 1745462530
transform 1 0 3796 0 1 1435
box -3 -3 3 3
use M3_M2  M3_M2_646
timestamp 1745462530
transform 1 0 3676 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_647
timestamp 1745462530
transform 1 0 3660 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_648
timestamp 1745462530
transform 1 0 3660 0 1 1435
box -3 -3 3 3
use M3_M2  M3_M2_649
timestamp 1745462530
transform 1 0 3500 0 1 1435
box -3 -3 3 3
use M3_M2  M3_M2_650
timestamp 1745462530
transform 1 0 3468 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_651
timestamp 1745462530
transform 1 0 4204 0 1 1475
box -3 -3 3 3
use M3_M2  M3_M2_652
timestamp 1745462530
transform 1 0 4044 0 1 1475
box -3 -3 3 3
use M3_M2  M3_M2_653
timestamp 1745462530
transform 1 0 3852 0 1 1895
box -3 -3 3 3
use M3_M2  M3_M2_654
timestamp 1745462530
transform 1 0 3844 0 1 1645
box -3 -3 3 3
use M3_M2  M3_M2_655
timestamp 1745462530
transform 1 0 3836 0 1 2045
box -3 -3 3 3
use M3_M2  M3_M2_656
timestamp 1745462530
transform 1 0 3836 0 1 1895
box -3 -3 3 3
use M3_M2  M3_M2_657
timestamp 1745462530
transform 1 0 3804 0 1 1645
box -3 -3 3 3
use M3_M2  M3_M2_658
timestamp 1745462530
transform 1 0 3796 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_659
timestamp 1745462530
transform 1 0 3772 0 1 2045
box -3 -3 3 3
use M3_M2  M3_M2_660
timestamp 1745462530
transform 1 0 3676 0 1 2045
box -3 -3 3 3
use M3_M2  M3_M2_661
timestamp 1745462530
transform 1 0 3636 0 1 1615
box -3 -3 3 3
use M3_M2  M3_M2_662
timestamp 1745462530
transform 1 0 3636 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_663
timestamp 1745462530
transform 1 0 3564 0 1 1615
box -3 -3 3 3
use M3_M2  M3_M2_664
timestamp 1745462530
transform 1 0 4300 0 1 1575
box -3 -3 3 3
use M3_M2  M3_M2_665
timestamp 1745462530
transform 1 0 4276 0 1 1845
box -3 -3 3 3
use M3_M2  M3_M2_666
timestamp 1745462530
transform 1 0 4276 0 1 1575
box -3 -3 3 3
use M3_M2  M3_M2_667
timestamp 1745462530
transform 1 0 4268 0 1 2005
box -3 -3 3 3
use M3_M2  M3_M2_668
timestamp 1745462530
transform 1 0 4204 0 1 2005
box -3 -3 3 3
use M3_M2  M3_M2_669
timestamp 1745462530
transform 1 0 4180 0 1 1845
box -3 -3 3 3
use M3_M2  M3_M2_670
timestamp 1745462530
transform 1 0 4156 0 1 1575
box -3 -3 3 3
use M3_M2  M3_M2_671
timestamp 1745462530
transform 1 0 4140 0 1 2005
box -3 -3 3 3
use M3_M2  M3_M2_672
timestamp 1745462530
transform 1 0 3980 0 1 1575
box -3 -3 3 3
use M3_M2  M3_M2_673
timestamp 1745462530
transform 1 0 4220 0 1 2375
box -3 -3 3 3
use M3_M2  M3_M2_674
timestamp 1745462530
transform 1 0 4140 0 1 2375
box -3 -3 3 3
use M3_M2  M3_M2_675
timestamp 1745462530
transform 1 0 3924 0 1 2375
box -3 -3 3 3
use M3_M2  M3_M2_676
timestamp 1745462530
transform 1 0 3604 0 1 2375
box -3 -3 3 3
use M3_M2  M3_M2_677
timestamp 1745462530
transform 1 0 3356 0 1 2375
box -3 -3 3 3
use M3_M2  M3_M2_678
timestamp 1745462530
transform 1 0 3356 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_679
timestamp 1745462530
transform 1 0 3236 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_680
timestamp 1745462530
transform 1 0 4084 0 1 2985
box -3 -3 3 3
use M3_M2  M3_M2_681
timestamp 1745462530
transform 1 0 4060 0 1 2985
box -3 -3 3 3
use M3_M2  M3_M2_682
timestamp 1745462530
transform 1 0 3836 0 1 2985
box -3 -3 3 3
use M3_M2  M3_M2_683
timestamp 1745462530
transform 1 0 3836 0 1 2895
box -3 -3 3 3
use M3_M2  M3_M2_684
timestamp 1745462530
transform 1 0 3692 0 1 2895
box -3 -3 3 3
use M3_M2  M3_M2_685
timestamp 1745462530
transform 1 0 3460 0 1 2905
box -3 -3 3 3
use M3_M2  M3_M2_686
timestamp 1745462530
transform 1 0 3164 0 1 2905
box -3 -3 3 3
use M3_M2  M3_M2_687
timestamp 1745462530
transform 1 0 1900 0 1 2845
box -3 -3 3 3
use M3_M2  M3_M2_688
timestamp 1745462530
transform 1 0 1828 0 1 2845
box -3 -3 3 3
use M3_M2  M3_M2_689
timestamp 1745462530
transform 1 0 1828 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_690
timestamp 1745462530
transform 1 0 1764 0 1 2845
box -3 -3 3 3
use M3_M2  M3_M2_691
timestamp 1745462530
transform 1 0 1764 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_692
timestamp 1745462530
transform 1 0 1612 0 1 2845
box -3 -3 3 3
use M3_M2  M3_M2_693
timestamp 1745462530
transform 1 0 1316 0 1 2835
box -3 -3 3 3
use M3_M2  M3_M2_694
timestamp 1745462530
transform 1 0 1276 0 1 2835
box -3 -3 3 3
use M3_M2  M3_M2_695
timestamp 1745462530
transform 1 0 1996 0 1 2205
box -3 -3 3 3
use M3_M2  M3_M2_696
timestamp 1745462530
transform 1 0 1916 0 1 2205
box -3 -3 3 3
use M3_M2  M3_M2_697
timestamp 1745462530
transform 1 0 1716 0 1 2205
box -3 -3 3 3
use M3_M2  M3_M2_698
timestamp 1745462530
transform 1 0 1652 0 1 2205
box -3 -3 3 3
use M3_M2  M3_M2_699
timestamp 1745462530
transform 1 0 1572 0 1 2205
box -3 -3 3 3
use M3_M2  M3_M2_700
timestamp 1745462530
transform 1 0 1308 0 1 2205
box -3 -3 3 3
use M3_M2  M3_M2_701
timestamp 1745462530
transform 1 0 1244 0 1 2205
box -3 -3 3 3
use M3_M2  M3_M2_702
timestamp 1745462530
transform 1 0 1916 0 1 2625
box -3 -3 3 3
use M3_M2  M3_M2_703
timestamp 1745462530
transform 1 0 1844 0 1 2625
box -3 -3 3 3
use M3_M2  M3_M2_704
timestamp 1745462530
transform 1 0 1716 0 1 2675
box -3 -3 3 3
use M3_M2  M3_M2_705
timestamp 1745462530
transform 1 0 1716 0 1 2625
box -3 -3 3 3
use M3_M2  M3_M2_706
timestamp 1745462530
transform 1 0 1692 0 1 2675
box -3 -3 3 3
use M3_M2  M3_M2_707
timestamp 1745462530
transform 1 0 1564 0 1 2675
box -3 -3 3 3
use M3_M2  M3_M2_708
timestamp 1745462530
transform 1 0 1284 0 1 2725
box -3 -3 3 3
use M3_M2  M3_M2_709
timestamp 1745462530
transform 1 0 1284 0 1 2675
box -3 -3 3 3
use M3_M2  M3_M2_710
timestamp 1745462530
transform 1 0 1236 0 1 2725
box -3 -3 3 3
use M3_M2  M3_M2_711
timestamp 1745462530
transform 1 0 484 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_712
timestamp 1745462530
transform 1 0 436 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_713
timestamp 1745462530
transform 1 0 380 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_714
timestamp 1745462530
transform 1 0 300 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_715
timestamp 1745462530
transform 1 0 244 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_716
timestamp 1745462530
transform 1 0 436 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_717
timestamp 1745462530
transform 1 0 356 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_718
timestamp 1745462530
transform 1 0 292 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_719
timestamp 1745462530
transform 1 0 228 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_720
timestamp 1745462530
transform 1 0 740 0 1 1665
box -3 -3 3 3
use M3_M2  M3_M2_721
timestamp 1745462530
transform 1 0 700 0 1 1665
box -3 -3 3 3
use M3_M2  M3_M2_722
timestamp 1745462530
transform 1 0 676 0 1 1665
box -3 -3 3 3
use M3_M2  M3_M2_723
timestamp 1745462530
transform 1 0 628 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_724
timestamp 1745462530
transform 1 0 628 0 1 1665
box -3 -3 3 3
use M3_M2  M3_M2_725
timestamp 1745462530
transform 1 0 588 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_726
timestamp 1745462530
transform 1 0 532 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_727
timestamp 1745462530
transform 1 0 500 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_728
timestamp 1745462530
transform 1 0 436 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_729
timestamp 1745462530
transform 1 0 372 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_730
timestamp 1745462530
transform 1 0 308 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_731
timestamp 1745462530
transform 1 0 244 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_732
timestamp 1745462530
transform 1 0 500 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_733
timestamp 1745462530
transform 1 0 428 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_734
timestamp 1745462530
transform 1 0 396 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_735
timestamp 1745462530
transform 1 0 332 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_736
timestamp 1745462530
transform 1 0 228 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_737
timestamp 1745462530
transform 1 0 964 0 1 1335
box -3 -3 3 3
use M3_M2  M3_M2_738
timestamp 1745462530
transform 1 0 876 0 1 1335
box -3 -3 3 3
use M3_M2  M3_M2_739
timestamp 1745462530
transform 1 0 860 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_740
timestamp 1745462530
transform 1 0 812 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_741
timestamp 1745462530
transform 1 0 780 0 1 1465
box -3 -3 3 3
use M3_M2  M3_M2_742
timestamp 1745462530
transform 1 0 780 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_743
timestamp 1745462530
transform 1 0 780 0 1 1335
box -3 -3 3 3
use M3_M2  M3_M2_744
timestamp 1745462530
transform 1 0 724 0 1 1465
box -3 -3 3 3
use M3_M2  M3_M2_745
timestamp 1745462530
transform 1 0 700 0 1 1335
box -3 -3 3 3
use M3_M2  M3_M2_746
timestamp 1745462530
transform 1 0 1708 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_747
timestamp 1745462530
transform 1 0 1644 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_748
timestamp 1745462530
transform 1 0 1508 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_749
timestamp 1745462530
transform 1 0 1484 0 1 235
box -3 -3 3 3
use M3_M2  M3_M2_750
timestamp 1745462530
transform 1 0 1180 0 1 235
box -3 -3 3 3
use M3_M2  M3_M2_751
timestamp 1745462530
transform 1 0 2020 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_752
timestamp 1745462530
transform 1 0 1964 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_753
timestamp 1745462530
transform 1 0 1964 0 1 875
box -3 -3 3 3
use M3_M2  M3_M2_754
timestamp 1745462530
transform 1 0 1812 0 1 875
box -3 -3 3 3
use M3_M2  M3_M2_755
timestamp 1745462530
transform 1 0 1804 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_756
timestamp 1745462530
transform 1 0 1612 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_757
timestamp 1745462530
transform 1 0 1436 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_758
timestamp 1745462530
transform 1 0 2044 0 1 1275
box -3 -3 3 3
use M3_M2  M3_M2_759
timestamp 1745462530
transform 1 0 2012 0 1 1275
box -3 -3 3 3
use M3_M2  M3_M2_760
timestamp 1745462530
transform 1 0 1852 0 1 1285
box -3 -3 3 3
use M3_M2  M3_M2_761
timestamp 1745462530
transform 1 0 1636 0 1 1285
box -3 -3 3 3
use M3_M2  M3_M2_762
timestamp 1745462530
transform 1 0 1604 0 1 1285
box -3 -3 3 3
use M3_M2  M3_M2_763
timestamp 1745462530
transform 1 0 1484 0 1 1285
box -3 -3 3 3
use M3_M2  M3_M2_764
timestamp 1745462530
transform 1 0 1436 0 1 1285
box -3 -3 3 3
use M3_M2  M3_M2_765
timestamp 1745462530
transform 1 0 2044 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_766
timestamp 1745462530
transform 1 0 2044 0 1 1335
box -3 -3 3 3
use M3_M2  M3_M2_767
timestamp 1745462530
transform 1 0 2012 0 1 1335
box -3 -3 3 3
use M3_M2  M3_M2_768
timestamp 1745462530
transform 1 0 1948 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_769
timestamp 1745462530
transform 1 0 1852 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_770
timestamp 1745462530
transform 1 0 1676 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_771
timestamp 1745462530
transform 1 0 1612 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_772
timestamp 1745462530
transform 1 0 1540 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_773
timestamp 1745462530
transform 1 0 2916 0 1 205
box -3 -3 3 3
use M3_M2  M3_M2_774
timestamp 1745462530
transform 1 0 2860 0 1 405
box -3 -3 3 3
use M3_M2  M3_M2_775
timestamp 1745462530
transform 1 0 2804 0 1 405
box -3 -3 3 3
use M3_M2  M3_M2_776
timestamp 1745462530
transform 1 0 2804 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_777
timestamp 1745462530
transform 1 0 2756 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_778
timestamp 1745462530
transform 1 0 2548 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_779
timestamp 1745462530
transform 1 0 2548 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_780
timestamp 1745462530
transform 1 0 2380 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_781
timestamp 1745462530
transform 1 0 2316 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_782
timestamp 1745462530
transform 1 0 2252 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_783
timestamp 1745462530
transform 1 0 2900 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_784
timestamp 1745462530
transform 1 0 2740 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_785
timestamp 1745462530
transform 1 0 2572 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_786
timestamp 1745462530
transform 1 0 2364 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_787
timestamp 1745462530
transform 1 0 2364 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_788
timestamp 1745462530
transform 1 0 2300 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_789
timestamp 1745462530
transform 1 0 2852 0 1 1065
box -3 -3 3 3
use M3_M2  M3_M2_790
timestamp 1745462530
transform 1 0 2692 0 1 1065
box -3 -3 3 3
use M3_M2  M3_M2_791
timestamp 1745462530
transform 1 0 2684 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_792
timestamp 1745462530
transform 1 0 2636 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_793
timestamp 1745462530
transform 1 0 2372 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_794
timestamp 1745462530
transform 1 0 2324 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_795
timestamp 1745462530
transform 1 0 2860 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_796
timestamp 1745462530
transform 1 0 2820 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_797
timestamp 1745462530
transform 1 0 2820 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_798
timestamp 1745462530
transform 1 0 2788 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_799
timestamp 1745462530
transform 1 0 2788 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_800
timestamp 1745462530
transform 1 0 2676 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_801
timestamp 1745462530
transform 1 0 2652 0 1 1435
box -3 -3 3 3
use M3_M2  M3_M2_802
timestamp 1745462530
transform 1 0 2628 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_803
timestamp 1745462530
transform 1 0 2620 0 1 1435
box -3 -3 3 3
use M3_M2  M3_M2_804
timestamp 1745462530
transform 1 0 2412 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_805
timestamp 1745462530
transform 1 0 3452 0 1 295
box -3 -3 3 3
use M3_M2  M3_M2_806
timestamp 1745462530
transform 1 0 3396 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_807
timestamp 1745462530
transform 1 0 3340 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_808
timestamp 1745462530
transform 1 0 3324 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_809
timestamp 1745462530
transform 1 0 3284 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_810
timestamp 1745462530
transform 1 0 3228 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_811
timestamp 1745462530
transform 1 0 4324 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_812
timestamp 1745462530
transform 1 0 4260 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_813
timestamp 1745462530
transform 1 0 4244 0 1 845
box -3 -3 3 3
use M3_M2  M3_M2_814
timestamp 1745462530
transform 1 0 4204 0 1 845
box -3 -3 3 3
use M3_M2  M3_M2_815
timestamp 1745462530
transform 1 0 4164 0 1 845
box -3 -3 3 3
use M3_M2  M3_M2_816
timestamp 1745462530
transform 1 0 4068 0 1 845
box -3 -3 3 3
use M3_M2  M3_M2_817
timestamp 1745462530
transform 1 0 3972 0 1 845
box -3 -3 3 3
use M3_M2  M3_M2_818
timestamp 1745462530
transform 1 0 4236 0 1 1055
box -3 -3 3 3
use M3_M2  M3_M2_819
timestamp 1745462530
transform 1 0 4164 0 1 1065
box -3 -3 3 3
use M3_M2  M3_M2_820
timestamp 1745462530
transform 1 0 4084 0 1 1065
box -3 -3 3 3
use M3_M2  M3_M2_821
timestamp 1745462530
transform 1 0 3820 0 1 1065
box -3 -3 3 3
use M3_M2  M3_M2_822
timestamp 1745462530
transform 1 0 3468 0 1 1065
box -3 -3 3 3
use M3_M2  M3_M2_823
timestamp 1745462530
transform 1 0 3404 0 1 1065
box -3 -3 3 3
use M3_M2  M3_M2_824
timestamp 1745462530
transform 1 0 3940 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_825
timestamp 1745462530
transform 1 0 3892 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_826
timestamp 1745462530
transform 1 0 3796 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_827
timestamp 1745462530
transform 1 0 3628 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_828
timestamp 1745462530
transform 1 0 3476 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_829
timestamp 1745462530
transform 1 0 3388 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_830
timestamp 1745462530
transform 1 0 4236 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_831
timestamp 1745462530
transform 1 0 4228 0 1 1405
box -3 -3 3 3
use M3_M2  M3_M2_832
timestamp 1745462530
transform 1 0 4164 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_833
timestamp 1745462530
transform 1 0 4132 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_834
timestamp 1745462530
transform 1 0 4100 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_835
timestamp 1745462530
transform 1 0 3892 0 1 1775
box -3 -3 3 3
use M3_M2  M3_M2_836
timestamp 1745462530
transform 1 0 3868 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_837
timestamp 1745462530
transform 1 0 3732 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_838
timestamp 1745462530
transform 1 0 3620 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_839
timestamp 1745462530
transform 1 0 3620 0 1 2165
box -3 -3 3 3
use M3_M2  M3_M2_840
timestamp 1745462530
transform 1 0 3596 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_841
timestamp 1745462530
transform 1 0 3380 0 1 2165
box -3 -3 3 3
use M3_M2  M3_M2_842
timestamp 1745462530
transform 1 0 3292 0 1 1775
box -3 -3 3 3
use M3_M2  M3_M2_843
timestamp 1745462530
transform 1 0 3268 0 1 2165
box -3 -3 3 3
use M3_M2  M3_M2_844
timestamp 1745462530
transform 1 0 3132 0 1 2205
box -3 -3 3 3
use M3_M2  M3_M2_845
timestamp 1745462530
transform 1 0 2980 0 1 1875
box -3 -3 3 3
use M3_M2  M3_M2_846
timestamp 1745462530
transform 1 0 2884 0 1 1875
box -3 -3 3 3
use M3_M2  M3_M2_847
timestamp 1745462530
transform 1 0 2852 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_848
timestamp 1745462530
transform 1 0 2828 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_849
timestamp 1745462530
transform 1 0 2804 0 1 1875
box -3 -3 3 3
use M3_M2  M3_M2_850
timestamp 1745462530
transform 1 0 2948 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_851
timestamp 1745462530
transform 1 0 2788 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_852
timestamp 1745462530
transform 1 0 2716 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_853
timestamp 1745462530
transform 1 0 2700 0 1 2095
box -3 -3 3 3
use M3_M2  M3_M2_854
timestamp 1745462530
transform 1 0 2684 0 1 2095
box -3 -3 3 3
use M3_M2  M3_M2_855
timestamp 1745462530
transform 1 0 2684 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_856
timestamp 1745462530
transform 1 0 2652 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_857
timestamp 1745462530
transform 1 0 2652 0 1 2095
box -3 -3 3 3
use M3_M2  M3_M2_858
timestamp 1745462530
transform 1 0 4204 0 1 2695
box -3 -3 3 3
use M3_M2  M3_M2_859
timestamp 1745462530
transform 1 0 3884 0 1 2705
box -3 -3 3 3
use M3_M2  M3_M2_860
timestamp 1745462530
transform 1 0 3692 0 1 2705
box -3 -3 3 3
use M3_M2  M3_M2_861
timestamp 1745462530
transform 1 0 3460 0 1 2705
box -3 -3 3 3
use M3_M2  M3_M2_862
timestamp 1745462530
transform 1 0 3292 0 1 2705
box -3 -3 3 3
use M3_M2  M3_M2_863
timestamp 1745462530
transform 1 0 3916 0 1 2905
box -3 -3 3 3
use M3_M2  M3_M2_864
timestamp 1745462530
transform 1 0 3780 0 1 2915
box -3 -3 3 3
use M3_M2  M3_M2_865
timestamp 1745462530
transform 1 0 3708 0 1 2915
box -3 -3 3 3
use M3_M2  M3_M2_866
timestamp 1745462530
transform 1 0 3244 0 1 2915
box -3 -3 3 3
use M3_M2  M3_M2_867
timestamp 1745462530
transform 1 0 3020 0 1 2915
box -3 -3 3 3
use M3_M2  M3_M2_868
timestamp 1745462530
transform 1 0 4164 0 1 2855
box -3 -3 3 3
use M3_M2  M3_M2_869
timestamp 1745462530
transform 1 0 4100 0 1 2855
box -3 -3 3 3
use M3_M2  M3_M2_870
timestamp 1745462530
transform 1 0 3996 0 1 2855
box -3 -3 3 3
use M3_M2  M3_M2_871
timestamp 1745462530
transform 1 0 3876 0 1 2855
box -3 -3 3 3
use M3_M2  M3_M2_872
timestamp 1745462530
transform 1 0 3644 0 1 2855
box -3 -3 3 3
use M3_M2  M3_M2_873
timestamp 1745462530
transform 1 0 3412 0 1 2855
box -3 -3 3 3
use M3_M2  M3_M2_874
timestamp 1745462530
transform 1 0 3268 0 1 2855
box -3 -3 3 3
use M3_M2  M3_M2_875
timestamp 1745462530
transform 1 0 4244 0 1 2975
box -3 -3 3 3
use M3_M2  M3_M2_876
timestamp 1745462530
transform 1 0 4188 0 1 2975
box -3 -3 3 3
use M3_M2  M3_M2_877
timestamp 1745462530
transform 1 0 3748 0 1 2975
box -3 -3 3 3
use M3_M2  M3_M2_878
timestamp 1745462530
transform 1 0 3556 0 1 2985
box -3 -3 3 3
use M3_M2  M3_M2_879
timestamp 1745462530
transform 1 0 3316 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_880
timestamp 1745462530
transform 1 0 3220 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_881
timestamp 1745462530
transform 1 0 4228 0 1 2485
box -3 -3 3 3
use M3_M2  M3_M2_882
timestamp 1745462530
transform 1 0 3948 0 1 2485
box -3 -3 3 3
use M3_M2  M3_M2_883
timestamp 1745462530
transform 1 0 3852 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_884
timestamp 1745462530
transform 1 0 3852 0 1 2485
box -3 -3 3 3
use M3_M2  M3_M2_885
timestamp 1745462530
transform 1 0 3676 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_886
timestamp 1745462530
transform 1 0 3492 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_887
timestamp 1745462530
transform 1 0 3300 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_888
timestamp 1745462530
transform 1 0 3012 0 1 2565
box -3 -3 3 3
use M3_M2  M3_M2_889
timestamp 1745462530
transform 1 0 2892 0 1 2565
box -3 -3 3 3
use M3_M2  M3_M2_890
timestamp 1745462530
transform 1 0 2812 0 1 2565
box -3 -3 3 3
use M3_M2  M3_M2_891
timestamp 1745462530
transform 1 0 2812 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_892
timestamp 1745462530
transform 1 0 2788 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_893
timestamp 1745462530
transform 1 0 2708 0 1 2835
box -3 -3 3 3
use M3_M2  M3_M2_894
timestamp 1745462530
transform 1 0 2668 0 1 2835
box -3 -3 3 3
use M3_M2  M3_M2_895
timestamp 1745462530
transform 1 0 2628 0 1 2835
box -3 -3 3 3
use M3_M2  M3_M2_896
timestamp 1745462530
transform 1 0 2516 0 1 2835
box -3 -3 3 3
use M3_M2  M3_M2_897
timestamp 1745462530
transform 1 0 1308 0 1 3085
box -3 -3 3 3
use M3_M2  M3_M2_898
timestamp 1745462530
transform 1 0 1124 0 1 3495
box -3 -3 3 3
use M3_M2  M3_M2_899
timestamp 1745462530
transform 1 0 1084 0 1 3085
box -3 -3 3 3
use M3_M2  M3_M2_900
timestamp 1745462530
transform 1 0 1068 0 1 3495
box -3 -3 3 3
use M3_M2  M3_M2_901
timestamp 1745462530
transform 1 0 1068 0 1 3455
box -3 -3 3 3
use M3_M2  M3_M2_902
timestamp 1745462530
transform 1 0 1060 0 1 3615
box -3 -3 3 3
use M3_M2  M3_M2_903
timestamp 1745462530
transform 1 0 1060 0 1 3325
box -3 -3 3 3
use M3_M2  M3_M2_904
timestamp 1745462530
transform 1 0 1028 0 1 3325
box -3 -3 3 3
use M3_M2  M3_M2_905
timestamp 1745462530
transform 1 0 1004 0 1 3455
box -3 -3 3 3
use M3_M2  M3_M2_906
timestamp 1745462530
transform 1 0 988 0 1 3615
box -3 -3 3 3
use M3_M2  M3_M2_907
timestamp 1745462530
transform 1 0 980 0 1 3325
box -3 -3 3 3
use M3_M2  M3_M2_908
timestamp 1745462530
transform 1 0 1348 0 1 3265
box -3 -3 3 3
use M3_M2  M3_M2_909
timestamp 1745462530
transform 1 0 1300 0 1 3265
box -3 -3 3 3
use M3_M2  M3_M2_910
timestamp 1745462530
transform 1 0 1268 0 1 3265
box -3 -3 3 3
use M3_M2  M3_M2_911
timestamp 1745462530
transform 1 0 1100 0 1 3425
box -3 -3 3 3
use M3_M2  M3_M2_912
timestamp 1745462530
transform 1 0 844 0 1 3425
box -3 -3 3 3
use M3_M2  M3_M2_913
timestamp 1745462530
transform 1 0 948 0 1 3535
box -3 -3 3 3
use M3_M2  M3_M2_914
timestamp 1745462530
transform 1 0 860 0 1 3535
box -3 -3 3 3
use M3_M2  M3_M2_915
timestamp 1745462530
transform 1 0 988 0 1 3485
box -3 -3 3 3
use M3_M2  M3_M2_916
timestamp 1745462530
transform 1 0 820 0 1 3485
box -3 -3 3 3
use M3_M2  M3_M2_917
timestamp 1745462530
transform 1 0 1708 0 1 3245
box -3 -3 3 3
use M3_M2  M3_M2_918
timestamp 1745462530
transform 1 0 1516 0 1 3245
box -3 -3 3 3
use M3_M2  M3_M2_919
timestamp 1745462530
transform 1 0 1516 0 1 3185
box -3 -3 3 3
use M3_M2  M3_M2_920
timestamp 1745462530
transform 1 0 1436 0 1 3185
box -3 -3 3 3
use M3_M2  M3_M2_921
timestamp 1745462530
transform 1 0 1404 0 1 3305
box -3 -3 3 3
use M3_M2  M3_M2_922
timestamp 1745462530
transform 1 0 1372 0 1 3305
box -3 -3 3 3
use M3_M2  M3_M2_923
timestamp 1745462530
transform 1 0 1356 0 1 3185
box -3 -3 3 3
use M3_M2  M3_M2_924
timestamp 1745462530
transform 1 0 1356 0 1 3175
box -3 -3 3 3
use M3_M2  M3_M2_925
timestamp 1745462530
transform 1 0 1204 0 1 3175
box -3 -3 3 3
use M3_M2  M3_M2_926
timestamp 1745462530
transform 1 0 1588 0 1 3425
box -3 -3 3 3
use M3_M2  M3_M2_927
timestamp 1745462530
transform 1 0 1540 0 1 3425
box -3 -3 3 3
use M3_M2  M3_M2_928
timestamp 1745462530
transform 1 0 1740 0 1 3285
box -3 -3 3 3
use M3_M2  M3_M2_929
timestamp 1745462530
transform 1 0 1692 0 1 3285
box -3 -3 3 3
use M3_M2  M3_M2_930
timestamp 1745462530
transform 1 0 1684 0 1 3295
box -3 -3 3 3
use M3_M2  M3_M2_931
timestamp 1745462530
transform 1 0 1660 0 1 3295
box -3 -3 3 3
use M3_M2  M3_M2_932
timestamp 1745462530
transform 1 0 1628 0 1 3295
box -3 -3 3 3
use M3_M2  M3_M2_933
timestamp 1745462530
transform 1 0 1292 0 1 3295
box -3 -3 3 3
use M3_M2  M3_M2_934
timestamp 1745462530
transform 1 0 1268 0 1 3215
box -3 -3 3 3
use M3_M2  M3_M2_935
timestamp 1745462530
transform 1 0 1084 0 1 3215
box -3 -3 3 3
use M3_M2  M3_M2_936
timestamp 1745462530
transform 1 0 1732 0 1 3175
box -3 -3 3 3
use M3_M2  M3_M2_937
timestamp 1745462530
transform 1 0 1716 0 1 3175
box -3 -3 3 3
use M3_M2  M3_M2_938
timestamp 1745462530
transform 1 0 1668 0 1 3285
box -3 -3 3 3
use M3_M2  M3_M2_939
timestamp 1745462530
transform 1 0 1668 0 1 3175
box -3 -3 3 3
use M3_M2  M3_M2_940
timestamp 1745462530
transform 1 0 1620 0 1 3285
box -3 -3 3 3
use M3_M2  M3_M2_941
timestamp 1745462530
transform 1 0 1604 0 1 3175
box -3 -3 3 3
use M3_M2  M3_M2_942
timestamp 1745462530
transform 1 0 2588 0 1 3345
box -3 -3 3 3
use M3_M2  M3_M2_943
timestamp 1745462530
transform 1 0 2548 0 1 3345
box -3 -3 3 3
use M3_M2  M3_M2_944
timestamp 1745462530
transform 1 0 2532 0 1 3065
box -3 -3 3 3
use M3_M2  M3_M2_945
timestamp 1745462530
transform 1 0 2468 0 1 3205
box -3 -3 3 3
use M3_M2  M3_M2_946
timestamp 1745462530
transform 1 0 2468 0 1 3065
box -3 -3 3 3
use M3_M2  M3_M2_947
timestamp 1745462530
transform 1 0 2460 0 1 3485
box -3 -3 3 3
use M3_M2  M3_M2_948
timestamp 1745462530
transform 1 0 2428 0 1 3205
box -3 -3 3 3
use M3_M2  M3_M2_949
timestamp 1745462530
transform 1 0 2420 0 1 3485
box -3 -3 3 3
use M3_M2  M3_M2_950
timestamp 1745462530
transform 1 0 2156 0 1 3575
box -3 -3 3 3
use M3_M2  M3_M2_951
timestamp 1745462530
transform 1 0 2156 0 1 3485
box -3 -3 3 3
use M3_M2  M3_M2_952
timestamp 1745462530
transform 1 0 2124 0 1 3575
box -3 -3 3 3
use M3_M2  M3_M2_953
timestamp 1745462530
transform 1 0 3524 0 1 3555
box -3 -3 3 3
use M3_M2  M3_M2_954
timestamp 1745462530
transform 1 0 3492 0 1 3385
box -3 -3 3 3
use M3_M2  M3_M2_955
timestamp 1745462530
transform 1 0 3484 0 1 3555
box -3 -3 3 3
use M3_M2  M3_M2_956
timestamp 1745462530
transform 1 0 3452 0 1 3105
box -3 -3 3 3
use M3_M2  M3_M2_957
timestamp 1745462530
transform 1 0 3420 0 1 3385
box -3 -3 3 3
use M3_M2  M3_M2_958
timestamp 1745462530
transform 1 0 3380 0 1 3385
box -3 -3 3 3
use M3_M2  M3_M2_959
timestamp 1745462530
transform 1 0 3316 0 1 3105
box -3 -3 3 3
use M3_M2  M3_M2_960
timestamp 1745462530
transform 1 0 3308 0 1 3385
box -3 -3 3 3
use M3_M2  M3_M2_961
timestamp 1745462530
transform 1 0 3252 0 1 3385
box -3 -3 3 3
use M3_M2  M3_M2_962
timestamp 1745462530
transform 1 0 3140 0 1 3105
box -3 -3 3 3
use M3_M2  M3_M2_963
timestamp 1745462530
transform 1 0 1964 0 1 3085
box -3 -3 3 3
use M3_M2  M3_M2_964
timestamp 1745462530
transform 1 0 1908 0 1 3135
box -3 -3 3 3
use M3_M2  M3_M2_965
timestamp 1745462530
transform 1 0 1908 0 1 3085
box -3 -3 3 3
use M3_M2  M3_M2_966
timestamp 1745462530
transform 1 0 1884 0 1 2935
box -3 -3 3 3
use M3_M2  M3_M2_967
timestamp 1745462530
transform 1 0 1876 0 1 2775
box -3 -3 3 3
use M3_M2  M3_M2_968
timestamp 1745462530
transform 1 0 1828 0 1 2775
box -3 -3 3 3
use M3_M2  M3_M2_969
timestamp 1745462530
transform 1 0 1732 0 1 2935
box -3 -3 3 3
use M3_M2  M3_M2_970
timestamp 1745462530
transform 1 0 1724 0 1 3205
box -3 -3 3 3
use M3_M2  M3_M2_971
timestamp 1745462530
transform 1 0 1724 0 1 3145
box -3 -3 3 3
use M3_M2  M3_M2_972
timestamp 1745462530
transform 1 0 1548 0 1 3205
box -3 -3 3 3
use M3_M2  M3_M2_973
timestamp 1745462530
transform 1 0 1532 0 1 3205
box -3 -3 3 3
use M3_M2  M3_M2_974
timestamp 1745462530
transform 1 0 3620 0 1 3375
box -3 -3 3 3
use M3_M2  M3_M2_975
timestamp 1745462530
transform 1 0 3620 0 1 3055
box -3 -3 3 3
use M3_M2  M3_M2_976
timestamp 1745462530
transform 1 0 3580 0 1 3585
box -3 -3 3 3
use M3_M2  M3_M2_977
timestamp 1745462530
transform 1 0 3580 0 1 3475
box -3 -3 3 3
use M3_M2  M3_M2_978
timestamp 1745462530
transform 1 0 3580 0 1 3375
box -3 -3 3 3
use M3_M2  M3_M2_979
timestamp 1745462530
transform 1 0 3524 0 1 3375
box -3 -3 3 3
use M3_M2  M3_M2_980
timestamp 1745462530
transform 1 0 3492 0 1 3055
box -3 -3 3 3
use M3_M2  M3_M2_981
timestamp 1745462530
transform 1 0 3404 0 1 3585
box -3 -3 3 3
use M3_M2  M3_M2_982
timestamp 1745462530
transform 1 0 3404 0 1 3475
box -3 -3 3 3
use M3_M2  M3_M2_983
timestamp 1745462530
transform 1 0 3364 0 1 3055
box -3 -3 3 3
use M3_M2  M3_M2_984
timestamp 1745462530
transform 1 0 3348 0 1 3475
box -3 -3 3 3
use M3_M2  M3_M2_985
timestamp 1745462530
transform 1 0 3348 0 1 3445
box -3 -3 3 3
use M3_M2  M3_M2_986
timestamp 1745462530
transform 1 0 3276 0 1 3585
box -3 -3 3 3
use M3_M2  M3_M2_987
timestamp 1745462530
transform 1 0 3228 0 1 3445
box -3 -3 3 3
use M3_M2  M3_M2_988
timestamp 1745462530
transform 1 0 1644 0 1 3445
box -3 -3 3 3
use M3_M2  M3_M2_989
timestamp 1745462530
transform 1 0 2900 0 1 3465
box -3 -3 3 3
use M3_M2  M3_M2_990
timestamp 1745462530
transform 1 0 2812 0 1 3465
box -3 -3 3 3
use M3_M2  M3_M2_991
timestamp 1745462530
transform 1 0 2732 0 1 3665
box -3 -3 3 3
use M3_M2  M3_M2_992
timestamp 1745462530
transform 1 0 2708 0 1 3665
box -3 -3 3 3
use M3_M2  M3_M2_993
timestamp 1745462530
transform 1 0 2668 0 1 3955
box -3 -3 3 3
use M3_M2  M3_M2_994
timestamp 1745462530
transform 1 0 2500 0 1 4085
box -3 -3 3 3
use M3_M2  M3_M2_995
timestamp 1745462530
transform 1 0 2500 0 1 3955
box -3 -3 3 3
use M3_M2  M3_M2_996
timestamp 1745462530
transform 1 0 1588 0 1 3485
box -3 -3 3 3
use M3_M2  M3_M2_997
timestamp 1745462530
transform 1 0 1564 0 1 3225
box -3 -3 3 3
use M3_M2  M3_M2_998
timestamp 1745462530
transform 1 0 1500 0 1 3225
box -3 -3 3 3
use M3_M2  M3_M2_999
timestamp 1745462530
transform 1 0 1484 0 1 4085
box -3 -3 3 3
use M3_M2  M3_M2_1000
timestamp 1745462530
transform 1 0 1484 0 1 3485
box -3 -3 3 3
use M3_M2  M3_M2_1001
timestamp 1745462530
transform 1 0 1636 0 1 3585
box -3 -3 3 3
use M3_M2  M3_M2_1002
timestamp 1745462530
transform 1 0 1620 0 1 3045
box -3 -3 3 3
use M3_M2  M3_M2_1003
timestamp 1745462530
transform 1 0 1604 0 1 3585
box -3 -3 3 3
use M3_M2  M3_M2_1004
timestamp 1745462530
transform 1 0 1580 0 1 3045
box -3 -3 3 3
use M3_M2  M3_M2_1005
timestamp 1745462530
transform 1 0 1532 0 1 3165
box -3 -3 3 3
use M3_M2  M3_M2_1006
timestamp 1745462530
transform 1 0 1452 0 1 3585
box -3 -3 3 3
use M3_M2  M3_M2_1007
timestamp 1745462530
transform 1 0 1452 0 1 3165
box -3 -3 3 3
use M3_M2  M3_M2_1008
timestamp 1745462530
transform 1 0 1420 0 1 3585
box -3 -3 3 3
use M3_M2  M3_M2_1009
timestamp 1745462530
transform 1 0 1420 0 1 3165
box -3 -3 3 3
use M3_M2  M3_M2_1010
timestamp 1745462530
transform 1 0 1836 0 1 3715
box -3 -3 3 3
use M3_M2  M3_M2_1011
timestamp 1745462530
transform 1 0 1788 0 1 3715
box -3 -3 3 3
use M3_M2  M3_M2_1012
timestamp 1745462530
transform 1 0 1676 0 1 3665
box -3 -3 3 3
use M3_M2  M3_M2_1013
timestamp 1745462530
transform 1 0 1660 0 1 3665
box -3 -3 3 3
use M3_M2  M3_M2_1014
timestamp 1745462530
transform 1 0 1588 0 1 3665
box -3 -3 3 3
use M3_M2  M3_M2_1015
timestamp 1745462530
transform 1 0 1428 0 1 3665
box -3 -3 3 3
use M3_M2  M3_M2_1016
timestamp 1745462530
transform 1 0 1324 0 1 2975
box -3 -3 3 3
use M3_M2  M3_M2_1017
timestamp 1745462530
transform 1 0 1308 0 1 3315
box -3 -3 3 3
use M3_M2  M3_M2_1018
timestamp 1745462530
transform 1 0 1284 0 1 3665
box -3 -3 3 3
use M3_M2  M3_M2_1019
timestamp 1745462530
transform 1 0 1252 0 1 3315
box -3 -3 3 3
use M3_M2  M3_M2_1020
timestamp 1745462530
transform 1 0 1252 0 1 2975
box -3 -3 3 3
use M3_M2  M3_M2_1021
timestamp 1745462530
transform 1 0 628 0 1 3235
box -3 -3 3 3
use M3_M2  M3_M2_1022
timestamp 1745462530
transform 1 0 572 0 1 3225
box -3 -3 3 3
use M3_M2  M3_M2_1023
timestamp 1745462530
transform 1 0 468 0 1 3225
box -3 -3 3 3
use M3_M2  M3_M2_1024
timestamp 1745462530
transform 1 0 468 0 1 3185
box -3 -3 3 3
use M3_M2  M3_M2_1025
timestamp 1745462530
transform 1 0 372 0 1 3185
box -3 -3 3 3
use M3_M2  M3_M2_1026
timestamp 1745462530
transform 1 0 260 0 1 3185
box -3 -3 3 3
use M3_M2  M3_M2_1027
timestamp 1745462530
transform 1 0 188 0 1 3225
box -3 -3 3 3
use M3_M2  M3_M2_1028
timestamp 1745462530
transform 1 0 140 0 1 3225
box -3 -3 3 3
use M3_M2  M3_M2_1029
timestamp 1745462530
transform 1 0 188 0 1 3115
box -3 -3 3 3
use M3_M2  M3_M2_1030
timestamp 1745462530
transform 1 0 148 0 1 3115
box -3 -3 3 3
use M3_M2  M3_M2_1031
timestamp 1745462530
transform 1 0 1844 0 1 3515
box -3 -3 3 3
use M3_M2  M3_M2_1032
timestamp 1745462530
transform 1 0 1844 0 1 3375
box -3 -3 3 3
use M3_M2  M3_M2_1033
timestamp 1745462530
transform 1 0 1772 0 1 3525
box -3 -3 3 3
use M3_M2  M3_M2_1034
timestamp 1745462530
transform 1 0 1748 0 1 3225
box -3 -3 3 3
use M3_M2  M3_M2_1035
timestamp 1745462530
transform 1 0 1740 0 1 3205
box -3 -3 3 3
use M3_M2  M3_M2_1036
timestamp 1745462530
transform 1 0 1740 0 1 3075
box -3 -3 3 3
use M3_M2  M3_M2_1037
timestamp 1745462530
transform 1 0 1732 0 1 3375
box -3 -3 3 3
use M3_M2  M3_M2_1038
timestamp 1745462530
transform 1 0 1716 0 1 3525
box -3 -3 3 3
use M3_M2  M3_M2_1039
timestamp 1745462530
transform 1 0 1692 0 1 3375
box -3 -3 3 3
use M3_M2  M3_M2_1040
timestamp 1745462530
transform 1 0 1636 0 1 3075
box -3 -3 3 3
use M3_M2  M3_M2_1041
timestamp 1745462530
transform 1 0 1628 0 1 3375
box -3 -3 3 3
use M3_M2  M3_M2_1042
timestamp 1745462530
transform 1 0 1028 0 1 2805
box -3 -3 3 3
use M3_M2  M3_M2_1043
timestamp 1745462530
transform 1 0 988 0 1 2805
box -3 -3 3 3
use M3_M2  M3_M2_1044
timestamp 1745462530
transform 1 0 988 0 1 2765
box -3 -3 3 3
use M3_M2  M3_M2_1045
timestamp 1745462530
transform 1 0 884 0 1 2765
box -3 -3 3 3
use M3_M2  M3_M2_1046
timestamp 1745462530
transform 1 0 1268 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_1047
timestamp 1745462530
transform 1 0 1204 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_1048
timestamp 1745462530
transform 1 0 1204 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_1049
timestamp 1745462530
transform 1 0 1164 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_1050
timestamp 1745462530
transform 1 0 1260 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_1051
timestamp 1745462530
transform 1 0 1220 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_1052
timestamp 1745462530
transform 1 0 1284 0 1 2575
box -3 -3 3 3
use M3_M2  M3_M2_1053
timestamp 1745462530
transform 1 0 1260 0 1 2715
box -3 -3 3 3
use M3_M2  M3_M2_1054
timestamp 1745462530
transform 1 0 1260 0 1 2575
box -3 -3 3 3
use M3_M2  M3_M2_1055
timestamp 1745462530
transform 1 0 1220 0 1 2715
box -3 -3 3 3
use M3_M2  M3_M2_1056
timestamp 1745462530
transform 1 0 1228 0 1 2165
box -3 -3 3 3
use M3_M2  M3_M2_1057
timestamp 1745462530
transform 1 0 1212 0 1 2165
box -3 -3 3 3
use M3_M2  M3_M2_1058
timestamp 1745462530
transform 1 0 1140 0 1 2165
box -3 -3 3 3
use M3_M2  M3_M2_1059
timestamp 1745462530
transform 1 0 1212 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_1060
timestamp 1745462530
transform 1 0 1164 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_1061
timestamp 1745462530
transform 1 0 1188 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_1062
timestamp 1745462530
transform 1 0 1156 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_1063
timestamp 1745462530
transform 1 0 868 0 1 2645
box -3 -3 3 3
use M3_M2  M3_M2_1064
timestamp 1745462530
transform 1 0 860 0 1 2835
box -3 -3 3 3
use M3_M2  M3_M2_1065
timestamp 1745462530
transform 1 0 836 0 1 2835
box -3 -3 3 3
use M3_M2  M3_M2_1066
timestamp 1745462530
transform 1 0 828 0 1 2645
box -3 -3 3 3
use M3_M2  M3_M2_1067
timestamp 1745462530
transform 1 0 900 0 1 2675
box -3 -3 3 3
use M3_M2  M3_M2_1068
timestamp 1745462530
transform 1 0 884 0 1 2885
box -3 -3 3 3
use M3_M2  M3_M2_1069
timestamp 1745462530
transform 1 0 868 0 1 2675
box -3 -3 3 3
use M3_M2  M3_M2_1070
timestamp 1745462530
transform 1 0 244 0 1 2765
box -3 -3 3 3
use M3_M2  M3_M2_1071
timestamp 1745462530
transform 1 0 188 0 1 2885
box -3 -3 3 3
use M3_M2  M3_M2_1072
timestamp 1745462530
transform 1 0 188 0 1 2765
box -3 -3 3 3
use M3_M2  M3_M2_1073
timestamp 1745462530
transform 1 0 220 0 1 2335
box -3 -3 3 3
use M3_M2  M3_M2_1074
timestamp 1745462530
transform 1 0 172 0 1 2335
box -3 -3 3 3
use M3_M2  M3_M2_1075
timestamp 1745462530
transform 1 0 236 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_1076
timestamp 1745462530
transform 1 0 196 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_1077
timestamp 1745462530
transform 1 0 572 0 1 1035
box -3 -3 3 3
use M3_M2  M3_M2_1078
timestamp 1745462530
transform 1 0 300 0 1 1035
box -3 -3 3 3
use M3_M2  M3_M2_1079
timestamp 1745462530
transform 1 0 292 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_1080
timestamp 1745462530
transform 1 0 252 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_1081
timestamp 1745462530
transform 1 0 196 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_1082
timestamp 1745462530
transform 1 0 660 0 1 845
box -3 -3 3 3
use M3_M2  M3_M2_1083
timestamp 1745462530
transform 1 0 340 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_1084
timestamp 1745462530
transform 1 0 340 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_1085
timestamp 1745462530
transform 1 0 308 0 1 845
box -3 -3 3 3
use M3_M2  M3_M2_1086
timestamp 1745462530
transform 1 0 308 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_1087
timestamp 1745462530
transform 1 0 260 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_1088
timestamp 1745462530
transform 1 0 220 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_1089
timestamp 1745462530
transform 1 0 308 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_1090
timestamp 1745462530
transform 1 0 236 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_1091
timestamp 1745462530
transform 1 0 748 0 1 575
box -3 -3 3 3
use M3_M2  M3_M2_1092
timestamp 1745462530
transform 1 0 708 0 1 575
box -3 -3 3 3
use M3_M2  M3_M2_1093
timestamp 1745462530
transform 1 0 236 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_1094
timestamp 1745462530
transform 1 0 204 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_1095
timestamp 1745462530
transform 1 0 1196 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_1096
timestamp 1745462530
transform 1 0 1156 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_1097
timestamp 1745462530
transform 1 0 1100 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_1098
timestamp 1745462530
transform 1 0 1100 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_1099
timestamp 1745462530
transform 1 0 1332 0 1 535
box -3 -3 3 3
use M3_M2  M3_M2_1100
timestamp 1745462530
transform 1 0 1204 0 1 535
box -3 -3 3 3
use M3_M2  M3_M2_1101
timestamp 1745462530
transform 1 0 1140 0 1 535
box -3 -3 3 3
use M3_M2  M3_M2_1102
timestamp 1745462530
transform 1 0 1372 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_1103
timestamp 1745462530
transform 1 0 1316 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_1104
timestamp 1745462530
transform 1 0 1452 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_1105
timestamp 1745462530
transform 1 0 1420 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_1106
timestamp 1745462530
transform 1 0 1444 0 1 975
box -3 -3 3 3
use M3_M2  M3_M2_1107
timestamp 1745462530
transform 1 0 1404 0 1 975
box -3 -3 3 3
use M3_M2  M3_M2_1108
timestamp 1745462530
transform 1 0 1484 0 1 1335
box -3 -3 3 3
use M3_M2  M3_M2_1109
timestamp 1745462530
transform 1 0 1420 0 1 1335
box -3 -3 3 3
use M3_M2  M3_M2_1110
timestamp 1745462530
transform 1 0 1548 0 1 1415
box -3 -3 3 3
use M3_M2  M3_M2_1111
timestamp 1745462530
transform 1 0 1508 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_1112
timestamp 1745462530
transform 1 0 2324 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_1113
timestamp 1745462530
transform 1 0 2228 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_1114
timestamp 1745462530
transform 1 0 2476 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_1115
timestamp 1745462530
transform 1 0 2396 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_1116
timestamp 1745462530
transform 1 0 2396 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_1117
timestamp 1745462530
transform 1 0 2324 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_1118
timestamp 1745462530
transform 1 0 2204 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_1119
timestamp 1745462530
transform 1 0 2428 0 1 535
box -3 -3 3 3
use M3_M2  M3_M2_1120
timestamp 1745462530
transform 1 0 2348 0 1 535
box -3 -3 3 3
use M3_M2  M3_M2_1121
timestamp 1745462530
transform 1 0 2628 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_1122
timestamp 1745462530
transform 1 0 2596 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_1123
timestamp 1745462530
transform 1 0 3468 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_1124
timestamp 1745462530
transform 1 0 3428 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_1125
timestamp 1745462530
transform 1 0 3340 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_1126
timestamp 1745462530
transform 1 0 3548 0 1 455
box -3 -3 3 3
use M3_M2  M3_M2_1127
timestamp 1745462530
transform 1 0 3452 0 1 455
box -3 -3 3 3
use M3_M2  M3_M2_1128
timestamp 1745462530
transform 1 0 4012 0 1 495
box -3 -3 3 3
use M3_M2  M3_M2_1129
timestamp 1745462530
transform 1 0 3980 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_1130
timestamp 1745462530
transform 1 0 3980 0 1 495
box -3 -3 3 3
use M3_M2  M3_M2_1131
timestamp 1745462530
transform 1 0 3588 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_1132
timestamp 1745462530
transform 1 0 3444 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_1133
timestamp 1745462530
transform 1 0 3972 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_1134
timestamp 1745462530
transform 1 0 3940 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_1135
timestamp 1745462530
transform 1 0 3476 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_1136
timestamp 1745462530
transform 1 0 3428 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_1137
timestamp 1745462530
transform 1 0 4116 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_1138
timestamp 1745462530
transform 1 0 3964 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_1139
timestamp 1745462530
transform 1 0 3948 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_1140
timestamp 1745462530
transform 1 0 3564 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_1141
timestamp 1745462530
transform 1 0 3564 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_1142
timestamp 1745462530
transform 1 0 3532 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_1143
timestamp 1745462530
transform 1 0 4140 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_1144
timestamp 1745462530
transform 1 0 4100 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_1145
timestamp 1745462530
transform 1 0 3668 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_1146
timestamp 1745462530
transform 1 0 3596 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_1147
timestamp 1745462530
transform 1 0 3708 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_1148
timestamp 1745462530
transform 1 0 3620 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_1149
timestamp 1745462530
transform 1 0 3404 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_1150
timestamp 1745462530
transform 1 0 3356 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_1151
timestamp 1745462530
transform 1 0 2652 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_1152
timestamp 1745462530
transform 1 0 2612 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_1153
timestamp 1745462530
transform 1 0 3540 0 1 2775
box -3 -3 3 3
use M3_M2  M3_M2_1154
timestamp 1745462530
transform 1 0 3420 0 1 2785
box -3 -3 3 3
use M3_M2  M3_M2_1155
timestamp 1745462530
transform 1 0 3484 0 1 2435
box -3 -3 3 3
use M3_M2  M3_M2_1156
timestamp 1745462530
transform 1 0 3452 0 1 2435
box -3 -3 3 3
use M3_M2  M3_M2_1157
timestamp 1745462530
transform 1 0 3284 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_1158
timestamp 1745462530
transform 1 0 3236 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_1159
timestamp 1745462530
transform 1 0 3044 0 1 3025
box -3 -3 3 3
use M3_M2  M3_M2_1160
timestamp 1745462530
transform 1 0 2964 0 1 3045
box -3 -3 3 3
use M3_M2  M3_M2_1161
timestamp 1745462530
transform 1 0 2964 0 1 3025
box -3 -3 3 3
use M3_M2  M3_M2_1162
timestamp 1745462530
transform 1 0 2876 0 1 3045
box -3 -3 3 3
use M3_M2  M3_M2_1163
timestamp 1745462530
transform 1 0 2716 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_1164
timestamp 1745462530
transform 1 0 2692 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_1165
timestamp 1745462530
transform 1 0 900 0 1 2805
box -3 -3 3 3
use M3_M2  M3_M2_1166
timestamp 1745462530
transform 1 0 868 0 1 2805
box -3 -3 3 3
use M3_M2  M3_M2_1167
timestamp 1745462530
transform 1 0 1812 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_1168
timestamp 1745462530
transform 1 0 1796 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_1169
timestamp 1745462530
transform 1 0 1764 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_1170
timestamp 1745462530
transform 1 0 1828 0 1 1975
box -3 -3 3 3
use M3_M2  M3_M2_1171
timestamp 1745462530
transform 1 0 1748 0 1 1975
box -3 -3 3 3
use M3_M2  M3_M2_1172
timestamp 1745462530
transform 1 0 884 0 1 2785
box -3 -3 3 3
use M3_M2  M3_M2_1173
timestamp 1745462530
transform 1 0 820 0 1 2785
box -3 -3 3 3
use M3_M2  M3_M2_1174
timestamp 1745462530
transform 1 0 500 0 1 2785
box -3 -3 3 3
use M3_M2  M3_M2_1175
timestamp 1745462530
transform 1 0 468 0 1 2785
box -3 -3 3 3
use M3_M2  M3_M2_1176
timestamp 1745462530
transform 1 0 756 0 1 655
box -3 -3 3 3
use M3_M2  M3_M2_1177
timestamp 1745462530
transform 1 0 380 0 1 1465
box -3 -3 3 3
use M3_M2  M3_M2_1178
timestamp 1745462530
transform 1 0 340 0 1 1075
box -3 -3 3 3
use M3_M2  M3_M2_1179
timestamp 1745462530
transform 1 0 316 0 1 1465
box -3 -3 3 3
use M3_M2  M3_M2_1180
timestamp 1745462530
transform 1 0 316 0 1 655
box -3 -3 3 3
use M3_M2  M3_M2_1181
timestamp 1745462530
transform 1 0 172 0 1 655
box -3 -3 3 3
use M3_M2  M3_M2_1182
timestamp 1745462530
transform 1 0 164 0 1 1075
box -3 -3 3 3
use M3_M2  M3_M2_1183
timestamp 1745462530
transform 1 0 284 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_1184
timestamp 1745462530
transform 1 0 252 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_1185
timestamp 1745462530
transform 1 0 228 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_1186
timestamp 1745462530
transform 1 0 804 0 1 495
box -3 -3 3 3
use M3_M2  M3_M2_1187
timestamp 1745462530
transform 1 0 324 0 1 495
box -3 -3 3 3
use M3_M2  M3_M2_1188
timestamp 1745462530
transform 1 0 308 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_1189
timestamp 1745462530
transform 1 0 228 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_1190
timestamp 1745462530
transform 1 0 188 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_1191
timestamp 1745462530
transform 1 0 284 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_1192
timestamp 1745462530
transform 1 0 252 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_1193
timestamp 1745462530
transform 1 0 220 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_1194
timestamp 1745462530
transform 1 0 180 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_1195
timestamp 1745462530
transform 1 0 1988 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_1196
timestamp 1745462530
transform 1 0 1940 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_1197
timestamp 1745462530
transform 1 0 1644 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_1198
timestamp 1745462530
transform 1 0 2076 0 1 495
box -3 -3 3 3
use M3_M2  M3_M2_1199
timestamp 1745462530
transform 1 0 1948 0 1 495
box -3 -3 3 3
use M3_M2  M3_M2_1200
timestamp 1745462530
transform 1 0 2036 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_1201
timestamp 1745462530
transform 1 0 1964 0 1 605
box -3 -3 3 3
use M3_M2  M3_M2_1202
timestamp 1745462530
transform 1 0 2028 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_1203
timestamp 1745462530
transform 1 0 1972 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_1204
timestamp 1745462530
transform 1 0 2108 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_1205
timestamp 1745462530
transform 1 0 2052 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_1206
timestamp 1745462530
transform 1 0 2500 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_1207
timestamp 1745462530
transform 1 0 2404 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_1208
timestamp 1745462530
transform 1 0 2452 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_1209
timestamp 1745462530
transform 1 0 2316 0 1 725
box -3 -3 3 3
use M3_M2  M3_M2_1210
timestamp 1745462530
transform 1 0 2492 0 1 485
box -3 -3 3 3
use M3_M2  M3_M2_1211
timestamp 1745462530
transform 1 0 2356 0 1 485
box -3 -3 3 3
use M3_M2  M3_M2_1212
timestamp 1745462530
transform 1 0 2548 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_1213
timestamp 1745462530
transform 1 0 2500 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_1214
timestamp 1745462530
transform 1 0 2628 0 1 1065
box -3 -3 3 3
use M3_M2  M3_M2_1215
timestamp 1745462530
transform 1 0 2588 0 1 1065
box -3 -3 3 3
use M3_M2  M3_M2_1216
timestamp 1745462530
transform 1 0 2628 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_1217
timestamp 1745462530
transform 1 0 2588 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_1218
timestamp 1745462530
transform 1 0 3684 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_1219
timestamp 1745462530
transform 1 0 3628 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_1220
timestamp 1745462530
transform 1 0 3628 0 1 335
box -3 -3 3 3
use M3_M2  M3_M2_1221
timestamp 1745462530
transform 1 0 3532 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_1222
timestamp 1745462530
transform 1 0 3420 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_1223
timestamp 1745462530
transform 1 0 3764 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_1224
timestamp 1745462530
transform 1 0 3644 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_1225
timestamp 1745462530
transform 1 0 3612 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_1226
timestamp 1745462530
transform 1 0 4244 0 1 465
box -3 -3 3 3
use M3_M2  M3_M2_1227
timestamp 1745462530
transform 1 0 3732 0 1 465
box -3 -3 3 3
use M3_M2  M3_M2_1228
timestamp 1745462530
transform 1 0 3804 0 1 645
box -3 -3 3 3
use M3_M2  M3_M2_1229
timestamp 1745462530
transform 1 0 3700 0 1 645
box -3 -3 3 3
use M3_M2  M3_M2_1230
timestamp 1745462530
transform 1 0 4180 0 1 815
box -3 -3 3 3
use M3_M2  M3_M2_1231
timestamp 1745462530
transform 1 0 4132 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_1232
timestamp 1745462530
transform 1 0 3828 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_1233
timestamp 1745462530
transform 1 0 3788 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_1234
timestamp 1745462530
transform 1 0 3804 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_1235
timestamp 1745462530
transform 1 0 3764 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_1236
timestamp 1745462530
transform 1 0 4180 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_1237
timestamp 1745462530
transform 1 0 3900 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_1238
timestamp 1745462530
transform 1 0 3748 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_1239
timestamp 1745462530
transform 1 0 4244 0 1 1435
box -3 -3 3 3
use M3_M2  M3_M2_1240
timestamp 1745462530
transform 1 0 3900 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_1241
timestamp 1745462530
transform 1 0 3788 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_1242
timestamp 1745462530
transform 1 0 3876 0 1 1535
box -3 -3 3 3
use M3_M2  M3_M2_1243
timestamp 1745462530
transform 1 0 3852 0 1 1535
box -3 -3 3 3
use M3_M2  M3_M2_1244
timestamp 1745462530
transform 1 0 3836 0 1 1535
box -3 -3 3 3
use M3_M2  M3_M2_1245
timestamp 1745462530
transform 1 0 4012 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_1246
timestamp 1745462530
transform 1 0 3940 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_1247
timestamp 1745462530
transform 1 0 3892 0 1 2755
box -3 -3 3 3
use M3_M2  M3_M2_1248
timestamp 1745462530
transform 1 0 3804 0 1 2755
box -3 -3 3 3
use M3_M2  M3_M2_1249
timestamp 1745462530
transform 1 0 3772 0 1 2755
box -3 -3 3 3
use M3_M2  M3_M2_1250
timestamp 1745462530
transform 1 0 3884 0 1 2765
box -3 -3 3 3
use M3_M2  M3_M2_1251
timestamp 1745462530
transform 1 0 3844 0 1 2765
box -3 -3 3 3
use M3_M2  M3_M2_1252
timestamp 1745462530
transform 1 0 3820 0 1 2765
box -3 -3 3 3
use M3_M2  M3_M2_1253
timestamp 1745462530
transform 1 0 3908 0 1 2475
box -3 -3 3 3
use M3_M2  M3_M2_1254
timestamp 1745462530
transform 1 0 3868 0 1 2545
box -3 -3 3 3
use M3_M2  M3_M2_1255
timestamp 1745462530
transform 1 0 3868 0 1 2475
box -3 -3 3 3
use M3_M2  M3_M2_1256
timestamp 1745462530
transform 1 0 3820 0 1 2545
box -3 -3 3 3
use M3_M2  M3_M2_1257
timestamp 1745462530
transform 1 0 3956 0 1 2355
box -3 -3 3 3
use M3_M2  M3_M2_1258
timestamp 1745462530
transform 1 0 3900 0 1 2355
box -3 -3 3 3
use M3_M2  M3_M2_1259
timestamp 1745462530
transform 1 0 3868 0 1 3035
box -3 -3 3 3
use M3_M2  M3_M2_1260
timestamp 1745462530
transform 1 0 3836 0 1 3035
box -3 -3 3 3
use M3_M2  M3_M2_1261
timestamp 1745462530
transform 1 0 3012 0 1 3065
box -3 -3 3 3
use M3_M2  M3_M2_1262
timestamp 1745462530
transform 1 0 2924 0 1 3065
box -3 -3 3 3
use M3_M2  M3_M2_1263
timestamp 1745462530
transform 1 0 2884 0 1 3095
box -3 -3 3 3
use M3_M2  M3_M2_1264
timestamp 1745462530
transform 1 0 2844 0 1 3095
box -3 -3 3 3
use M3_M2  M3_M2_1265
timestamp 1745462530
transform 1 0 988 0 1 2625
box -3 -3 3 3
use M3_M2  M3_M2_1266
timestamp 1745462530
transform 1 0 916 0 1 2625
box -3 -3 3 3
use M3_M2  M3_M2_1267
timestamp 1745462530
transform 1 0 724 0 1 2625
box -3 -3 3 3
use M3_M2  M3_M2_1268
timestamp 1745462530
transform 1 0 1772 0 1 2835
box -3 -3 3 3
use M3_M2  M3_M2_1269
timestamp 1745462530
transform 1 0 1700 0 1 2835
box -3 -3 3 3
use M3_M2  M3_M2_1270
timestamp 1745462530
transform 1 0 1732 0 1 2185
box -3 -3 3 3
use M3_M2  M3_M2_1271
timestamp 1745462530
transform 1 0 1668 0 1 2185
box -3 -3 3 3
use M3_M2  M3_M2_1272
timestamp 1745462530
transform 1 0 1764 0 1 2705
box -3 -3 3 3
use M3_M2  M3_M2_1273
timestamp 1745462530
transform 1 0 1764 0 1 2545
box -3 -3 3 3
use M3_M2  M3_M2_1274
timestamp 1745462530
transform 1 0 1708 0 1 2705
box -3 -3 3 3
use M3_M2  M3_M2_1275
timestamp 1745462530
transform 1 0 1668 0 1 2705
box -3 -3 3 3
use M3_M2  M3_M2_1276
timestamp 1745462530
transform 1 0 1668 0 1 2535
box -3 -3 3 3
use M3_M2  M3_M2_1277
timestamp 1745462530
transform 1 0 1676 0 1 2125
box -3 -3 3 3
use M3_M2  M3_M2_1278
timestamp 1745462530
transform 1 0 1620 0 1 2125
box -3 -3 3 3
use M3_M2  M3_M2_1279
timestamp 1745462530
transform 1 0 1588 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_1280
timestamp 1745462530
transform 1 0 1532 0 1 1935
box -3 -3 3 3
use M3_M2  M3_M2_1281
timestamp 1745462530
transform 1 0 652 0 1 2685
box -3 -3 3 3
use M3_M2  M3_M2_1282
timestamp 1745462530
transform 1 0 596 0 1 2685
box -3 -3 3 3
use M3_M2  M3_M2_1283
timestamp 1745462530
transform 1 0 564 0 1 2645
box -3 -3 3 3
use M3_M2  M3_M2_1284
timestamp 1745462530
transform 1 0 452 0 1 2715
box -3 -3 3 3
use M3_M2  M3_M2_1285
timestamp 1745462530
transform 1 0 452 0 1 2645
box -3 -3 3 3
use M3_M2  M3_M2_1286
timestamp 1745462530
transform 1 0 420 0 1 2715
box -3 -3 3 3
use M3_M2  M3_M2_1287
timestamp 1745462530
transform 1 0 636 0 1 2645
box -3 -3 3 3
use M3_M2  M3_M2_1288
timestamp 1745462530
transform 1 0 548 0 1 2635
box -3 -3 3 3
use M3_M2  M3_M2_1289
timestamp 1745462530
transform 1 0 748 0 1 2575
box -3 -3 3 3
use M3_M2  M3_M2_1290
timestamp 1745462530
transform 1 0 604 0 1 2575
box -3 -3 3 3
use M3_M2  M3_M2_1291
timestamp 1745462530
transform 1 0 364 0 1 2575
box -3 -3 3 3
use M3_M2  M3_M2_1292
timestamp 1745462530
transform 1 0 548 0 1 535
box -3 -3 3 3
use M3_M2  M3_M2_1293
timestamp 1745462530
transform 1 0 380 0 1 535
box -3 -3 3 3
use M3_M2  M3_M2_1294
timestamp 1745462530
transform 1 0 380 0 1 455
box -3 -3 3 3
use M3_M2  M3_M2_1295
timestamp 1745462530
transform 1 0 300 0 1 455
box -3 -3 3 3
use M3_M2  M3_M2_1296
timestamp 1745462530
transform 1 0 1876 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_1297
timestamp 1745462530
transform 1 0 1780 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_1298
timestamp 1745462530
transform 1 0 1748 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_1299
timestamp 1745462530
transform 1 0 1852 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_1300
timestamp 1745462530
transform 1 0 1796 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_1301
timestamp 1745462530
transform 1 0 2052 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_1302
timestamp 1745462530
transform 1 0 2012 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_1303
timestamp 1745462530
transform 1 0 2020 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_1304
timestamp 1745462530
transform 1 0 1980 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_1305
timestamp 1745462530
transform 1 0 1956 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_1306
timestamp 1745462530
transform 1 0 1924 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_1307
timestamp 1745462530
transform 1 0 2276 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_1308
timestamp 1745462530
transform 1 0 2260 0 1 325
box -3 -3 3 3
use M3_M2  M3_M2_1309
timestamp 1745462530
transform 1 0 2220 0 1 325
box -3 -3 3 3
use M3_M2  M3_M2_1310
timestamp 1745462530
transform 1 0 2204 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_1311
timestamp 1745462530
transform 1 0 2212 0 1 605
box -3 -3 3 3
use M3_M2  M3_M2_1312
timestamp 1745462530
transform 1 0 2180 0 1 605
box -3 -3 3 3
use M3_M2  M3_M2_1313
timestamp 1745462530
transform 1 0 2412 0 1 465
box -3 -3 3 3
use M3_M2  M3_M2_1314
timestamp 1745462530
transform 1 0 2332 0 1 155
box -3 -3 3 3
use M3_M2  M3_M2_1315
timestamp 1745462530
transform 1 0 2276 0 1 465
box -3 -3 3 3
use M3_M2  M3_M2_1316
timestamp 1745462530
transform 1 0 2276 0 1 155
box -3 -3 3 3
use M3_M2  M3_M2_1317
timestamp 1745462530
transform 1 0 2388 0 1 405
box -3 -3 3 3
use M3_M2  M3_M2_1318
timestamp 1745462530
transform 1 0 2252 0 1 405
box -3 -3 3 3
use M3_M2  M3_M2_1319
timestamp 1745462530
transform 1 0 2220 0 1 405
box -3 -3 3 3
use M3_M2  M3_M2_1320
timestamp 1745462530
transform 1 0 2324 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_1321
timestamp 1745462530
transform 1 0 2284 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_1322
timestamp 1745462530
transform 1 0 2396 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_1323
timestamp 1745462530
transform 1 0 2356 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_1324
timestamp 1745462530
transform 1 0 3828 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_1325
timestamp 1745462530
transform 1 0 3516 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_1326
timestamp 1745462530
transform 1 0 4244 0 1 255
box -3 -3 3 3
use M3_M2  M3_M2_1327
timestamp 1745462530
transform 1 0 4196 0 1 415
box -3 -3 3 3
use M3_M2  M3_M2_1328
timestamp 1745462530
transform 1 0 4196 0 1 255
box -3 -3 3 3
use M3_M2  M3_M2_1329
timestamp 1745462530
transform 1 0 3948 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_1330
timestamp 1745462530
transform 1 0 3940 0 1 415
box -3 -3 3 3
use M3_M2  M3_M2_1331
timestamp 1745462530
transform 1 0 3908 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_1332
timestamp 1745462530
transform 1 0 4268 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_1333
timestamp 1745462530
transform 1 0 4196 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_1334
timestamp 1745462530
transform 1 0 4268 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_1335
timestamp 1745462530
transform 1 0 3604 0 1 1415
box -3 -3 3 3
use M3_M2  M3_M2_1336
timestamp 1745462530
transform 1 0 3516 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_1337
timestamp 1745462530
transform 1 0 3516 0 1 1415
box -3 -3 3 3
use M3_M2  M3_M2_1338
timestamp 1745462530
transform 1 0 3356 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_1339
timestamp 1745462530
transform 1 0 3716 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_1340
timestamp 1745462530
transform 1 0 3644 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_1341
timestamp 1745462530
transform 1 0 3644 0 1 1405
box -3 -3 3 3
use M3_M2  M3_M2_1342
timestamp 1745462530
transform 1 0 3572 0 1 1405
box -3 -3 3 3
use M3_M2  M3_M2_1343
timestamp 1745462530
transform 1 0 4276 0 1 1495
box -3 -3 3 3
use M3_M2  M3_M2_1344
timestamp 1745462530
transform 1 0 3644 0 1 1495
box -3 -3 3 3
use M3_M2  M3_M2_1345
timestamp 1745462530
transform 1 0 3420 0 1 1495
box -3 -3 3 3
use M3_M2  M3_M2_1346
timestamp 1745462530
transform 1 0 3684 0 1 1575
box -3 -3 3 3
use M3_M2  M3_M2_1347
timestamp 1745462530
transform 1 0 3620 0 1 1575
box -3 -3 3 3
use M3_M2  M3_M2_1348
timestamp 1745462530
transform 1 0 4220 0 1 2585
box -3 -3 3 3
use M3_M2  M3_M2_1349
timestamp 1745462530
transform 1 0 4156 0 1 2585
box -3 -3 3 3
use M3_M2  M3_M2_1350
timestamp 1745462530
transform 1 0 4116 0 1 2585
box -3 -3 3 3
use M3_M2  M3_M2_1351
timestamp 1745462530
transform 1 0 4204 0 1 2295
box -3 -3 3 3
use M3_M2  M3_M2_1352
timestamp 1745462530
transform 1 0 4132 0 1 2295
box -3 -3 3 3
use M3_M2  M3_M2_1353
timestamp 1745462530
transform 1 0 4108 0 1 2295
box -3 -3 3 3
use M3_M2  M3_M2_1354
timestamp 1745462530
transform 1 0 2892 0 1 2405
box -3 -3 3 3
use M3_M2  M3_M2_1355
timestamp 1745462530
transform 1 0 2844 0 1 2405
box -3 -3 3 3
use M3_M2  M3_M2_1356
timestamp 1745462530
transform 1 0 2692 0 1 3035
box -3 -3 3 3
use M3_M2  M3_M2_1357
timestamp 1745462530
transform 1 0 2644 0 1 3035
box -3 -3 3 3
use M3_M2  M3_M2_1358
timestamp 1745462530
transform 1 0 2612 0 1 3035
box -3 -3 3 3
use M3_M2  M3_M2_1359
timestamp 1745462530
transform 1 0 2636 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_1360
timestamp 1745462530
transform 1 0 2604 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_1361
timestamp 1745462530
transform 1 0 980 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_1362
timestamp 1745462530
transform 1 0 740 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_1363
timestamp 1745462530
transform 1 0 1388 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_1364
timestamp 1745462530
transform 1 0 1364 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_1365
timestamp 1745462530
transform 1 0 1340 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_1366
timestamp 1745462530
transform 1 0 1324 0 1 2535
box -3 -3 3 3
use M3_M2  M3_M2_1367
timestamp 1745462530
transform 1 0 1292 0 1 2525
box -3 -3 3 3
use M3_M2  M3_M2_1368
timestamp 1745462530
transform 1 0 1292 0 1 2385
box -3 -3 3 3
use M3_M2  M3_M2_1369
timestamp 1745462530
transform 1 0 1276 0 1 2385
box -3 -3 3 3
use M3_M2  M3_M2_1370
timestamp 1745462530
transform 1 0 1316 0 1 2265
box -3 -3 3 3
use M3_M2  M3_M2_1371
timestamp 1745462530
transform 1 0 1316 0 1 2055
box -3 -3 3 3
use M3_M2  M3_M2_1372
timestamp 1745462530
transform 1 0 1292 0 1 2055
box -3 -3 3 3
use M3_M2  M3_M2_1373
timestamp 1745462530
transform 1 0 1260 0 1 2265
box -3 -3 3 3
use M3_M2  M3_M2_1374
timestamp 1745462530
transform 1 0 1260 0 1 2465
box -3 -3 3 3
use M3_M2  M3_M2_1375
timestamp 1745462530
transform 1 0 1220 0 1 2465
box -3 -3 3 3
use M3_M2  M3_M2_1376
timestamp 1745462530
transform 1 0 1276 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_1377
timestamp 1745462530
transform 1 0 1260 0 1 2075
box -3 -3 3 3
use M3_M2  M3_M2_1378
timestamp 1745462530
transform 1 0 1220 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_1379
timestamp 1745462530
transform 1 0 1172 0 1 2185
box -3 -3 3 3
use M3_M2  M3_M2_1380
timestamp 1745462530
transform 1 0 1172 0 1 2075
box -3 -3 3 3
use M3_M2  M3_M2_1381
timestamp 1745462530
transform 1 0 1148 0 1 2185
box -3 -3 3 3
use M3_M2  M3_M2_1382
timestamp 1745462530
transform 1 0 676 0 1 2805
box -3 -3 3 3
use M3_M2  M3_M2_1383
timestamp 1745462530
transform 1 0 580 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_1384
timestamp 1745462530
transform 1 0 412 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_1385
timestamp 1745462530
transform 1 0 372 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_1386
timestamp 1745462530
transform 1 0 756 0 1 2835
box -3 -3 3 3
use M3_M2  M3_M2_1387
timestamp 1745462530
transform 1 0 604 0 1 2835
box -3 -3 3 3
use M3_M2  M3_M2_1388
timestamp 1745462530
transform 1 0 604 0 1 2815
box -3 -3 3 3
use M3_M2  M3_M2_1389
timestamp 1745462530
transform 1 0 316 0 1 2815
box -3 -3 3 3
use M3_M2  M3_M2_1390
timestamp 1745462530
transform 1 0 620 0 1 1375
box -3 -3 3 3
use M3_M2  M3_M2_1391
timestamp 1745462530
transform 1 0 620 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_1392
timestamp 1745462530
transform 1 0 548 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_1393
timestamp 1745462530
transform 1 0 548 0 1 675
box -3 -3 3 3
use M3_M2  M3_M2_1394
timestamp 1745462530
transform 1 0 540 0 1 1375
box -3 -3 3 3
use M3_M2  M3_M2_1395
timestamp 1745462530
transform 1 0 516 0 1 675
box -3 -3 3 3
use M3_M2  M3_M2_1396
timestamp 1745462530
transform 1 0 484 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_1397
timestamp 1745462530
transform 1 0 412 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_1398
timestamp 1745462530
transform 1 0 596 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_1399
timestamp 1745462530
transform 1 0 396 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_1400
timestamp 1745462530
transform 1 0 428 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_1401
timestamp 1745462530
transform 1 0 380 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_1402
timestamp 1745462530
transform 1 0 660 0 1 115
box -3 -3 3 3
use M3_M2  M3_M2_1403
timestamp 1745462530
transform 1 0 628 0 1 115
box -3 -3 3 3
use M3_M2  M3_M2_1404
timestamp 1745462530
transform 1 0 1380 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_1405
timestamp 1745462530
transform 1 0 1188 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_1406
timestamp 1745462530
transform 1 0 1452 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_1407
timestamp 1745462530
transform 1 0 1364 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_1408
timestamp 1745462530
transform 1 0 1476 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_1409
timestamp 1745462530
transform 1 0 1444 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_1410
timestamp 1745462530
transform 1 0 1620 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_1411
timestamp 1745462530
transform 1 0 1572 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_1412
timestamp 1745462530
transform 1 0 1612 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_1413
timestamp 1745462530
transform 1 0 1548 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_1414
timestamp 1745462530
transform 1 0 2948 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_1415
timestamp 1745462530
transform 1 0 2884 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_1416
timestamp 1745462530
transform 1 0 3108 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_1417
timestamp 1745462530
transform 1 0 2924 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_1418
timestamp 1745462530
transform 1 0 2900 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_1419
timestamp 1745462530
transform 1 0 2860 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_1420
timestamp 1745462530
transform 1 0 2828 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_1421
timestamp 1745462530
transform 1 0 2700 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_1422
timestamp 1745462530
transform 1 0 3028 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_1423
timestamp 1745462530
transform 1 0 2844 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_1424
timestamp 1745462530
transform 1 0 2924 0 1 865
box -3 -3 3 3
use M3_M2  M3_M2_1425
timestamp 1745462530
transform 1 0 2892 0 1 865
box -3 -3 3 3
use M3_M2  M3_M2_1426
timestamp 1745462530
transform 1 0 3292 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_1427
timestamp 1745462530
transform 1 0 3292 0 1 325
box -3 -3 3 3
use M3_M2  M3_M2_1428
timestamp 1745462530
transform 1 0 3228 0 1 325
box -3 -3 3 3
use M3_M2  M3_M2_1429
timestamp 1745462530
transform 1 0 3212 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_1430
timestamp 1745462530
transform 1 0 3396 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_1431
timestamp 1745462530
transform 1 0 3244 0 1 535
box -3 -3 3 3
use M3_M2  M3_M2_1432
timestamp 1745462530
transform 1 0 3196 0 1 535
box -3 -3 3 3
use M3_M2  M3_M2_1433
timestamp 1745462530
transform 1 0 4100 0 1 445
box -3 -3 3 3
use M3_M2  M3_M2_1434
timestamp 1745462530
transform 1 0 3388 0 1 495
box -3 -3 3 3
use M3_M2  M3_M2_1435
timestamp 1745462530
transform 1 0 3388 0 1 445
box -3 -3 3 3
use M3_M2  M3_M2_1436
timestamp 1745462530
transform 1 0 3228 0 1 495
box -3 -3 3 3
use M3_M2  M3_M2_1437
timestamp 1745462530
transform 1 0 3388 0 1 605
box -3 -3 3 3
use M3_M2  M3_M2_1438
timestamp 1745462530
transform 1 0 3388 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_1439
timestamp 1745462530
transform 1 0 3364 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_1440
timestamp 1745462530
transform 1 0 3348 0 1 605
box -3 -3 3 3
use M3_M2  M3_M2_1441
timestamp 1745462530
transform 1 0 4084 0 1 815
box -3 -3 3 3
use M3_M2  M3_M2_1442
timestamp 1745462530
transform 1 0 4036 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_1443
timestamp 1745462530
transform 1 0 3420 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_1444
timestamp 1745462530
transform 1 0 3380 0 1 1065
box -3 -3 3 3
use M3_M2  M3_M2_1445
timestamp 1745462530
transform 1 0 3380 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_1446
timestamp 1745462530
transform 1 0 3300 0 1 1055
box -3 -3 3 3
use M3_M2  M3_M2_1447
timestamp 1745462530
transform 1 0 3396 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_1448
timestamp 1745462530
transform 1 0 3340 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_1449
timestamp 1745462530
transform 1 0 4108 0 1 1335
box -3 -3 3 3
use M3_M2  M3_M2_1450
timestamp 1745462530
transform 1 0 4036 0 1 1335
box -3 -3 3 3
use M3_M2  M3_M2_1451
timestamp 1745462530
transform 1 0 3428 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_1452
timestamp 1745462530
transform 1 0 3428 0 1 1335
box -3 -3 3 3
use M3_M2  M3_M2_1453
timestamp 1745462530
transform 1 0 3332 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_1454
timestamp 1745462530
transform 1 0 3540 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_1455
timestamp 1745462530
transform 1 0 3444 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_1456
timestamp 1745462530
transform 1 0 3412 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_1457
timestamp 1745462530
transform 1 0 4092 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_1458
timestamp 1745462530
transform 1 0 4044 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_1459
timestamp 1745462530
transform 1 0 3492 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_1460
timestamp 1745462530
transform 1 0 3356 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_1461
timestamp 1745462530
transform 1 0 3596 0 1 1575
box -3 -3 3 3
use M3_M2  M3_M2_1462
timestamp 1745462530
transform 1 0 3468 0 1 1575
box -3 -3 3 3
use M3_M2  M3_M2_1463
timestamp 1745462530
transform 1 0 3428 0 1 1575
box -3 -3 3 3
use M3_M2  M3_M2_1464
timestamp 1745462530
transform 1 0 4188 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_1465
timestamp 1745462530
transform 1 0 4156 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_1466
timestamp 1745462530
transform 1 0 3308 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_1467
timestamp 1745462530
transform 1 0 3268 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_1468
timestamp 1745462530
transform 1 0 3300 0 1 2695
box -3 -3 3 3
use M3_M2  M3_M2_1469
timestamp 1745462530
transform 1 0 3204 0 1 2695
box -3 -3 3 3
use M3_M2  M3_M2_1470
timestamp 1745462530
transform 1 0 3268 0 1 2805
box -3 -3 3 3
use M3_M2  M3_M2_1471
timestamp 1745462530
transform 1 0 3180 0 1 2805
box -3 -3 3 3
use M3_M2  M3_M2_1472
timestamp 1745462530
transform 1 0 3308 0 1 2455
box -3 -3 3 3
use M3_M2  M3_M2_1473
timestamp 1745462530
transform 1 0 3260 0 1 2455
box -3 -3 3 3
use M3_M2  M3_M2_1474
timestamp 1745462530
transform 1 0 3220 0 1 2455
box -3 -3 3 3
use M3_M2  M3_M2_1475
timestamp 1745462530
transform 1 0 3260 0 1 2385
box -3 -3 3 3
use M3_M2  M3_M2_1476
timestamp 1745462530
transform 1 0 3204 0 1 2385
box -3 -3 3 3
use M3_M2  M3_M2_1477
timestamp 1745462530
transform 1 0 2820 0 1 3025
box -3 -3 3 3
use M3_M2  M3_M2_1478
timestamp 1745462530
transform 1 0 2764 0 1 3045
box -3 -3 3 3
use M3_M2  M3_M2_1479
timestamp 1745462530
transform 1 0 2764 0 1 3025
box -3 -3 3 3
use M3_M2  M3_M2_1480
timestamp 1745462530
transform 1 0 2676 0 1 3085
box -3 -3 3 3
use M3_M2  M3_M2_1481
timestamp 1745462530
transform 1 0 2676 0 1 3045
box -3 -3 3 3
use M3_M2  M3_M2_1482
timestamp 1745462530
transform 1 0 2644 0 1 3085
box -3 -3 3 3
use M3_M2  M3_M2_1483
timestamp 1745462530
transform 1 0 2820 0 1 2715
box -3 -3 3 3
use M3_M2  M3_M2_1484
timestamp 1745462530
transform 1 0 2788 0 1 2715
box -3 -3 3 3
use M3_M2  M3_M2_1485
timestamp 1745462530
transform 1 0 1620 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_1486
timestamp 1745462530
transform 1 0 1580 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_1487
timestamp 1745462530
transform 1 0 1572 0 1 2245
box -3 -3 3 3
use M3_M2  M3_M2_1488
timestamp 1745462530
transform 1 0 1540 0 1 2245
box -3 -3 3 3
use M3_M2  M3_M2_1489
timestamp 1745462530
transform 1 0 1572 0 1 2635
box -3 -3 3 3
use M3_M2  M3_M2_1490
timestamp 1745462530
transform 1 0 1556 0 1 2445
box -3 -3 3 3
use M3_M2  M3_M2_1491
timestamp 1745462530
transform 1 0 1532 0 1 2635
box -3 -3 3 3
use M3_M2  M3_M2_1492
timestamp 1745462530
transform 1 0 1476 0 1 2445
box -3 -3 3 3
use M3_M2  M3_M2_1493
timestamp 1745462530
transform 1 0 1388 0 1 2365
box -3 -3 3 3
use M3_M2  M3_M2_1494
timestamp 1745462530
transform 1 0 1372 0 1 2365
box -3 -3 3 3
use M3_M2  M3_M2_1495
timestamp 1745462530
transform 1 0 1412 0 1 2065
box -3 -3 3 3
use M3_M2  M3_M2_1496
timestamp 1745462530
transform 1 0 1356 0 1 2065
box -3 -3 3 3
use M3_M2  M3_M2_1497
timestamp 1745462530
transform 1 0 740 0 1 2725
box -3 -3 3 3
use M3_M2  M3_M2_1498
timestamp 1745462530
transform 1 0 644 0 1 2725
box -3 -3 3 3
use M3_M2  M3_M2_1499
timestamp 1745462530
transform 1 0 292 0 1 2725
box -3 -3 3 3
use M3_M2  M3_M2_1500
timestamp 1745462530
transform 1 0 292 0 1 2705
box -3 -3 3 3
use M3_M2  M3_M2_1501
timestamp 1745462530
transform 1 0 204 0 1 2705
box -3 -3 3 3
use M3_M2  M3_M2_1502
timestamp 1745462530
transform 1 0 772 0 1 2745
box -3 -3 3 3
use M3_M2  M3_M2_1503
timestamp 1745462530
transform 1 0 724 0 1 2745
box -3 -3 3 3
use M3_M2  M3_M2_1504
timestamp 1745462530
transform 1 0 716 0 1 2845
box -3 -3 3 3
use M3_M2  M3_M2_1505
timestamp 1745462530
transform 1 0 236 0 1 2805
box -3 -3 3 3
use M3_M2  M3_M2_1506
timestamp 1745462530
transform 1 0 204 0 1 2845
box -3 -3 3 3
use M3_M2  M3_M2_1507
timestamp 1745462530
transform 1 0 204 0 1 2805
box -3 -3 3 3
use M3_M2  M3_M2_1508
timestamp 1745462530
transform 1 0 948 0 1 2705
box -3 -3 3 3
use M3_M2  M3_M2_1509
timestamp 1745462530
transform 1 0 700 0 1 2705
box -3 -3 3 3
use M3_M2  M3_M2_1510
timestamp 1745462530
transform 1 0 228 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_1511
timestamp 1745462530
transform 1 0 196 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_1512
timestamp 1745462530
transform 1 0 556 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_1513
timestamp 1745462530
transform 1 0 492 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_1514
timestamp 1745462530
transform 1 0 484 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_1515
timestamp 1745462530
transform 1 0 468 0 1 1535
box -3 -3 3 3
use M3_M2  M3_M2_1516
timestamp 1745462530
transform 1 0 468 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_1517
timestamp 1745462530
transform 1 0 308 0 1 1535
box -3 -3 3 3
use M3_M2  M3_M2_1518
timestamp 1745462530
transform 1 0 204 0 1 1535
box -3 -3 3 3
use M3_M2  M3_M2_1519
timestamp 1745462530
transform 1 0 444 0 1 1005
box -3 -3 3 3
use M3_M2  M3_M2_1520
timestamp 1745462530
transform 1 0 420 0 1 1005
box -3 -3 3 3
use M3_M2  M3_M2_1521
timestamp 1745462530
transform 1 0 564 0 1 685
box -3 -3 3 3
use M3_M2  M3_M2_1522
timestamp 1745462530
transform 1 0 564 0 1 235
box -3 -3 3 3
use M3_M2  M3_M2_1523
timestamp 1745462530
transform 1 0 548 0 1 235
box -3 -3 3 3
use M3_M2  M3_M2_1524
timestamp 1745462530
transform 1 0 532 0 1 685
box -3 -3 3 3
use M3_M2  M3_M2_1525
timestamp 1745462530
transform 1 0 444 0 1 235
box -3 -3 3 3
use M3_M2  M3_M2_1526
timestamp 1745462530
transform 1 0 844 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_1527
timestamp 1745462530
transform 1 0 804 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_1528
timestamp 1745462530
transform 1 0 1132 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_1529
timestamp 1745462530
transform 1 0 1116 0 1 535
box -3 -3 3 3
use M3_M2  M3_M2_1530
timestamp 1745462530
transform 1 0 1076 0 1 535
box -3 -3 3 3
use M3_M2  M3_M2_1531
timestamp 1745462530
transform 1 0 1076 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_1532
timestamp 1745462530
transform 1 0 1060 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_1533
timestamp 1745462530
transform 1 0 1004 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_1534
timestamp 1745462530
transform 1 0 1388 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_1535
timestamp 1745462530
transform 1 0 1268 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_1536
timestamp 1745462530
transform 1 0 1220 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_1537
timestamp 1745462530
transform 1 0 1220 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_1538
timestamp 1745462530
transform 1 0 1084 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_1539
timestamp 1745462530
transform 1 0 1284 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_1540
timestamp 1745462530
transform 1 0 1252 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_1541
timestamp 1745462530
transform 1 0 1444 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_1542
timestamp 1745462530
transform 1 0 1404 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_1543
timestamp 1745462530
transform 1 0 1436 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_1544
timestamp 1745462530
transform 1 0 1396 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_1545
timestamp 1745462530
transform 1 0 2052 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_1546
timestamp 1745462530
transform 1 0 2012 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_1547
timestamp 1745462530
transform 1 0 2788 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_1548
timestamp 1745462530
transform 1 0 2740 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_1549
timestamp 1745462530
transform 1 0 2708 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_1550
timestamp 1745462530
transform 1 0 2740 0 1 495
box -3 -3 3 3
use M3_M2  M3_M2_1551
timestamp 1745462530
transform 1 0 2716 0 1 495
box -3 -3 3 3
use M3_M2  M3_M2_1552
timestamp 1745462530
transform 1 0 2708 0 1 285
box -3 -3 3 3
use M3_M2  M3_M2_1553
timestamp 1745462530
transform 1 0 2652 0 1 285
box -3 -3 3 3
use M3_M2  M3_M2_1554
timestamp 1745462530
transform 1 0 2796 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_1555
timestamp 1745462530
transform 1 0 2732 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_1556
timestamp 1745462530
transform 1 0 3612 0 1 535
box -3 -3 3 3
use M3_M2  M3_M2_1557
timestamp 1745462530
transform 1 0 3588 0 1 535
box -3 -3 3 3
use M3_M2  M3_M2_1558
timestamp 1745462530
transform 1 0 3588 0 1 275
box -3 -3 3 3
use M3_M2  M3_M2_1559
timestamp 1745462530
transform 1 0 3292 0 1 275
box -3 -3 3 3
use M3_M2  M3_M2_1560
timestamp 1745462530
transform 1 0 3612 0 1 285
box -3 -3 3 3
use M3_M2  M3_M2_1561
timestamp 1745462530
transform 1 0 3564 0 1 285
box -3 -3 3 3
use M3_M2  M3_M2_1562
timestamp 1745462530
transform 1 0 3772 0 1 235
box -3 -3 3 3
use M3_M2  M3_M2_1563
timestamp 1745462530
transform 1 0 3692 0 1 235
box -3 -3 3 3
use M3_M2  M3_M2_1564
timestamp 1745462530
transform 1 0 4348 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_1565
timestamp 1745462530
transform 1 0 4268 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_1566
timestamp 1745462530
transform 1 0 4180 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_1567
timestamp 1745462530
transform 1 0 4140 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_1568
timestamp 1745462530
transform 1 0 3636 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_1569
timestamp 1745462530
transform 1 0 3596 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_1570
timestamp 1745462530
transform 1 0 4244 0 1 1815
box -3 -3 3 3
use M3_M2  M3_M2_1571
timestamp 1745462530
transform 1 0 3868 0 1 1855
box -3 -3 3 3
use M3_M2  M3_M2_1572
timestamp 1745462530
transform 1 0 3868 0 1 1815
box -3 -3 3 3
use M3_M2  M3_M2_1573
timestamp 1745462530
transform 1 0 3796 0 1 1935
box -3 -3 3 3
use M3_M2  M3_M2_1574
timestamp 1745462530
transform 1 0 3788 0 1 1855
box -3 -3 3 3
use M3_M2  M3_M2_1575
timestamp 1745462530
transform 1 0 3596 0 1 1935
box -3 -3 3 3
use M3_M2  M3_M2_1576
timestamp 1745462530
transform 1 0 4244 0 1 1865
box -3 -3 3 3
use M3_M2  M3_M2_1577
timestamp 1745462530
transform 1 0 3788 0 1 1865
box -3 -3 3 3
use M3_M2  M3_M2_1578
timestamp 1745462530
transform 1 0 3684 0 1 1865
box -3 -3 3 3
use M3_M2  M3_M2_1579
timestamp 1745462530
transform 1 0 3668 0 1 1865
box -3 -3 3 3
use M3_M2  M3_M2_1580
timestamp 1745462530
transform 1 0 3620 0 1 1865
box -3 -3 3 3
use M3_M2  M3_M2_1581
timestamp 1745462530
transform 1 0 3804 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_1582
timestamp 1745462530
transform 1 0 3740 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_1583
timestamp 1745462530
transform 1 0 3700 0 1 2775
box -3 -3 3 3
use M3_M2  M3_M2_1584
timestamp 1745462530
transform 1 0 3620 0 1 2775
box -3 -3 3 3
use M3_M2  M3_M2_1585
timestamp 1745462530
transform 1 0 3588 0 1 2775
box -3 -3 3 3
use M3_M2  M3_M2_1586
timestamp 1745462530
transform 1 0 3644 0 1 2805
box -3 -3 3 3
use M3_M2  M3_M2_1587
timestamp 1745462530
transform 1 0 3612 0 1 2805
box -3 -3 3 3
use M3_M2  M3_M2_1588
timestamp 1745462530
transform 1 0 3684 0 1 2435
box -3 -3 3 3
use M3_M2  M3_M2_1589
timestamp 1745462530
transform 1 0 3612 0 1 2435
box -3 -3 3 3
use M3_M2  M3_M2_1590
timestamp 1745462530
transform 1 0 3548 0 1 2435
box -3 -3 3 3
use M3_M2  M3_M2_1591
timestamp 1745462530
transform 1 0 3644 0 1 2455
box -3 -3 3 3
use M3_M2  M3_M2_1592
timestamp 1745462530
transform 1 0 3572 0 1 2455
box -3 -3 3 3
use M3_M2  M3_M2_1593
timestamp 1745462530
transform 1 0 3532 0 1 2455
box -3 -3 3 3
use M3_M2  M3_M2_1594
timestamp 1745462530
transform 1 0 3556 0 1 3525
box -3 -3 3 3
use M3_M2  M3_M2_1595
timestamp 1745462530
transform 1 0 3524 0 1 3525
box -3 -3 3 3
use M3_M2  M3_M2_1596
timestamp 1745462530
transform 1 0 3500 0 1 3365
box -3 -3 3 3
use M3_M2  M3_M2_1597
timestamp 1745462530
transform 1 0 3476 0 1 3175
box -3 -3 3 3
use M3_M2  M3_M2_1598
timestamp 1745462530
transform 1 0 3460 0 1 3175
box -3 -3 3 3
use M3_M2  M3_M2_1599
timestamp 1745462530
transform 1 0 3452 0 1 3365
box -3 -3 3 3
use M3_M2  M3_M2_1600
timestamp 1745462530
transform 1 0 3340 0 1 3525
box -3 -3 3 3
use M3_M2  M3_M2_1601
timestamp 1745462530
transform 1 0 3332 0 1 3545
box -3 -3 3 3
use M3_M2  M3_M2_1602
timestamp 1745462530
transform 1 0 3276 0 1 3545
box -3 -3 3 3
use M3_M2  M3_M2_1603
timestamp 1745462530
transform 1 0 3244 0 1 3175
box -3 -3 3 3
use M3_M2  M3_M2_1604
timestamp 1745462530
transform 1 0 3164 0 1 3175
box -3 -3 3 3
use M3_M2  M3_M2_1605
timestamp 1745462530
transform 1 0 3508 0 1 3465
box -3 -3 3 3
use M3_M2  M3_M2_1606
timestamp 1745462530
transform 1 0 3484 0 1 3465
box -3 -3 3 3
use M3_M2  M3_M2_1607
timestamp 1745462530
transform 1 0 3476 0 1 3395
box -3 -3 3 3
use M3_M2  M3_M2_1608
timestamp 1745462530
transform 1 0 3404 0 1 3395
box -3 -3 3 3
use M3_M2  M3_M2_1609
timestamp 1745462530
transform 1 0 3356 0 1 3395
box -3 -3 3 3
use M3_M2  M3_M2_1610
timestamp 1745462530
transform 1 0 3332 0 1 3265
box -3 -3 3 3
use M3_M2  M3_M2_1611
timestamp 1745462530
transform 1 0 3284 0 1 3265
box -3 -3 3 3
use M3_M2  M3_M2_1612
timestamp 1745462530
transform 1 0 3252 0 1 3145
box -3 -3 3 3
use M3_M2  M3_M2_1613
timestamp 1745462530
transform 1 0 3204 0 1 3145
box -3 -3 3 3
use M3_M2  M3_M2_1614
timestamp 1745462530
transform 1 0 2796 0 1 3135
box -3 -3 3 3
use M3_M2  M3_M2_1615
timestamp 1745462530
transform 1 0 2636 0 1 3495
box -3 -3 3 3
use M3_M2  M3_M2_1616
timestamp 1745462530
transform 1 0 2588 0 1 3495
box -3 -3 3 3
use M3_M2  M3_M2_1617
timestamp 1745462530
transform 1 0 2524 0 1 3225
box -3 -3 3 3
use M3_M2  M3_M2_1618
timestamp 1745462530
transform 1 0 2524 0 1 3135
box -3 -3 3 3
use M3_M2  M3_M2_1619
timestamp 1745462530
transform 1 0 2476 0 1 3225
box -3 -3 3 3
use M3_M2  M3_M2_1620
timestamp 1745462530
transform 1 0 2468 0 1 3495
box -3 -3 3 3
use M3_M2  M3_M2_1621
timestamp 1745462530
transform 1 0 2420 0 1 3135
box -3 -3 3 3
use M3_M2  M3_M2_1622
timestamp 1745462530
transform 1 0 2860 0 1 3525
box -3 -3 3 3
use M3_M2  M3_M2_1623
timestamp 1745462530
transform 1 0 2836 0 1 3195
box -3 -3 3 3
use M3_M2  M3_M2_1624
timestamp 1745462530
transform 1 0 2796 0 1 3525
box -3 -3 3 3
use M3_M2  M3_M2_1625
timestamp 1745462530
transform 1 0 2772 0 1 3195
box -3 -3 3 3
use M3_M2  M3_M2_1626
timestamp 1745462530
transform 1 0 2740 0 1 3305
box -3 -3 3 3
use M3_M2  M3_M2_1627
timestamp 1745462530
transform 1 0 2716 0 1 3305
box -3 -3 3 3
use M3_M2  M3_M2_1628
timestamp 1745462530
transform 1 0 2700 0 1 3525
box -3 -3 3 3
use M3_M2  M3_M2_1629
timestamp 1745462530
transform 1 0 3076 0 1 3095
box -3 -3 3 3
use M3_M2  M3_M2_1630
timestamp 1745462530
transform 1 0 3036 0 1 3095
box -3 -3 3 3
use M3_M2  M3_M2_1631
timestamp 1745462530
transform 1 0 2988 0 1 3085
box -3 -3 3 3
use M3_M2  M3_M2_1632
timestamp 1745462530
transform 1 0 2916 0 1 3085
box -3 -3 3 3
use M3_M2  M3_M2_1633
timestamp 1745462530
transform 1 0 3044 0 1 3525
box -3 -3 3 3
use M3_M2  M3_M2_1634
timestamp 1745462530
transform 1 0 3028 0 1 3405
box -3 -3 3 3
use M3_M2  M3_M2_1635
timestamp 1745462530
transform 1 0 3004 0 1 3525
box -3 -3 3 3
use M3_M2  M3_M2_1636
timestamp 1745462530
transform 1 0 2972 0 1 3525
box -3 -3 3 3
use M3_M2  M3_M2_1637
timestamp 1745462530
transform 1 0 2932 0 1 3175
box -3 -3 3 3
use M3_M2  M3_M2_1638
timestamp 1745462530
transform 1 0 2884 0 1 3175
box -3 -3 3 3
use M3_M2  M3_M2_1639
timestamp 1745462530
transform 1 0 2868 0 1 3405
box -3 -3 3 3
use M3_M2  M3_M2_1640
timestamp 1745462530
transform 1 0 2852 0 1 3175
box -3 -3 3 3
use M3_M2  M3_M2_1641
timestamp 1745462530
transform 1 0 3564 0 1 3365
box -3 -3 3 3
use M3_M2  M3_M2_1642
timestamp 1745462530
transform 1 0 3548 0 1 3545
box -3 -3 3 3
use M3_M2  M3_M2_1643
timestamp 1745462530
transform 1 0 3516 0 1 3365
box -3 -3 3 3
use M3_M2  M3_M2_1644
timestamp 1745462530
transform 1 0 3484 0 1 3195
box -3 -3 3 3
use M3_M2  M3_M2_1645
timestamp 1745462530
transform 1 0 3364 0 1 3545
box -3 -3 3 3
use M3_M2  M3_M2_1646
timestamp 1745462530
transform 1 0 3324 0 1 3195
box -3 -3 3 3
use M3_M2  M3_M2_1647
timestamp 1745462530
transform 1 0 3228 0 1 3525
box -3 -3 3 3
use M3_M2  M3_M2_1648
timestamp 1745462530
transform 1 0 3212 0 1 3195
box -3 -3 3 3
use M3_M2  M3_M2_1649
timestamp 1745462530
transform 1 0 3204 0 1 3525
box -3 -3 3 3
use M3_M2  M3_M2_1650
timestamp 1745462530
transform 1 0 3468 0 1 3345
box -3 -3 3 3
use M3_M2  M3_M2_1651
timestamp 1745462530
transform 1 0 3428 0 1 3345
box -3 -3 3 3
use M3_M2  M3_M2_1652
timestamp 1745462530
transform 1 0 3380 0 1 3155
box -3 -3 3 3
use M3_M2  M3_M2_1653
timestamp 1745462530
transform 1 0 3356 0 1 3345
box -3 -3 3 3
use M3_M2  M3_M2_1654
timestamp 1745462530
transform 1 0 3196 0 1 3155
box -3 -3 3 3
use M3_M2  M3_M2_1655
timestamp 1745462530
transform 1 0 3188 0 1 3525
box -3 -3 3 3
use M3_M2  M3_M2_1656
timestamp 1745462530
transform 1 0 3132 0 1 3175
box -3 -3 3 3
use M3_M2  M3_M2_1657
timestamp 1745462530
transform 1 0 3124 0 1 3285
box -3 -3 3 3
use M3_M2  M3_M2_1658
timestamp 1745462530
transform 1 0 3124 0 1 3155
box -3 -3 3 3
use M3_M2  M3_M2_1659
timestamp 1745462530
transform 1 0 3116 0 1 3175
box -3 -3 3 3
use M3_M2  M3_M2_1660
timestamp 1745462530
transform 1 0 3108 0 1 3525
box -3 -3 3 3
use M3_M2  M3_M2_1661
timestamp 1745462530
transform 1 0 3108 0 1 3285
box -3 -3 3 3
use M3_M2  M3_M2_1662
timestamp 1745462530
transform 1 0 2812 0 1 3095
box -3 -3 3 3
use M3_M2  M3_M2_1663
timestamp 1745462530
transform 1 0 2532 0 1 3525
box -3 -3 3 3
use M3_M2  M3_M2_1664
timestamp 1745462530
transform 1 0 2516 0 1 3095
box -3 -3 3 3
use M3_M2  M3_M2_1665
timestamp 1745462530
transform 1 0 2444 0 1 3525
box -3 -3 3 3
use M3_M2  M3_M2_1666
timestamp 1745462530
transform 1 0 2436 0 1 3095
box -3 -3 3 3
use M3_M2  M3_M2_1667
timestamp 1745462530
transform 1 0 2404 0 1 3535
box -3 -3 3 3
use M3_M2  M3_M2_1668
timestamp 1745462530
transform 1 0 2652 0 1 2805
box -3 -3 3 3
use M3_M2  M3_M2_1669
timestamp 1745462530
transform 1 0 2564 0 1 2805
box -3 -3 3 3
use M3_M2  M3_M2_1670
timestamp 1745462530
transform 1 0 1876 0 1 3865
box -3 -3 3 3
use M3_M2  M3_M2_1671
timestamp 1745462530
transform 1 0 1828 0 1 3865
box -3 -3 3 3
use M3_M2  M3_M2_1672
timestamp 1745462530
transform 1 0 1828 0 1 3845
box -3 -3 3 3
use M3_M2  M3_M2_1673
timestamp 1745462530
transform 1 0 1772 0 1 3835
box -3 -3 3 3
use M3_M2  M3_M2_1674
timestamp 1745462530
transform 1 0 1772 0 1 3785
box -3 -3 3 3
use M3_M2  M3_M2_1675
timestamp 1745462530
transform 1 0 1724 0 1 3785
box -3 -3 3 3
use M3_M2  M3_M2_1676
timestamp 1745462530
transform 1 0 1700 0 1 3785
box -3 -3 3 3
use M3_M2  M3_M2_1677
timestamp 1745462530
transform 1 0 1860 0 1 3835
box -3 -3 3 3
use M3_M2  M3_M2_1678
timestamp 1745462530
transform 1 0 1812 0 1 3835
box -3 -3 3 3
use M3_M2  M3_M2_1679
timestamp 1745462530
transform 1 0 1812 0 1 3775
box -3 -3 3 3
use M3_M2  M3_M2_1680
timestamp 1745462530
transform 1 0 1756 0 1 3775
box -3 -3 3 3
use M3_M2  M3_M2_1681
timestamp 1745462530
transform 1 0 2620 0 1 3785
box -3 -3 3 3
use M3_M2  M3_M2_1682
timestamp 1745462530
transform 1 0 2580 0 1 3795
box -3 -3 3 3
use M3_M2  M3_M2_1683
timestamp 1745462530
transform 1 0 2532 0 1 3795
box -3 -3 3 3
use M3_M2  M3_M2_1684
timestamp 1745462530
transform 1 0 2532 0 1 3775
box -3 -3 3 3
use M3_M2  M3_M2_1685
timestamp 1745462530
transform 1 0 2500 0 1 3775
box -3 -3 3 3
use M3_M2  M3_M2_1686
timestamp 1745462530
transform 1 0 2076 0 1 3885
box -3 -3 3 3
use M3_M2  M3_M2_1687
timestamp 1745462530
transform 1 0 2076 0 1 3775
box -3 -3 3 3
use M3_M2  M3_M2_1688
timestamp 1745462530
transform 1 0 2052 0 1 3775
box -3 -3 3 3
use M3_M2  M3_M2_1689
timestamp 1745462530
transform 1 0 2020 0 1 3885
box -3 -3 3 3
use M3_M2  M3_M2_1690
timestamp 1745462530
transform 1 0 2652 0 1 3775
box -3 -3 3 3
use M3_M2  M3_M2_1691
timestamp 1745462530
transform 1 0 2612 0 1 3775
box -3 -3 3 3
use M3_M2  M3_M2_1692
timestamp 1745462530
transform 1 0 2612 0 1 3755
box -3 -3 3 3
use M3_M2  M3_M2_1693
timestamp 1745462530
transform 1 0 2588 0 1 3755
box -3 -3 3 3
use M3_M2  M3_M2_1694
timestamp 1745462530
transform 1 0 2476 0 1 3755
box -3 -3 3 3
use M3_M2  M3_M2_1695
timestamp 1745462530
transform 1 0 2084 0 1 3755
box -3 -3 3 3
use M3_M2  M3_M2_1696
timestamp 1745462530
transform 1 0 2060 0 1 3755
box -3 -3 3 3
use M3_M2  M3_M2_1697
timestamp 1745462530
transform 1 0 1892 0 1 3325
box -3 -3 3 3
use M3_M2  M3_M2_1698
timestamp 1745462530
transform 1 0 1604 0 1 3315
box -3 -3 3 3
use M3_M2  M3_M2_1699
timestamp 1745462530
transform 1 0 1596 0 1 3625
box -3 -3 3 3
use M3_M2  M3_M2_1700
timestamp 1745462530
transform 1 0 1556 0 1 3625
box -3 -3 3 3
use M3_M2  M3_M2_1701
timestamp 1745462530
transform 1 0 1508 0 1 3625
box -3 -3 3 3
use M3_M2  M3_M2_1702
timestamp 1745462530
transform 1 0 1484 0 1 3625
box -3 -3 3 3
use M3_M2  M3_M2_1703
timestamp 1745462530
transform 1 0 3580 0 1 4045
box -3 -3 3 3
use M3_M2  M3_M2_1704
timestamp 1745462530
transform 1 0 3556 0 1 4045
box -3 -3 3 3
use M3_M2  M3_M2_1705
timestamp 1745462530
transform 1 0 3460 0 1 4045
box -3 -3 3 3
use M3_M2  M3_M2_1706
timestamp 1745462530
transform 1 0 3460 0 1 4005
box -3 -3 3 3
use M3_M2  M3_M2_1707
timestamp 1745462530
transform 1 0 3076 0 1 4085
box -3 -3 3 3
use M3_M2  M3_M2_1708
timestamp 1745462530
transform 1 0 3076 0 1 4005
box -3 -3 3 3
use M3_M2  M3_M2_1709
timestamp 1745462530
transform 1 0 2700 0 1 4085
box -3 -3 3 3
use M3_M2  M3_M2_1710
timestamp 1745462530
transform 1 0 2692 0 1 4135
box -3 -3 3 3
use M3_M2  M3_M2_1711
timestamp 1745462530
transform 1 0 2644 0 1 4085
box -3 -3 3 3
use M3_M2  M3_M2_1712
timestamp 1745462530
transform 1 0 2372 0 1 4135
box -3 -3 3 3
use M3_M2  M3_M2_1713
timestamp 1745462530
transform 1 0 2268 0 1 4125
box -3 -3 3 3
use M3_M2  M3_M2_1714
timestamp 1745462530
transform 1 0 2260 0 1 4095
box -3 -3 3 3
use M3_M2  M3_M2_1715
timestamp 1745462530
transform 1 0 2148 0 1 4095
box -3 -3 3 3
use M3_M2  M3_M2_1716
timestamp 1745462530
transform 1 0 3524 0 1 3825
box -3 -3 3 3
use M3_M2  M3_M2_1717
timestamp 1745462530
transform 1 0 3476 0 1 3825
box -3 -3 3 3
use M3_M2  M3_M2_1718
timestamp 1745462530
transform 1 0 3236 0 1 3815
box -3 -3 3 3
use M3_M2  M3_M2_1719
timestamp 1745462530
transform 1 0 3044 0 1 3805
box -3 -3 3 3
use M3_M2  M3_M2_1720
timestamp 1745462530
transform 1 0 3044 0 1 3785
box -3 -3 3 3
use M3_M2  M3_M2_1721
timestamp 1745462530
transform 1 0 3036 0 1 3965
box -3 -3 3 3
use M3_M2  M3_M2_1722
timestamp 1745462530
transform 1 0 2916 0 1 3785
box -3 -3 3 3
use M3_M2  M3_M2_1723
timestamp 1745462530
transform 1 0 2916 0 1 3765
box -3 -3 3 3
use M3_M2  M3_M2_1724
timestamp 1745462530
transform 1 0 2764 0 1 3995
box -3 -3 3 3
use M3_M2  M3_M2_1725
timestamp 1745462530
transform 1 0 2764 0 1 3985
box -3 -3 3 3
use M3_M2  M3_M2_1726
timestamp 1745462530
transform 1 0 2668 0 1 3775
box -3 -3 3 3
use M3_M2  M3_M2_1727
timestamp 1745462530
transform 1 0 2316 0 1 3985
box -3 -3 3 3
use M3_M2  M3_M2_1728
timestamp 1745462530
transform 1 0 2156 0 1 3985
box -3 -3 3 3
use M3_M2  M3_M2_1729
timestamp 1745462530
transform 1 0 2156 0 1 3935
box -3 -3 3 3
use M3_M2  M3_M2_1730
timestamp 1745462530
transform 1 0 1980 0 1 3935
box -3 -3 3 3
use M3_M2  M3_M2_1731
timestamp 1745462530
transform 1 0 1980 0 1 3815
box -3 -3 3 3
use M3_M2  M3_M2_1732
timestamp 1745462530
transform 1 0 1884 0 1 3815
box -3 -3 3 3
use M3_M2  M3_M2_1733
timestamp 1745462530
transform 1 0 1884 0 1 3775
box -3 -3 3 3
use M3_M2  M3_M2_1734
timestamp 1745462530
transform 1 0 1828 0 1 3775
box -3 -3 3 3
use M3_M2  M3_M2_1735
timestamp 1745462530
transform 1 0 1980 0 1 2775
box -3 -3 3 3
use M3_M2  M3_M2_1736
timestamp 1745462530
transform 1 0 1924 0 1 2775
box -3 -3 3 3
use M3_M2  M3_M2_1737
timestamp 1745462530
transform 1 0 1988 0 1 2585
box -3 -3 3 3
use M3_M2  M3_M2_1738
timestamp 1745462530
transform 1 0 1924 0 1 2585
box -3 -3 3 3
use M3_M2  M3_M2_1739
timestamp 1745462530
transform 1 0 2004 0 1 2085
box -3 -3 3 3
use M3_M2  M3_M2_1740
timestamp 1745462530
transform 1 0 1980 0 1 2085
box -3 -3 3 3
use M3_M2  M3_M2_1741
timestamp 1745462530
transform 1 0 1836 0 1 2085
box -3 -3 3 3
use M3_M2  M3_M2_1742
timestamp 1745462530
transform 1 0 1828 0 1 2385
box -3 -3 3 3
use M3_M2  M3_M2_1743
timestamp 1745462530
transform 1 0 1772 0 1 2385
box -3 -3 3 3
use M3_M2  M3_M2_1744
timestamp 1745462530
transform 1 0 1772 0 1 2355
box -3 -3 3 3
use M3_M2  M3_M2_1745
timestamp 1745462530
transform 1 0 1732 0 1 2355
box -3 -3 3 3
use M3_M2  M3_M2_1746
timestamp 1745462530
transform 1 0 1852 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_1747
timestamp 1745462530
transform 1 0 1748 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_1748
timestamp 1745462530
transform 1 0 700 0 1 2555
box -3 -3 3 3
use M3_M2  M3_M2_1749
timestamp 1745462530
transform 1 0 636 0 1 2555
box -3 -3 3 3
use M3_M2  M3_M2_1750
timestamp 1745462530
transform 1 0 396 0 1 2555
box -3 -3 3 3
use M3_M2  M3_M2_1751
timestamp 1745462530
transform 1 0 660 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_1752
timestamp 1745462530
transform 1 0 612 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_1753
timestamp 1745462530
transform 1 0 572 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_1754
timestamp 1745462530
transform 1 0 708 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_1755
timestamp 1745462530
transform 1 0 644 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_1756
timestamp 1745462530
transform 1 0 236 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_1757
timestamp 1745462530
transform 1 0 204 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_1758
timestamp 1745462530
transform 1 0 988 0 1 2445
box -3 -3 3 3
use M3_M2  M3_M2_1759
timestamp 1745462530
transform 1 0 908 0 1 2445
box -3 -3 3 3
use M3_M2  M3_M2_1760
timestamp 1745462530
transform 1 0 852 0 1 2435
box -3 -3 3 3
use M3_M2  M3_M2_1761
timestamp 1745462530
transform 1 0 820 0 1 2435
box -3 -3 3 3
use M3_M2  M3_M2_1762
timestamp 1745462530
transform 1 0 700 0 1 2435
box -3 -3 3 3
use M3_M2  M3_M2_1763
timestamp 1745462530
transform 1 0 556 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_1764
timestamp 1745462530
transform 1 0 372 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_1765
timestamp 1745462530
transform 1 0 356 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_1766
timestamp 1745462530
transform 1 0 348 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_1767
timestamp 1745462530
transform 1 0 332 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_1768
timestamp 1745462530
transform 1 0 316 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_1769
timestamp 1745462530
transform 1 0 580 0 1 665
box -3 -3 3 3
use M3_M2  M3_M2_1770
timestamp 1745462530
transform 1 0 492 0 1 685
box -3 -3 3 3
use M3_M2  M3_M2_1771
timestamp 1745462530
transform 1 0 492 0 1 665
box -3 -3 3 3
use M3_M2  M3_M2_1772
timestamp 1745462530
transform 1 0 284 0 1 685
box -3 -3 3 3
use M3_M2  M3_M2_1773
timestamp 1745462530
transform 1 0 620 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_1774
timestamp 1745462530
transform 1 0 492 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_1775
timestamp 1745462530
transform 1 0 732 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_1776
timestamp 1745462530
transform 1 0 700 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_1777
timestamp 1745462530
transform 1 0 1628 0 1 485
box -3 -3 3 3
use M3_M2  M3_M2_1778
timestamp 1745462530
transform 1 0 1508 0 1 485
box -3 -3 3 3
use M3_M2  M3_M2_1779
timestamp 1745462530
transform 1 0 1700 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_1780
timestamp 1745462530
transform 1 0 1612 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_1781
timestamp 1745462530
transform 1 0 1748 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_1782
timestamp 1745462530
transform 1 0 1700 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_1783
timestamp 1745462530
transform 1 0 1812 0 1 1035
box -3 -3 3 3
use M3_M2  M3_M2_1784
timestamp 1745462530
transform 1 0 1764 0 1 1035
box -3 -3 3 3
use M3_M2  M3_M2_1785
timestamp 1745462530
transform 1 0 1860 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_1786
timestamp 1745462530
transform 1 0 1820 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_1787
timestamp 1745462530
transform 1 0 1860 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_1788
timestamp 1745462530
transform 1 0 1764 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_1789
timestamp 1745462530
transform 1 0 2964 0 1 655
box -3 -3 3 3
use M3_M2  M3_M2_1790
timestamp 1745462530
transform 1 0 2924 0 1 655
box -3 -3 3 3
use M3_M2  M3_M2_1791
timestamp 1745462530
transform 1 0 2892 0 1 655
box -3 -3 3 3
use M3_M2  M3_M2_1792
timestamp 1745462530
transform 1 0 3060 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_1793
timestamp 1745462530
transform 1 0 2876 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_1794
timestamp 1745462530
transform 1 0 2948 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_1795
timestamp 1745462530
transform 1 0 2892 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_1796
timestamp 1745462530
transform 1 0 2956 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_1797
timestamp 1745462530
transform 1 0 2940 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_1798
timestamp 1745462530
transform 1 0 3916 0 1 495
box -3 -3 3 3
use M3_M2  M3_M2_1799
timestamp 1745462530
transform 1 0 3780 0 1 495
box -3 -3 3 3
use M3_M2  M3_M2_1800
timestamp 1745462530
transform 1 0 3780 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_1801
timestamp 1745462530
transform 1 0 3380 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_1802
timestamp 1745462530
transform 1 0 3908 0 1 265
box -3 -3 3 3
use M3_M2  M3_M2_1803
timestamp 1745462530
transform 1 0 3764 0 1 265
box -3 -3 3 3
use M3_M2  M3_M2_1804
timestamp 1745462530
transform 1 0 4172 0 1 245
box -3 -3 3 3
use M3_M2  M3_M2_1805
timestamp 1745462530
transform 1 0 4100 0 1 245
box -3 -3 3 3
use M3_M2  M3_M2_1806
timestamp 1745462530
transform 1 0 3932 0 1 245
box -3 -3 3 3
use M3_M2  M3_M2_1807
timestamp 1745462530
transform 1 0 4020 0 1 335
box -3 -3 3 3
use M3_M2  M3_M2_1808
timestamp 1745462530
transform 1 0 3916 0 1 335
box -3 -3 3 3
use M3_M2  M3_M2_1809
timestamp 1745462530
transform 1 0 4180 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_1810
timestamp 1745462530
transform 1 0 4148 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_1811
timestamp 1745462530
transform 1 0 4260 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_1812
timestamp 1745462530
transform 1 0 4132 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_1813
timestamp 1745462530
transform 1 0 4044 0 1 1855
box -3 -3 3 3
use M3_M2  M3_M2_1814
timestamp 1745462530
transform 1 0 4044 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_1815
timestamp 1745462530
transform 1 0 3900 0 1 1855
box -3 -3 3 3
use M3_M2  M3_M2_1816
timestamp 1745462530
transform 1 0 3916 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_1817
timestamp 1745462530
transform 1 0 3884 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_1818
timestamp 1745462530
transform 1 0 4268 0 1 2085
box -3 -3 3 3
use M3_M2  M3_M2_1819
timestamp 1745462530
transform 1 0 4204 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_1820
timestamp 1745462530
transform 1 0 4108 0 1 2085
box -3 -3 3 3
use M3_M2  M3_M2_1821
timestamp 1745462530
transform 1 0 4108 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_1822
timestamp 1745462530
transform 1 0 4068 0 1 2085
box -3 -3 3 3
use M3_M2  M3_M2_1823
timestamp 1745462530
transform 1 0 3940 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_1824
timestamp 1745462530
transform 1 0 4236 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_1825
timestamp 1745462530
transform 1 0 4212 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_1826
timestamp 1745462530
transform 1 0 4212 0 1 2755
box -3 -3 3 3
use M3_M2  M3_M2_1827
timestamp 1745462530
transform 1 0 4148 0 1 2755
box -3 -3 3 3
use M3_M2  M3_M2_1828
timestamp 1745462530
transform 1 0 4116 0 1 2755
box -3 -3 3 3
use M3_M2  M3_M2_1829
timestamp 1745462530
transform 1 0 4244 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_1830
timestamp 1745462530
transform 1 0 4180 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_1831
timestamp 1745462530
transform 1 0 4252 0 1 2435
box -3 -3 3 3
use M3_M2  M3_M2_1832
timestamp 1745462530
transform 1 0 4164 0 1 2435
box -3 -3 3 3
use M3_M2  M3_M2_1833
timestamp 1745462530
transform 1 0 3372 0 1 3465
box -3 -3 3 3
use M3_M2  M3_M2_1834
timestamp 1745462530
transform 1 0 3356 0 1 3465
box -3 -3 3 3
use M3_M2  M3_M2_1835
timestamp 1745462530
transform 1 0 3100 0 1 3465
box -3 -3 3 3
use M3_M2  M3_M2_1836
timestamp 1745462530
transform 1 0 3052 0 1 3465
box -3 -3 3 3
use M3_M2  M3_M2_1837
timestamp 1745462530
transform 1 0 2924 0 1 3525
box -3 -3 3 3
use M3_M2  M3_M2_1838
timestamp 1745462530
transform 1 0 2924 0 1 3465
box -3 -3 3 3
use M3_M2  M3_M2_1839
timestamp 1745462530
transform 1 0 2884 0 1 3525
box -3 -3 3 3
use M3_M2  M3_M2_1840
timestamp 1745462530
transform 1 0 2492 0 1 3535
box -3 -3 3 3
use M3_M2  M3_M2_1841
timestamp 1745462530
transform 1 0 2436 0 1 3535
box -3 -3 3 3
use M3_M2  M3_M2_1842
timestamp 1745462530
transform 1 0 3260 0 1 3545
box -3 -3 3 3
use M3_M2  M3_M2_1843
timestamp 1745462530
transform 1 0 3156 0 1 3535
box -3 -3 3 3
use M3_M2  M3_M2_1844
timestamp 1745462530
transform 1 0 3012 0 1 3605
box -3 -3 3 3
use M3_M2  M3_M2_1845
timestamp 1745462530
transform 1 0 3004 0 1 3545
box -3 -3 3 3
use M3_M2  M3_M2_1846
timestamp 1745462530
transform 1 0 2804 0 1 3625
box -3 -3 3 3
use M3_M2  M3_M2_1847
timestamp 1745462530
transform 1 0 2780 0 1 3605
box -3 -3 3 3
use M3_M2  M3_M2_1848
timestamp 1745462530
transform 1 0 2444 0 1 3605
box -3 -3 3 3
use M3_M2  M3_M2_1849
timestamp 1745462530
transform 1 0 2396 0 1 3365
box -3 -3 3 3
use M3_M2  M3_M2_1850
timestamp 1745462530
transform 1 0 2356 0 1 3365
box -3 -3 3 3
use M3_M2  M3_M2_1851
timestamp 1745462530
transform 1 0 2348 0 1 3605
box -3 -3 3 3
use M3_M2  M3_M2_1852
timestamp 1745462530
transform 1 0 3516 0 1 4145
box -3 -3 3 3
use M3_M2  M3_M2_1853
timestamp 1745462530
transform 1 0 3476 0 1 4145
box -3 -3 3 3
use M3_M2  M3_M2_1854
timestamp 1745462530
transform 1 0 3556 0 1 3405
box -3 -3 3 3
use M3_M2  M3_M2_1855
timestamp 1745462530
transform 1 0 3516 0 1 3495
box -3 -3 3 3
use M3_M2  M3_M2_1856
timestamp 1745462530
transform 1 0 3516 0 1 3405
box -3 -3 3 3
use M3_M2  M3_M2_1857
timestamp 1745462530
transform 1 0 3476 0 1 3495
box -3 -3 3 3
use M3_M2  M3_M2_1858
timestamp 1745462530
transform 1 0 3428 0 1 3495
box -3 -3 3 3
use M3_M2  M3_M2_1859
timestamp 1745462530
transform 1 0 3428 0 1 3425
box -3 -3 3 3
use M3_M2  M3_M2_1860
timestamp 1745462530
transform 1 0 2892 0 1 3425
box -3 -3 3 3
use M3_M2  M3_M2_1861
timestamp 1745462530
transform 1 0 2724 0 1 3425
box -3 -3 3 3
use M3_M2  M3_M2_1862
timestamp 1745462530
transform 1 0 2644 0 1 3425
box -3 -3 3 3
use M3_M2  M3_M2_1863
timestamp 1745462530
transform 1 0 2532 0 1 3425
box -3 -3 3 3
use M3_M2  M3_M2_1864
timestamp 1745462530
transform 1 0 2532 0 1 3405
box -3 -3 3 3
use M3_M2  M3_M2_1865
timestamp 1745462530
transform 1 0 2484 0 1 3405
box -3 -3 3 3
use M3_M2  M3_M2_1866
timestamp 1745462530
transform 1 0 4332 0 1 3745
box -3 -3 3 3
use M3_M2  M3_M2_1867
timestamp 1745462530
transform 1 0 4292 0 1 3745
box -3 -3 3 3
use M3_M2  M3_M2_1868
timestamp 1745462530
transform 1 0 4244 0 1 3745
box -3 -3 3 3
use M3_M2  M3_M2_1869
timestamp 1745462530
transform 1 0 4220 0 1 3745
box -3 -3 3 3
use M3_M2  M3_M2_1870
timestamp 1745462530
transform 1 0 2044 0 1 3915
box -3 -3 3 3
use M3_M2  M3_M2_1871
timestamp 1745462530
transform 1 0 2012 0 1 3915
box -3 -3 3 3
use M3_M2  M3_M2_1872
timestamp 1745462530
transform 1 0 3332 0 1 3145
box -3 -3 3 3
use M3_M2  M3_M2_1873
timestamp 1745462530
transform 1 0 3292 0 1 3145
box -3 -3 3 3
use M3_M2  M3_M2_1874
timestamp 1745462530
transform 1 0 3268 0 1 3085
box -3 -3 3 3
use M3_M2  M3_M2_1875
timestamp 1745462530
transform 1 0 3212 0 1 3085
box -3 -3 3 3
use M3_M2  M3_M2_1876
timestamp 1745462530
transform 1 0 3204 0 1 3205
box -3 -3 3 3
use M3_M2  M3_M2_1877
timestamp 1745462530
transform 1 0 2876 0 1 3205
box -3 -3 3 3
use M3_M2  M3_M2_1878
timestamp 1745462530
transform 1 0 2844 0 1 3255
box -3 -3 3 3
use M3_M2  M3_M2_1879
timestamp 1745462530
transform 1 0 2684 0 1 3255
box -3 -3 3 3
use M3_M2  M3_M2_1880
timestamp 1745462530
transform 1 0 2596 0 1 3255
box -3 -3 3 3
use M3_M2  M3_M2_1881
timestamp 1745462530
transform 1 0 2404 0 1 3245
box -3 -3 3 3
use M3_M2  M3_M2_1882
timestamp 1745462530
transform 1 0 4252 0 1 3185
box -3 -3 3 3
use M3_M2  M3_M2_1883
timestamp 1745462530
transform 1 0 4204 0 1 3185
box -3 -3 3 3
use M3_M2  M3_M2_1884
timestamp 1745462530
transform 1 0 3844 0 1 3735
box -3 -3 3 3
use M3_M2  M3_M2_1885
timestamp 1745462530
transform 1 0 3812 0 1 3735
box -3 -3 3 3
use M3_M2  M3_M2_1886
timestamp 1745462530
transform 1 0 2756 0 1 3015
box -3 -3 3 3
use M3_M2  M3_M2_1887
timestamp 1745462530
transform 1 0 2708 0 1 3015
box -3 -3 3 3
use M3_M2  M3_M2_1888
timestamp 1745462530
transform 1 0 2676 0 1 3025
box -3 -3 3 3
use M3_M2  M3_M2_1889
timestamp 1745462530
transform 1 0 2556 0 1 3025
box -3 -3 3 3
use M3_M2  M3_M2_1890
timestamp 1745462530
transform 1 0 3492 0 1 3305
box -3 -3 3 3
use M3_M2  M3_M2_1891
timestamp 1745462530
transform 1 0 3444 0 1 3305
box -3 -3 3 3
use M3_M2  M3_M2_1892
timestamp 1745462530
transform 1 0 3388 0 1 3305
box -3 -3 3 3
use M3_M2  M3_M2_1893
timestamp 1745462530
transform 1 0 3348 0 1 3305
box -3 -3 3 3
use M3_M2  M3_M2_1894
timestamp 1745462530
transform 1 0 2916 0 1 3305
box -3 -3 3 3
use M3_M2  M3_M2_1895
timestamp 1745462530
transform 1 0 2756 0 1 3335
box -3 -3 3 3
use M3_M2  M3_M2_1896
timestamp 1745462530
transform 1 0 2756 0 1 3305
box -3 -3 3 3
use M3_M2  M3_M2_1897
timestamp 1745462530
transform 1 0 2748 0 1 3175
box -3 -3 3 3
use M3_M2  M3_M2_1898
timestamp 1745462530
transform 1 0 2724 0 1 3335
box -3 -3 3 3
use M3_M2  M3_M2_1899
timestamp 1745462530
transform 1 0 2716 0 1 3175
box -3 -3 3 3
use M3_M2  M3_M2_1900
timestamp 1745462530
transform 1 0 2564 0 1 3335
box -3 -3 3 3
use M3_M2  M3_M2_1901
timestamp 1745462530
transform 1 0 2500 0 1 3335
box -3 -3 3 3
use M3_M2  M3_M2_1902
timestamp 1745462530
transform 1 0 4100 0 1 3545
box -3 -3 3 3
use M3_M2  M3_M2_1903
timestamp 1745462530
transform 1 0 4060 0 1 3545
box -3 -3 3 3
use M3_M2  M3_M2_1904
timestamp 1745462530
transform 1 0 4076 0 1 3585
box -3 -3 3 3
use M3_M2  M3_M2_1905
timestamp 1745462530
transform 1 0 4044 0 1 3585
box -3 -3 3 3
use M3_M2  M3_M2_1906
timestamp 1745462530
transform 1 0 3468 0 1 3095
box -3 -3 3 3
use M3_M2  M3_M2_1907
timestamp 1745462530
transform 1 0 3412 0 1 3185
box -3 -3 3 3
use M3_M2  M3_M2_1908
timestamp 1745462530
transform 1 0 3412 0 1 3095
box -3 -3 3 3
use M3_M2  M3_M2_1909
timestamp 1745462530
transform 1 0 3348 0 1 3185
box -3 -3 3 3
use M3_M2  M3_M2_1910
timestamp 1745462530
transform 1 0 2844 0 1 3185
box -3 -3 3 3
use M3_M2  M3_M2_1911
timestamp 1745462530
transform 1 0 2748 0 1 3185
box -3 -3 3 3
use M3_M2  M3_M2_1912
timestamp 1745462530
transform 1 0 2540 0 1 3185
box -3 -3 3 3
use M3_M2  M3_M2_1913
timestamp 1745462530
transform 1 0 1908 0 1 3955
box -3 -3 3 3
use M3_M2  M3_M2_1914
timestamp 1745462530
transform 1 0 1892 0 1 3955
box -3 -3 3 3
use M3_M2  M3_M2_1915
timestamp 1745462530
transform 1 0 4252 0 1 3345
box -3 -3 3 3
use M3_M2  M3_M2_1916
timestamp 1745462530
transform 1 0 4212 0 1 3345
box -3 -3 3 3
use M3_M2  M3_M2_1917
timestamp 1745462530
transform 1 0 4252 0 1 3395
box -3 -3 3 3
use M3_M2  M3_M2_1918
timestamp 1745462530
transform 1 0 4204 0 1 3395
box -3 -3 3 3
use M3_M2  M3_M2_1919
timestamp 1745462530
transform 1 0 3980 0 1 3225
box -3 -3 3 3
use M3_M2  M3_M2_1920
timestamp 1745462530
transform 1 0 3948 0 1 3225
box -3 -3 3 3
use M3_M2  M3_M2_1921
timestamp 1745462530
transform 1 0 3564 0 1 3535
box -3 -3 3 3
use M3_M2  M3_M2_1922
timestamp 1745462530
transform 1 0 3540 0 1 3535
box -3 -3 3 3
use M3_M2  M3_M2_1923
timestamp 1745462530
transform 1 0 3500 0 1 3535
box -3 -3 3 3
use M3_M2  M3_M2_1924
timestamp 1745462530
transform 1 0 3444 0 1 3555
box -3 -3 3 3
use M3_M2  M3_M2_1925
timestamp 1745462530
transform 1 0 3444 0 1 3535
box -3 -3 3 3
use M3_M2  M3_M2_1926
timestamp 1745462530
transform 1 0 2956 0 1 3555
box -3 -3 3 3
use M3_M2  M3_M2_1927
timestamp 1745462530
transform 1 0 2732 0 1 3545
box -3 -3 3 3
use M3_M2  M3_M2_1928
timestamp 1745462530
transform 1 0 2692 0 1 3545
box -3 -3 3 3
use M3_M2  M3_M2_1929
timestamp 1745462530
transform 1 0 2604 0 1 3545
box -3 -3 3 3
use M3_M2  M3_M2_1930
timestamp 1745462530
transform 1 0 2548 0 1 3545
box -3 -3 3 3
use M3_M2  M3_M2_1931
timestamp 1745462530
transform 1 0 3012 0 1 3975
box -3 -3 3 3
use M3_M2  M3_M2_1932
timestamp 1745462530
transform 1 0 2972 0 1 3975
box -3 -3 3 3
use M3_M2  M3_M2_1933
timestamp 1745462530
transform 1 0 3788 0 1 4035
box -3 -3 3 3
use M3_M2  M3_M2_1934
timestamp 1745462530
transform 1 0 3756 0 1 4035
box -3 -3 3 3
use M3_M2  M3_M2_1935
timestamp 1745462530
transform 1 0 3716 0 1 3965
box -3 -3 3 3
use M3_M2  M3_M2_1936
timestamp 1745462530
transform 1 0 3684 0 1 3965
box -3 -3 3 3
use M3_M2  M3_M2_1937
timestamp 1745462530
transform 1 0 3740 0 1 4105
box -3 -3 3 3
use M3_M2  M3_M2_1938
timestamp 1745462530
transform 1 0 3700 0 1 4105
box -3 -3 3 3
use M3_M2  M3_M2_1939
timestamp 1745462530
transform 1 0 3204 0 1 3365
box -3 -3 3 3
use M3_M2  M3_M2_1940
timestamp 1745462530
transform 1 0 3164 0 1 3365
box -3 -3 3 3
use M3_M2  M3_M2_1941
timestamp 1745462530
transform 1 0 3116 0 1 3365
box -3 -3 3 3
use M3_M2  M3_M2_1942
timestamp 1745462530
transform 1 0 3036 0 1 3365
box -3 -3 3 3
use M3_M2  M3_M2_1943
timestamp 1745462530
transform 1 0 2852 0 1 3365
box -3 -3 3 3
use M3_M2  M3_M2_1944
timestamp 1745462530
transform 1 0 2644 0 1 3365
box -3 -3 3 3
use M3_M2  M3_M2_1945
timestamp 1745462530
transform 1 0 2620 0 1 3365
box -3 -3 3 3
use M3_M2  M3_M2_1946
timestamp 1745462530
transform 1 0 2596 0 1 3365
box -3 -3 3 3
use M3_M2  M3_M2_1947
timestamp 1745462530
transform 1 0 3140 0 1 3865
box -3 -3 3 3
use M3_M2  M3_M2_1948
timestamp 1745462530
transform 1 0 3028 0 1 3865
box -3 -3 3 3
use M3_M2  M3_M2_1949
timestamp 1745462530
transform 1 0 1748 0 1 3815
box -3 -3 3 3
use M3_M2  M3_M2_1950
timestamp 1745462530
transform 1 0 1604 0 1 3815
box -3 -3 3 3
use M3_M2  M3_M2_1951
timestamp 1745462530
transform 1 0 2804 0 1 3945
box -3 -3 3 3
use M3_M2  M3_M2_1952
timestamp 1745462530
transform 1 0 2796 0 1 3725
box -3 -3 3 3
use M3_M2  M3_M2_1953
timestamp 1745462530
transform 1 0 2780 0 1 3725
box -3 -3 3 3
use M3_M2  M3_M2_1954
timestamp 1745462530
transform 1 0 2772 0 1 3945
box -3 -3 3 3
use M3_M2  M3_M2_1955
timestamp 1745462530
transform 1 0 1724 0 1 3715
box -3 -3 3 3
use M3_M2  M3_M2_1956
timestamp 1745462530
transform 1 0 1580 0 1 3715
box -3 -3 3 3
use M3_M2  M3_M2_1957
timestamp 1745462530
transform 1 0 4084 0 1 3315
box -3 -3 3 3
use M3_M2  M3_M2_1958
timestamp 1745462530
transform 1 0 4052 0 1 3315
box -3 -3 3 3
use M3_M2  M3_M2_1959
timestamp 1745462530
transform 1 0 1828 0 1 3955
box -3 -3 3 3
use M3_M2  M3_M2_1960
timestamp 1745462530
transform 1 0 1708 0 1 3955
box -3 -3 3 3
use M3_M2  M3_M2_1961
timestamp 1745462530
transform 1 0 1836 0 1 3795
box -3 -3 3 3
use M3_M2  M3_M2_1962
timestamp 1745462530
transform 1 0 1740 0 1 3795
box -3 -3 3 3
use M3_M2  M3_M2_1963
timestamp 1745462530
transform 1 0 1716 0 1 3905
box -3 -3 3 3
use M3_M2  M3_M2_1964
timestamp 1745462530
transform 1 0 1668 0 1 3905
box -3 -3 3 3
use M3_M2  M3_M2_1965
timestamp 1745462530
transform 1 0 1500 0 1 3905
box -3 -3 3 3
use M3_M2  M3_M2_1966
timestamp 1745462530
transform 1 0 1684 0 1 3855
box -3 -3 3 3
use M3_M2  M3_M2_1967
timestamp 1745462530
transform 1 0 1612 0 1 3855
box -3 -3 3 3
use M3_M2  M3_M2_1968
timestamp 1745462530
transform 1 0 1884 0 1 3915
box -3 -3 3 3
use M3_M2  M3_M2_1969
timestamp 1745462530
transform 1 0 1844 0 1 3915
box -3 -3 3 3
use M3_M2  M3_M2_1970
timestamp 1745462530
transform 1 0 2044 0 1 3865
box -3 -3 3 3
use M3_M2  M3_M2_1971
timestamp 1745462530
transform 1 0 1948 0 1 3865
box -3 -3 3 3
use M3_M2  M3_M2_1972
timestamp 1745462530
transform 1 0 2076 0 1 3695
box -3 -3 3 3
use M3_M2  M3_M2_1973
timestamp 1745462530
transform 1 0 2036 0 1 3695
box -3 -3 3 3
use M3_M2  M3_M2_1974
timestamp 1745462530
transform 1 0 2876 0 1 3785
box -3 -3 3 3
use M3_M2  M3_M2_1975
timestamp 1745462530
transform 1 0 2660 0 1 3785
box -3 -3 3 3
use M3_M2  M3_M2_1976
timestamp 1745462530
transform 1 0 2708 0 1 3865
box -3 -3 3 3
use M3_M2  M3_M2_1977
timestamp 1745462530
transform 1 0 2692 0 1 3865
box -3 -3 3 3
use M3_M2  M3_M2_1978
timestamp 1745462530
transform 1 0 2692 0 1 3815
box -3 -3 3 3
use M3_M2  M3_M2_1979
timestamp 1745462530
transform 1 0 2564 0 1 3815
box -3 -3 3 3
use M3_M2  M3_M2_1980
timestamp 1745462530
transform 1 0 2068 0 1 3795
box -3 -3 3 3
use M3_M2  M3_M2_1981
timestamp 1745462530
transform 1 0 2020 0 1 3795
box -3 -3 3 3
use M3_M2  M3_M2_1982
timestamp 1745462530
transform 1 0 2044 0 1 3755
box -3 -3 3 3
use M3_M2  M3_M2_1983
timestamp 1745462530
transform 1 0 2004 0 1 3755
box -3 -3 3 3
use M3_M2  M3_M2_1984
timestamp 1745462530
transform 1 0 3980 0 1 3585
box -3 -3 3 3
use M3_M2  M3_M2_1985
timestamp 1745462530
transform 1 0 3916 0 1 3585
box -3 -3 3 3
use M3_M2  M3_M2_1986
timestamp 1745462530
transform 1 0 2940 0 1 3885
box -3 -3 3 3
use M3_M2  M3_M2_1987
timestamp 1745462530
transform 1 0 2900 0 1 3885
box -3 -3 3 3
use M3_M2  M3_M2_1988
timestamp 1745462530
transform 1 0 2900 0 1 3755
box -3 -3 3 3
use M3_M2  M3_M2_1989
timestamp 1745462530
transform 1 0 2628 0 1 3755
box -3 -3 3 3
use M3_M2  M3_M2_1990
timestamp 1745462530
transform 1 0 2612 0 1 3945
box -3 -3 3 3
use M3_M2  M3_M2_1991
timestamp 1745462530
transform 1 0 2556 0 1 3945
box -3 -3 3 3
use M3_M2  M3_M2_1992
timestamp 1745462530
transform 1 0 2524 0 1 3945
box -3 -3 3 3
use M3_M2  M3_M2_1993
timestamp 1745462530
transform 1 0 2308 0 1 4095
box -3 -3 3 3
use M3_M2  M3_M2_1994
timestamp 1745462530
transform 1 0 2276 0 1 4095
box -3 -3 3 3
use M3_M2  M3_M2_1995
timestamp 1745462530
transform 1 0 2508 0 1 4145
box -3 -3 3 3
use M3_M2  M3_M2_1996
timestamp 1745462530
transform 1 0 2460 0 1 4145
box -3 -3 3 3
use M3_M2  M3_M2_1997
timestamp 1745462530
transform 1 0 2364 0 1 4145
box -3 -3 3 3
use M3_M2  M3_M2_1998
timestamp 1745462530
transform 1 0 3732 0 1 4115
box -3 -3 3 3
use M3_M2  M3_M2_1999
timestamp 1745462530
transform 1 0 3452 0 1 4115
box -3 -3 3 3
use M3_M2  M3_M2_2000
timestamp 1745462530
transform 1 0 3724 0 1 3955
box -3 -3 3 3
use M3_M2  M3_M2_2001
timestamp 1745462530
transform 1 0 3588 0 1 3955
box -3 -3 3 3
use M3_M2  M3_M2_2002
timestamp 1745462530
transform 1 0 3908 0 1 4145
box -3 -3 3 3
use M3_M2  M3_M2_2003
timestamp 1745462530
transform 1 0 3876 0 1 4145
box -3 -3 3 3
use M3_M2  M3_M2_2004
timestamp 1745462530
transform 1 0 3556 0 1 4145
box -3 -3 3 3
use M3_M2  M3_M2_2005
timestamp 1745462530
transform 1 0 3772 0 1 4015
box -3 -3 3 3
use M3_M2  M3_M2_2006
timestamp 1745462530
transform 1 0 3572 0 1 4015
box -3 -3 3 3
use M3_M2  M3_M2_2007
timestamp 1745462530
transform 1 0 3068 0 1 4045
box -3 -3 3 3
use M3_M2  M3_M2_2008
timestamp 1745462530
transform 1 0 3004 0 1 4045
box -3 -3 3 3
use M3_M2  M3_M2_2009
timestamp 1745462530
transform 1 0 2228 0 1 4145
box -3 -3 3 3
use M3_M2  M3_M2_2010
timestamp 1745462530
transform 1 0 2204 0 1 4145
box -3 -3 3 3
use M3_M2  M3_M2_2011
timestamp 1745462530
transform 1 0 2196 0 1 4105
box -3 -3 3 3
use M3_M2  M3_M2_2012
timestamp 1745462530
transform 1 0 2172 0 1 4105
box -3 -3 3 3
use M3_M2  M3_M2_2013
timestamp 1745462530
transform 1 0 2428 0 1 4195
box -3 -3 3 3
use M3_M2  M3_M2_2014
timestamp 1745462530
transform 1 0 2388 0 1 4195
box -3 -3 3 3
use M3_M2  M3_M2_2015
timestamp 1745462530
transform 1 0 2348 0 1 4195
box -3 -3 3 3
use M3_M2  M3_M2_2016
timestamp 1745462530
transform 1 0 3420 0 1 4115
box -3 -3 3 3
use M3_M2  M3_M2_2017
timestamp 1745462530
transform 1 0 3308 0 1 4115
box -3 -3 3 3
use M3_M2  M3_M2_2018
timestamp 1745462530
transform 1 0 3204 0 1 4115
box -3 -3 3 3
use M3_M2  M3_M2_2019
timestamp 1745462530
transform 1 0 3596 0 1 4005
box -3 -3 3 3
use M3_M2  M3_M2_2020
timestamp 1745462530
transform 1 0 3524 0 1 4005
box -3 -3 3 3
use M3_M2  M3_M2_2021
timestamp 1745462530
transform 1 0 3532 0 1 4125
box -3 -3 3 3
use M3_M2  M3_M2_2022
timestamp 1745462530
transform 1 0 3508 0 1 4215
box -3 -3 3 3
use M3_M2  M3_M2_2023
timestamp 1745462530
transform 1 0 3428 0 1 4215
box -3 -3 3 3
use M3_M2  M3_M2_2024
timestamp 1745462530
transform 1 0 3428 0 1 4125
box -3 -3 3 3
use M3_M2  M3_M2_2025
timestamp 1745462530
transform 1 0 3396 0 1 4125
box -3 -3 3 3
use M3_M2  M3_M2_2026
timestamp 1745462530
transform 1 0 3564 0 1 4105
box -3 -3 3 3
use M3_M2  M3_M2_2027
timestamp 1745462530
transform 1 0 3508 0 1 4105
box -3 -3 3 3
use M3_M2  M3_M2_2028
timestamp 1745462530
transform 1 0 3084 0 1 4195
box -3 -3 3 3
use M3_M2  M3_M2_2029
timestamp 1745462530
transform 1 0 3044 0 1 4195
box -3 -3 3 3
use M3_M2  M3_M2_2030
timestamp 1745462530
transform 1 0 2780 0 1 4105
box -3 -3 3 3
use M3_M2  M3_M2_2031
timestamp 1745462530
transform 1 0 2764 0 1 4105
box -3 -3 3 3
use M3_M2  M3_M2_2032
timestamp 1745462530
transform 1 0 2660 0 1 4105
box -3 -3 3 3
use M3_M2  M3_M2_2033
timestamp 1745462530
transform 1 0 2396 0 1 4005
box -3 -3 3 3
use M3_M2  M3_M2_2034
timestamp 1745462530
transform 1 0 2348 0 1 4005
box -3 -3 3 3
use M3_M2  M3_M2_2035
timestamp 1745462530
transform 1 0 3684 0 1 3815
box -3 -3 3 3
use M3_M2  M3_M2_2036
timestamp 1745462530
transform 1 0 3684 0 1 3775
box -3 -3 3 3
use M3_M2  M3_M2_2037
timestamp 1745462530
transform 1 0 3612 0 1 3775
box -3 -3 3 3
use M3_M2  M3_M2_2038
timestamp 1745462530
transform 1 0 3564 0 1 3815
box -3 -3 3 3
use M3_M2  M3_M2_2039
timestamp 1745462530
transform 1 0 3620 0 1 3935
box -3 -3 3 3
use M3_M2  M3_M2_2040
timestamp 1745462530
transform 1 0 3476 0 1 3935
box -3 -3 3 3
use M3_M2  M3_M2_2041
timestamp 1745462530
transform 1 0 3652 0 1 3785
box -3 -3 3 3
use M3_M2  M3_M2_2042
timestamp 1745462530
transform 1 0 3508 0 1 3785
box -3 -3 3 3
use M3_M2  M3_M2_2043
timestamp 1745462530
transform 1 0 3108 0 1 3935
box -3 -3 3 3
use M3_M2  M3_M2_2044
timestamp 1745462530
transform 1 0 3092 0 1 3935
box -3 -3 3 3
use M3_M2  M3_M2_2045
timestamp 1745462530
transform 1 0 2860 0 1 3935
box -3 -3 3 3
use M3_M2  M3_M2_2046
timestamp 1745462530
transform 1 0 2796 0 1 3935
box -3 -3 3 3
use M3_M2  M3_M2_2047
timestamp 1745462530
transform 1 0 2788 0 1 3955
box -3 -3 3 3
use M3_M2  M3_M2_2048
timestamp 1745462530
transform 1 0 2708 0 1 3955
box -3 -3 3 3
use M3_M2  M3_M2_2049
timestamp 1745462530
transform 1 0 2124 0 1 3985
box -3 -3 3 3
use M3_M2  M3_M2_2050
timestamp 1745462530
transform 1 0 2100 0 1 3985
box -3 -3 3 3
use M3_M2  M3_M2_2051
timestamp 1745462530
transform 1 0 2404 0 1 3895
box -3 -3 3 3
use M3_M2  M3_M2_2052
timestamp 1745462530
transform 1 0 2372 0 1 3895
box -3 -3 3 3
use M3_M2  M3_M2_2053
timestamp 1745462530
transform 1 0 2332 0 1 3895
box -3 -3 3 3
use M3_M2  M3_M2_2054
timestamp 1745462530
transform 1 0 3228 0 1 3935
box -3 -3 3 3
use M3_M2  M3_M2_2055
timestamp 1745462530
transform 1 0 3180 0 1 3935
box -3 -3 3 3
use M3_M2  M3_M2_2056
timestamp 1745462530
transform 1 0 3516 0 1 3815
box -3 -3 3 3
use M3_M2  M3_M2_2057
timestamp 1745462530
transform 1 0 3396 0 1 3815
box -3 -3 3 3
use M3_M2  M3_M2_2058
timestamp 1745462530
transform 1 0 3468 0 1 3915
box -3 -3 3 3
use M3_M2  M3_M2_2059
timestamp 1745462530
transform 1 0 3316 0 1 3915
box -3 -3 3 3
use M3_M2  M3_M2_2060
timestamp 1745462530
transform 1 0 3484 0 1 3865
box -3 -3 3 3
use M3_M2  M3_M2_2061
timestamp 1745462530
transform 1 0 3420 0 1 3865
box -3 -3 3 3
use M3_M2  M3_M2_2062
timestamp 1745462530
transform 1 0 2268 0 1 3825
box -3 -3 3 3
use M3_M2  M3_M2_2063
timestamp 1745462530
transform 1 0 2236 0 1 3825
box -3 -3 3 3
use M3_M2  M3_M2_2064
timestamp 1745462530
transform 1 0 2180 0 1 3825
box -3 -3 3 3
use M3_M2  M3_M2_2065
timestamp 1745462530
transform 1 0 2140 0 1 3825
box -3 -3 3 3
use M3_M2  M3_M2_2066
timestamp 1745462530
transform 1 0 484 0 1 4015
box -3 -3 3 3
use M3_M2  M3_M2_2067
timestamp 1745462530
transform 1 0 420 0 1 4025
box -3 -3 3 3
use M3_M2  M3_M2_2068
timestamp 1745462530
transform 1 0 340 0 1 4025
box -3 -3 3 3
use M3_M2  M3_M2_2069
timestamp 1745462530
transform 1 0 452 0 1 4035
box -3 -3 3 3
use M3_M2  M3_M2_2070
timestamp 1745462530
transform 1 0 316 0 1 4035
box -3 -3 3 3
use M3_M2  M3_M2_2071
timestamp 1745462530
transform 1 0 1284 0 1 3825
box -3 -3 3 3
use M3_M2  M3_M2_2072
timestamp 1745462530
transform 1 0 1228 0 1 3835
box -3 -3 3 3
use M3_M2  M3_M2_2073
timestamp 1745462530
transform 1 0 468 0 1 3835
box -3 -3 3 3
use M3_M2  M3_M2_2074
timestamp 1745462530
transform 1 0 468 0 1 3795
box -3 -3 3 3
use M3_M2  M3_M2_2075
timestamp 1745462530
transform 1 0 204 0 1 3795
box -3 -3 3 3
use M3_M2  M3_M2_2076
timestamp 1745462530
transform 1 0 1580 0 1 3465
box -3 -3 3 3
use M3_M2  M3_M2_2077
timestamp 1745462530
transform 1 0 1540 0 1 3465
box -3 -3 3 3
use M3_M2  M3_M2_2078
timestamp 1745462530
transform 1 0 1556 0 1 3515
box -3 -3 3 3
use M3_M2  M3_M2_2079
timestamp 1745462530
transform 1 0 1508 0 1 3515
box -3 -3 3 3
use M3_M2  M3_M2_2080
timestamp 1745462530
transform 1 0 1444 0 1 3635
box -3 -3 3 3
use M3_M2  M3_M2_2081
timestamp 1745462530
transform 1 0 1340 0 1 3635
box -3 -3 3 3
use M3_M2  M3_M2_2082
timestamp 1745462530
transform 1 0 1460 0 1 3405
box -3 -3 3 3
use M3_M2  M3_M2_2083
timestamp 1745462530
transform 1 0 1444 0 1 3405
box -3 -3 3 3
use M3_M2  M3_M2_2084
timestamp 1745462530
transform 1 0 1012 0 1 4125
box -3 -3 3 3
use M3_M2  M3_M2_2085
timestamp 1745462530
transform 1 0 932 0 1 4125
box -3 -3 3 3
use M3_M2  M3_M2_2086
timestamp 1745462530
transform 1 0 3884 0 1 4195
box -3 -3 3 3
use M3_M2  M3_M2_2087
timestamp 1745462530
transform 1 0 3836 0 1 4195
box -3 -3 3 3
use M3_M2  M3_M2_2088
timestamp 1745462530
transform 1 0 3804 0 1 4195
box -3 -3 3 3
use M3_M2  M3_M2_2089
timestamp 1745462530
transform 1 0 3668 0 1 4195
box -3 -3 3 3
use M3_M2  M3_M2_2090
timestamp 1745462530
transform 1 0 3612 0 1 4195
box -3 -3 3 3
use M3_M2  M3_M2_2091
timestamp 1745462530
transform 1 0 3524 0 1 4195
box -3 -3 3 3
use M3_M2  M3_M2_2092
timestamp 1745462530
transform 1 0 3516 0 1 4165
box -3 -3 3 3
use M3_M2  M3_M2_2093
timestamp 1745462530
transform 1 0 3348 0 1 4085
box -3 -3 3 3
use M3_M2  M3_M2_2094
timestamp 1745462530
transform 1 0 3300 0 1 4165
box -3 -3 3 3
use M3_M2  M3_M2_2095
timestamp 1745462530
transform 1 0 3300 0 1 4085
box -3 -3 3 3
use M3_M2  M3_M2_2096
timestamp 1745462530
transform 1 0 3060 0 1 4165
box -3 -3 3 3
use M3_M2  M3_M2_2097
timestamp 1745462530
transform 1 0 3020 0 1 4165
box -3 -3 3 3
use M3_M2  M3_M2_2098
timestamp 1745462530
transform 1 0 2836 0 1 4165
box -3 -3 3 3
use M3_M2  M3_M2_2099
timestamp 1745462530
transform 1 0 2700 0 1 4165
box -3 -3 3 3
use M3_M2  M3_M2_2100
timestamp 1745462530
transform 1 0 2324 0 1 4165
box -3 -3 3 3
use M3_M2  M3_M2_2101
timestamp 1745462530
transform 1 0 2284 0 1 4275
box -3 -3 3 3
use M3_M2  M3_M2_2102
timestamp 1745462530
transform 1 0 2196 0 1 4275
box -3 -3 3 3
use M3_M2  M3_M2_2103
timestamp 1745462530
transform 1 0 2132 0 1 4095
box -3 -3 3 3
use M3_M2  M3_M2_2104
timestamp 1745462530
transform 1 0 2044 0 1 4095
box -3 -3 3 3
use M3_M2  M3_M2_2105
timestamp 1745462530
transform 1 0 1540 0 1 4105
box -3 -3 3 3
use M3_M2  M3_M2_2106
timestamp 1745462530
transform 1 0 3860 0 1 4255
box -3 -3 3 3
use M3_M2  M3_M2_2107
timestamp 1745462530
transform 1 0 3828 0 1 4255
box -3 -3 3 3
use M3_M2  M3_M2_2108
timestamp 1745462530
transform 1 0 3820 0 1 4065
box -3 -3 3 3
use M3_M2  M3_M2_2109
timestamp 1745462530
transform 1 0 3780 0 1 4065
box -3 -3 3 3
use M3_M2  M3_M2_2110
timestamp 1745462530
transform 1 0 3652 0 1 4065
box -3 -3 3 3
use M3_M2  M3_M2_2111
timestamp 1745462530
transform 1 0 3580 0 1 4065
box -3 -3 3 3
use M3_M2  M3_M2_2112
timestamp 1745462530
transform 1 0 3500 0 1 4255
box -3 -3 3 3
use M3_M2  M3_M2_2113
timestamp 1745462530
transform 1 0 3332 0 1 4305
box -3 -3 3 3
use M3_M2  M3_M2_2114
timestamp 1745462530
transform 1 0 3332 0 1 4255
box -3 -3 3 3
use M3_M2  M3_M2_2115
timestamp 1745462530
transform 1 0 3332 0 1 4065
box -3 -3 3 3
use M3_M2  M3_M2_2116
timestamp 1745462530
transform 1 0 3044 0 1 4305
box -3 -3 3 3
use M3_M2  M3_M2_2117
timestamp 1745462530
transform 1 0 3004 0 1 4305
box -3 -3 3 3
use M3_M2  M3_M2_2118
timestamp 1745462530
transform 1 0 2820 0 1 4295
box -3 -3 3 3
use M3_M2  M3_M2_2119
timestamp 1745462530
transform 1 0 2820 0 1 4275
box -3 -3 3 3
use M3_M2  M3_M2_2120
timestamp 1745462530
transform 1 0 2684 0 1 4275
box -3 -3 3 3
use M3_M2  M3_M2_2121
timestamp 1745462530
transform 1 0 2660 0 1 4275
box -3 -3 3 3
use M3_M2  M3_M2_2122
timestamp 1745462530
transform 1 0 2644 0 1 4185
box -3 -3 3 3
use M3_M2  M3_M2_2123
timestamp 1745462530
transform 1 0 2308 0 1 4185
box -3 -3 3 3
use M3_M2  M3_M2_2124
timestamp 1745462530
transform 1 0 2172 0 1 4185
box -3 -3 3 3
use M3_M2  M3_M2_2125
timestamp 1745462530
transform 1 0 2132 0 1 4185
box -3 -3 3 3
use M3_M2  M3_M2_2126
timestamp 1745462530
transform 1 0 2028 0 1 4185
box -3 -3 3 3
use M3_M2  M3_M2_2127
timestamp 1745462530
transform 1 0 2028 0 1 4065
box -3 -3 3 3
use M3_M2  M3_M2_2128
timestamp 1745462530
transform 1 0 1764 0 1 4065
box -3 -3 3 3
use M3_M2  M3_M2_2129
timestamp 1745462530
transform 1 0 1764 0 1 4025
box -3 -3 3 3
use M3_M2  M3_M2_2130
timestamp 1745462530
transform 1 0 1388 0 1 4085
box -3 -3 3 3
use M3_M2  M3_M2_2131
timestamp 1745462530
transform 1 0 1388 0 1 4025
box -3 -3 3 3
use M3_M2  M3_M2_2132
timestamp 1745462530
transform 1 0 1356 0 1 4085
box -3 -3 3 3
use M3_M2  M3_M2_2133
timestamp 1745462530
transform 1 0 1108 0 1 4025
box -3 -3 3 3
use M3_M2  M3_M2_2134
timestamp 1745462530
transform 1 0 1044 0 1 4025
box -3 -3 3 3
use M3_M2  M3_M2_2135
timestamp 1745462530
transform 1 0 980 0 1 4025
box -3 -3 3 3
use M3_M2  M3_M2_2136
timestamp 1745462530
transform 1 0 4148 0 1 3915
box -3 -3 3 3
use M3_M2  M3_M2_2137
timestamp 1745462530
transform 1 0 4140 0 1 4045
box -3 -3 3 3
use M3_M2  M3_M2_2138
timestamp 1745462530
transform 1 0 4124 0 1 4255
box -3 -3 3 3
use M3_M2  M3_M2_2139
timestamp 1745462530
transform 1 0 4124 0 1 4045
box -3 -3 3 3
use M3_M2  M3_M2_2140
timestamp 1745462530
transform 1 0 4116 0 1 3915
box -3 -3 3 3
use M3_M2  M3_M2_2141
timestamp 1745462530
transform 1 0 4092 0 1 3915
box -3 -3 3 3
use M3_M2  M3_M2_2142
timestamp 1745462530
transform 1 0 4020 0 1 4045
box -3 -3 3 3
use M3_M2  M3_M2_2143
timestamp 1745462530
transform 1 0 3956 0 1 4325
box -3 -3 3 3
use M3_M2  M3_M2_2144
timestamp 1745462530
transform 1 0 3956 0 1 4255
box -3 -3 3 3
use M3_M2  M3_M2_2145
timestamp 1745462530
transform 1 0 3940 0 1 4045
box -3 -3 3 3
use M3_M2  M3_M2_2146
timestamp 1745462530
transform 1 0 2956 0 1 4325
box -3 -3 3 3
use M3_M2  M3_M2_2147
timestamp 1745462530
transform 1 0 2932 0 1 4325
box -3 -3 3 3
use M3_M2  M3_M2_2148
timestamp 1745462530
transform 1 0 2932 0 1 4235
box -3 -3 3 3
use M3_M2  M3_M2_2149
timestamp 1745462530
transform 1 0 2636 0 1 4235
box -3 -3 3 3
use M3_M2  M3_M2_2150
timestamp 1745462530
transform 1 0 2580 0 1 4235
box -3 -3 3 3
use M3_M2  M3_M2_2151
timestamp 1745462530
transform 1 0 1988 0 1 4245
box -3 -3 3 3
use M3_M2  M3_M2_2152
timestamp 1745462530
transform 1 0 1988 0 1 4175
box -3 -3 3 3
use M3_M2  M3_M2_2153
timestamp 1745462530
transform 1 0 1964 0 1 4175
box -3 -3 3 3
use M3_M2  M3_M2_2154
timestamp 1745462530
transform 1 0 1916 0 1 4175
box -3 -3 3 3
use M3_M2  M3_M2_2155
timestamp 1745462530
transform 1 0 1876 0 1 4175
box -3 -3 3 3
use M3_M2  M3_M2_2156
timestamp 1745462530
transform 1 0 1412 0 1 4175
box -3 -3 3 3
use M3_M2  M3_M2_2157
timestamp 1745462530
transform 1 0 708 0 1 4115
box -3 -3 3 3
use M3_M2  M3_M2_2158
timestamp 1745462530
transform 1 0 644 0 1 4115
box -3 -3 3 3
use M3_M2  M3_M2_2159
timestamp 1745462530
transform 1 0 620 0 1 4195
box -3 -3 3 3
use M3_M2  M3_M2_2160
timestamp 1745462530
transform 1 0 580 0 1 4195
box -3 -3 3 3
use M3_M2  M3_M2_2161
timestamp 1745462530
transform 1 0 204 0 1 4225
box -3 -3 3 3
use M3_M2  M3_M2_2162
timestamp 1745462530
transform 1 0 180 0 1 4225
box -3 -3 3 3
use M3_M2  M3_M2_2163
timestamp 1745462530
transform 1 0 124 0 1 4225
box -3 -3 3 3
use M3_M2  M3_M2_2164
timestamp 1745462530
transform 1 0 132 0 1 3805
box -3 -3 3 3
use M3_M2  M3_M2_2165
timestamp 1745462530
transform 1 0 100 0 1 3805
box -3 -3 3 3
use M3_M2  M3_M2_2166
timestamp 1745462530
transform 1 0 180 0 1 3875
box -3 -3 3 3
use M3_M2  M3_M2_2167
timestamp 1745462530
transform 1 0 132 0 1 3875
box -3 -3 3 3
use M3_M2  M3_M2_2168
timestamp 1745462530
transform 1 0 116 0 1 3875
box -3 -3 3 3
use M3_M2  M3_M2_2169
timestamp 1745462530
transform 1 0 836 0 1 3965
box -3 -3 3 3
use M3_M2  M3_M2_2170
timestamp 1745462530
transform 1 0 780 0 1 3965
box -3 -3 3 3
use M3_M2  M3_M2_2171
timestamp 1745462530
transform 1 0 700 0 1 3965
box -3 -3 3 3
use M3_M2  M3_M2_2172
timestamp 1745462530
transform 1 0 396 0 1 3965
box -3 -3 3 3
use M3_M2  M3_M2_2173
timestamp 1745462530
transform 1 0 308 0 1 3965
box -3 -3 3 3
use M3_M2  M3_M2_2174
timestamp 1745462530
transform 1 0 228 0 1 3965
box -3 -3 3 3
use M3_M2  M3_M2_2175
timestamp 1745462530
transform 1 0 668 0 1 4135
box -3 -3 3 3
use M3_M2  M3_M2_2176
timestamp 1745462530
transform 1 0 652 0 1 4135
box -3 -3 3 3
use M3_M2  M3_M2_2177
timestamp 1745462530
transform 1 0 964 0 1 4145
box -3 -3 3 3
use M3_M2  M3_M2_2178
timestamp 1745462530
transform 1 0 892 0 1 4145
box -3 -3 3 3
use M3_M2  M3_M2_2179
timestamp 1745462530
transform 1 0 1004 0 1 4105
box -3 -3 3 3
use M3_M2  M3_M2_2180
timestamp 1745462530
transform 1 0 932 0 1 4105
box -3 -3 3 3
use M3_M2  M3_M2_2181
timestamp 1745462530
transform 1 0 820 0 1 4105
box -3 -3 3 3
use M3_M2  M3_M2_2182
timestamp 1745462530
transform 1 0 724 0 1 4105
box -3 -3 3 3
use M3_M2  M3_M2_2183
timestamp 1745462530
transform 1 0 1276 0 1 3515
box -3 -3 3 3
use M3_M2  M3_M2_2184
timestamp 1745462530
transform 1 0 1196 0 1 3745
box -3 -3 3 3
use M3_M2  M3_M2_2185
timestamp 1745462530
transform 1 0 1196 0 1 3535
box -3 -3 3 3
use M3_M2  M3_M2_2186
timestamp 1745462530
transform 1 0 1180 0 1 3525
box -3 -3 3 3
use M3_M2  M3_M2_2187
timestamp 1745462530
transform 1 0 1164 0 1 3745
box -3 -3 3 3
use M3_M2  M3_M2_2188
timestamp 1745462530
transform 1 0 956 0 1 4215
box -3 -3 3 3
use M3_M2  M3_M2_2189
timestamp 1745462530
transform 1 0 924 0 1 4215
box -3 -3 3 3
use M3_M2  M3_M2_2190
timestamp 1745462530
transform 1 0 828 0 1 4215
box -3 -3 3 3
use M3_M2  M3_M2_2191
timestamp 1745462530
transform 1 0 828 0 1 4145
box -3 -3 3 3
use M3_M2  M3_M2_2192
timestamp 1745462530
transform 1 0 708 0 1 3745
box -3 -3 3 3
use M3_M2  M3_M2_2193
timestamp 1745462530
transform 1 0 700 0 1 3815
box -3 -3 3 3
use M3_M2  M3_M2_2194
timestamp 1745462530
transform 1 0 524 0 1 3815
box -3 -3 3 3
use M3_M2  M3_M2_2195
timestamp 1745462530
transform 1 0 500 0 1 4145
box -3 -3 3 3
use M3_M2  M3_M2_2196
timestamp 1745462530
transform 1 0 364 0 1 4145
box -3 -3 3 3
use M3_M2  M3_M2_2197
timestamp 1745462530
transform 1 0 260 0 1 3875
box -3 -3 3 3
use M3_M2  M3_M2_2198
timestamp 1745462530
transform 1 0 260 0 1 3815
box -3 -3 3 3
use M3_M2  M3_M2_2199
timestamp 1745462530
transform 1 0 236 0 1 4145
box -3 -3 3 3
use M3_M2  M3_M2_2200
timestamp 1745462530
transform 1 0 236 0 1 3875
box -3 -3 3 3
use M3_M2  M3_M2_2201
timestamp 1745462530
transform 1 0 204 0 1 3875
box -3 -3 3 3
use M3_M2  M3_M2_2202
timestamp 1745462530
transform 1 0 1212 0 1 3465
box -3 -3 3 3
use M3_M2  M3_M2_2203
timestamp 1745462530
transform 1 0 1212 0 1 3385
box -3 -3 3 3
use M3_M2  M3_M2_2204
timestamp 1745462530
transform 1 0 1188 0 1 3465
box -3 -3 3 3
use M3_M2  M3_M2_2205
timestamp 1745462530
transform 1 0 1172 0 1 3385
box -3 -3 3 3
use M3_M2  M3_M2_2206
timestamp 1745462530
transform 1 0 1164 0 1 3725
box -3 -3 3 3
use M3_M2  M3_M2_2207
timestamp 1745462530
transform 1 0 852 0 1 3725
box -3 -3 3 3
use M3_M2  M3_M2_2208
timestamp 1745462530
transform 1 0 740 0 1 3725
box -3 -3 3 3
use M3_M2  M3_M2_2209
timestamp 1745462530
transform 1 0 700 0 1 3585
box -3 -3 3 3
use M3_M2  M3_M2_2210
timestamp 1745462530
transform 1 0 636 0 1 3585
box -3 -3 3 3
use M3_M2  M3_M2_2211
timestamp 1745462530
transform 1 0 604 0 1 3395
box -3 -3 3 3
use M3_M2  M3_M2_2212
timestamp 1745462530
transform 1 0 580 0 1 3585
box -3 -3 3 3
use M3_M2  M3_M2_2213
timestamp 1745462530
transform 1 0 516 0 1 3585
box -3 -3 3 3
use M3_M2  M3_M2_2214
timestamp 1745462530
transform 1 0 500 0 1 3395
box -3 -3 3 3
use M3_M2  M3_M2_2215
timestamp 1745462530
transform 1 0 452 0 1 3585
box -3 -3 3 3
use M3_M2  M3_M2_2216
timestamp 1745462530
transform 1 0 380 0 1 3395
box -3 -3 3 3
use M3_M2  M3_M2_2217
timestamp 1745462530
transform 1 0 1004 0 1 3105
box -3 -3 3 3
use M3_M2  M3_M2_2218
timestamp 1745462530
transform 1 0 972 0 1 3105
box -3 -3 3 3
use M3_M2  M3_M2_2219
timestamp 1745462530
transform 1 0 2164 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_2220
timestamp 1745462530
transform 1 0 908 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_2221
timestamp 1745462530
transform 1 0 2252 0 1 1865
box -3 -3 3 3
use M3_M2  M3_M2_2222
timestamp 1745462530
transform 1 0 2124 0 1 1855
box -3 -3 3 3
use M3_M2  M3_M2_2223
timestamp 1745462530
transform 1 0 2084 0 1 1855
box -3 -3 3 3
use M3_M2  M3_M2_2224
timestamp 1745462530
transform 1 0 1892 0 1 1855
box -3 -3 3 3
use M3_M2  M3_M2_2225
timestamp 1745462530
transform 1 0 1892 0 1 1835
box -3 -3 3 3
use M3_M2  M3_M2_2226
timestamp 1745462530
transform 1 0 1612 0 1 1835
box -3 -3 3 3
use M3_M2  M3_M2_2227
timestamp 1745462530
transform 1 0 2556 0 1 1465
box -3 -3 3 3
use M3_M2  M3_M2_2228
timestamp 1745462530
transform 1 0 2220 0 1 1465
box -3 -3 3 3
use M3_M2  M3_M2_2229
timestamp 1745462530
transform 1 0 2012 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_2230
timestamp 1745462530
transform 1 0 1980 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_2231
timestamp 1745462530
transform 1 0 1980 0 1 1535
box -3 -3 3 3
use M3_M2  M3_M2_2232
timestamp 1745462530
transform 1 0 1948 0 1 1535
box -3 -3 3 3
use M3_M2  M3_M2_2233
timestamp 1745462530
transform 1 0 2276 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_2234
timestamp 1745462530
transform 1 0 2244 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_2235
timestamp 1745462530
transform 1 0 2244 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_2236
timestamp 1745462530
transform 1 0 2004 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_2237
timestamp 1745462530
transform 1 0 1956 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_2238
timestamp 1745462530
transform 1 0 2204 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_2239
timestamp 1745462530
transform 1 0 2132 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_2240
timestamp 1745462530
transform 1 0 2124 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_2241
timestamp 1745462530
transform 1 0 2100 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_2242
timestamp 1745462530
transform 1 0 1572 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_2243
timestamp 1745462530
transform 1 0 1980 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_2244
timestamp 1745462530
transform 1 0 1436 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_2245
timestamp 1745462530
transform 1 0 1332 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_2246
timestamp 1745462530
transform 1 0 2268 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_2247
timestamp 1745462530
transform 1 0 2196 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_2248
timestamp 1745462530
transform 1 0 2164 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_2249
timestamp 1745462530
transform 1 0 2124 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_2250
timestamp 1745462530
transform 1 0 2124 0 1 1295
box -3 -3 3 3
use M3_M2  M3_M2_2251
timestamp 1745462530
transform 1 0 1804 0 1 1295
box -3 -3 3 3
use M3_M2  M3_M2_2252
timestamp 1745462530
transform 1 0 1636 0 1 3925
box -3 -3 3 3
use M3_M2  M3_M2_2253
timestamp 1745462530
transform 1 0 1340 0 1 3925
box -3 -3 3 3
use M3_M2  M3_M2_2254
timestamp 1745462530
transform 1 0 4284 0 1 4195
box -3 -3 3 3
use M3_M2  M3_M2_2255
timestamp 1745462530
transform 1 0 4284 0 1 4055
box -3 -3 3 3
use M3_M2  M3_M2_2256
timestamp 1745462530
transform 1 0 4180 0 1 4195
box -3 -3 3 3
use M3_M2  M3_M2_2257
timestamp 1745462530
transform 1 0 1652 0 1 4195
box -3 -3 3 3
use M3_M2  M3_M2_2258
timestamp 1745462530
transform 1 0 1652 0 1 4055
box -3 -3 3 3
use M3_M2  M3_M2_2259
timestamp 1745462530
transform 1 0 1556 0 1 4195
box -3 -3 3 3
use M3_M2  M3_M2_2260
timestamp 1745462530
transform 1 0 1404 0 1 4215
box -3 -3 3 3
use M3_M2  M3_M2_2261
timestamp 1745462530
transform 1 0 1364 0 1 3985
box -3 -3 3 3
use M3_M2  M3_M2_2262
timestamp 1745462530
transform 1 0 1308 0 1 4215
box -3 -3 3 3
use M3_M2  M3_M2_2263
timestamp 1745462530
transform 1 0 1260 0 1 4215
box -3 -3 3 3
use M3_M2  M3_M2_2264
timestamp 1745462530
transform 1 0 1220 0 1 3985
box -3 -3 3 3
use M3_M2  M3_M2_2265
timestamp 1745462530
transform 1 0 1212 0 1 4215
box -3 -3 3 3
use M3_M2  M3_M2_2266
timestamp 1745462530
transform 1 0 1116 0 1 4215
box -3 -3 3 3
use M3_M2  M3_M2_2267
timestamp 1745462530
transform 1 0 1108 0 1 3985
box -3 -3 3 3
use M3_M2  M3_M2_2268
timestamp 1745462530
transform 1 0 1020 0 1 4215
box -3 -3 3 3
use M3_M2  M3_M2_2269
timestamp 1745462530
transform 1 0 940 0 1 3985
box -3 -3 3 3
use M3_M2  M3_M2_2270
timestamp 1745462530
transform 1 0 820 0 1 3985
box -3 -3 3 3
use M3_M2  M3_M2_2271
timestamp 1745462530
transform 1 0 756 0 1 4195
box -3 -3 3 3
use M3_M2  M3_M2_2272
timestamp 1745462530
transform 1 0 748 0 1 3985
box -3 -3 3 3
use M3_M2  M3_M2_2273
timestamp 1745462530
transform 1 0 732 0 1 4195
box -3 -3 3 3
use M3_M2  M3_M2_2274
timestamp 1745462530
transform 1 0 644 0 1 3985
box -3 -3 3 3
use M3_M2  M3_M2_2275
timestamp 1745462530
transform 1 0 3356 0 1 3985
box -3 -3 3 3
use M3_M2  M3_M2_2276
timestamp 1745462530
transform 1 0 3252 0 1 3865
box -3 -3 3 3
use M3_M2  M3_M2_2277
timestamp 1745462530
transform 1 0 3244 0 1 3985
box -3 -3 3 3
use M3_M2  M3_M2_2278
timestamp 1745462530
transform 1 0 3220 0 1 3985
box -3 -3 3 3
use M3_M2  M3_M2_2279
timestamp 1745462530
transform 1 0 3220 0 1 3865
box -3 -3 3 3
use M3_M2  M3_M2_2280
timestamp 1745462530
transform 1 0 3124 0 1 4015
box -3 -3 3 3
use M3_M2  M3_M2_2281
timestamp 1745462530
transform 1 0 3124 0 1 3985
box -3 -3 3 3
use M3_M2  M3_M2_2282
timestamp 1745462530
transform 1 0 2492 0 1 4035
box -3 -3 3 3
use M3_M2  M3_M2_2283
timestamp 1745462530
transform 1 0 2492 0 1 4005
box -3 -3 3 3
use M3_M2  M3_M2_2284
timestamp 1745462530
transform 1 0 2068 0 1 4035
box -3 -3 3 3
use M3_M2  M3_M2_2285
timestamp 1745462530
transform 1 0 1356 0 1 4035
box -3 -3 3 3
use M3_M2  M3_M2_2286
timestamp 1745462530
transform 1 0 1356 0 1 3875
box -3 -3 3 3
use M3_M2  M3_M2_2287
timestamp 1745462530
transform 1 0 996 0 1 3875
box -3 -3 3 3
use M3_M2  M3_M2_2288
timestamp 1745462530
transform 1 0 996 0 1 3765
box -3 -3 3 3
use M3_M2  M3_M2_2289
timestamp 1745462530
transform 1 0 868 0 1 3755
box -3 -3 3 3
use M3_M2  M3_M2_2290
timestamp 1745462530
transform 1 0 556 0 1 3755
box -3 -3 3 3
use M3_M2  M3_M2_2291
timestamp 1745462530
transform 1 0 380 0 1 3755
box -3 -3 3 3
use M3_M2  M3_M2_2292
timestamp 1745462530
transform 1 0 356 0 1 4195
box -3 -3 3 3
use M3_M2  M3_M2_2293
timestamp 1745462530
transform 1 0 244 0 1 4195
box -3 -3 3 3
use M3_M2  M3_M2_2294
timestamp 1745462530
transform 1 0 3876 0 1 3975
box -3 -3 3 3
use M3_M2  M3_M2_2295
timestamp 1745462530
transform 1 0 3836 0 1 3975
box -3 -3 3 3
use M3_M2  M3_M2_2296
timestamp 1745462530
transform 1 0 3748 0 1 3975
box -3 -3 3 3
use M3_M2  M3_M2_2297
timestamp 1745462530
transform 1 0 3636 0 1 4295
box -3 -3 3 3
use M3_M2  M3_M2_2298
timestamp 1745462530
transform 1 0 3636 0 1 3975
box -3 -3 3 3
use M3_M2  M3_M2_2299
timestamp 1745462530
transform 1 0 3604 0 1 3975
box -3 -3 3 3
use M3_M2  M3_M2_2300
timestamp 1745462530
transform 1 0 3596 0 1 4165
box -3 -3 3 3
use M3_M2  M3_M2_2301
timestamp 1745462530
transform 1 0 3572 0 1 4295
box -3 -3 3 3
use M3_M2  M3_M2_2302
timestamp 1745462530
transform 1 0 3572 0 1 4165
box -3 -3 3 3
use M3_M2  M3_M2_2303
timestamp 1745462530
transform 1 0 3396 0 1 4295
box -3 -3 3 3
use M3_M2  M3_M2_2304
timestamp 1745462530
transform 1 0 3388 0 1 4195
box -3 -3 3 3
use M3_M2  M3_M2_2305
timestamp 1745462530
transform 1 0 3292 0 1 4195
box -3 -3 3 3
use M3_M2  M3_M2_2306
timestamp 1745462530
transform 1 0 3100 0 1 4195
box -3 -3 3 3
use M3_M2  M3_M2_2307
timestamp 1745462530
transform 1 0 3084 0 1 4125
box -3 -3 3 3
use M3_M2  M3_M2_2308
timestamp 1745462530
transform 1 0 2812 0 1 4125
box -3 -3 3 3
use M3_M2  M3_M2_2309
timestamp 1745462530
transform 1 0 2812 0 1 4065
box -3 -3 3 3
use M3_M2  M3_M2_2310
timestamp 1745462530
transform 1 0 2748 0 1 4065
box -3 -3 3 3
use M3_M2  M3_M2_2311
timestamp 1745462530
transform 1 0 2460 0 1 4065
box -3 -3 3 3
use M3_M2  M3_M2_2312
timestamp 1745462530
transform 1 0 2252 0 1 4065
box -3 -3 3 3
use M3_M2  M3_M2_2313
timestamp 1745462530
transform 1 0 3924 0 1 4265
box -3 -3 3 3
use M3_M2  M3_M2_2314
timestamp 1745462530
transform 1 0 3908 0 1 3955
box -3 -3 3 3
use M3_M2  M3_M2_2315
timestamp 1745462530
transform 1 0 3844 0 1 3955
box -3 -3 3 3
use M3_M2  M3_M2_2316
timestamp 1745462530
transform 1 0 3764 0 1 3955
box -3 -3 3 3
use M3_M2  M3_M2_2317
timestamp 1745462530
transform 1 0 3732 0 1 4305
box -3 -3 3 3
use M3_M2  M3_M2_2318
timestamp 1745462530
transform 1 0 3732 0 1 4265
box -3 -3 3 3
use M3_M2  M3_M2_2319
timestamp 1745462530
transform 1 0 3196 0 1 4285
box -3 -3 3 3
use M3_M2  M3_M2_2320
timestamp 1745462530
transform 1 0 2908 0 1 4185
box -3 -3 3 3
use M3_M2  M3_M2_2321
timestamp 1745462530
transform 1 0 2860 0 1 4185
box -3 -3 3 3
use M3_M2  M3_M2_2322
timestamp 1745462530
transform 1 0 2772 0 1 4185
box -3 -3 3 3
use M3_M2  M3_M2_2323
timestamp 1745462530
transform 1 0 2764 0 1 4315
box -3 -3 3 3
use M3_M2  M3_M2_2324
timestamp 1745462530
transform 1 0 2764 0 1 4285
box -3 -3 3 3
use M3_M2  M3_M2_2325
timestamp 1745462530
transform 1 0 2556 0 1 4195
box -3 -3 3 3
use M3_M2  M3_M2_2326
timestamp 1745462530
transform 1 0 2444 0 1 4315
box -3 -3 3 3
use M3_M2  M3_M2_2327
timestamp 1745462530
transform 1 0 2444 0 1 4195
box -3 -3 3 3
use M3_M2  M3_M2_2328
timestamp 1745462530
transform 1 0 2348 0 1 4315
box -3 -3 3 3
use M3_M2  M3_M2_2329
timestamp 1745462530
transform 1 0 2212 0 1 4315
box -3 -3 3 3
use M3_M2  M3_M2_2330
timestamp 1745462530
transform 1 0 2036 0 1 4315
box -3 -3 3 3
use M3_M2  M3_M2_2331
timestamp 1745462530
transform 1 0 4284 0 1 3925
box -3 -3 3 3
use M3_M2  M3_M2_2332
timestamp 1745462530
transform 1 0 4284 0 1 3575
box -3 -3 3 3
use M3_M2  M3_M2_2333
timestamp 1745462530
transform 1 0 4164 0 1 3575
box -3 -3 3 3
use M3_M2  M3_M2_2334
timestamp 1745462530
transform 1 0 4116 0 1 3575
box -3 -3 3 3
use M3_M2  M3_M2_2335
timestamp 1745462530
transform 1 0 4068 0 1 3575
box -3 -3 3 3
use M3_M2  M3_M2_2336
timestamp 1745462530
transform 1 0 3988 0 1 3995
box -3 -3 3 3
use M3_M2  M3_M2_2337
timestamp 1745462530
transform 1 0 3988 0 1 3925
box -3 -3 3 3
use M3_M2  M3_M2_2338
timestamp 1745462530
transform 1 0 3932 0 1 3575
box -3 -3 3 3
use M3_M2  M3_M2_2339
timestamp 1745462530
transform 1 0 2956 0 1 3995
box -3 -3 3 3
use M3_M2  M3_M2_2340
timestamp 1745462530
transform 1 0 2956 0 1 3955
box -3 -3 3 3
use M3_M2  M3_M2_2341
timestamp 1745462530
transform 1 0 2908 0 1 3955
box -3 -3 3 3
use M3_M2  M3_M2_2342
timestamp 1745462530
transform 1 0 2892 0 1 4015
box -3 -3 3 3
use M3_M2  M3_M2_2343
timestamp 1745462530
transform 1 0 2892 0 1 3955
box -3 -3 3 3
use M3_M2  M3_M2_2344
timestamp 1745462530
transform 1 0 2572 0 1 4015
box -3 -3 3 3
use M3_M2  M3_M2_2345
timestamp 1745462530
transform 1 0 1980 0 1 4015
box -3 -3 3 3
use M3_M2  M3_M2_2346
timestamp 1745462530
transform 1 0 1916 0 1 4015
box -3 -3 3 3
use M3_M2  M3_M2_2347
timestamp 1745462530
transform 1 0 4340 0 1 4155
box -3 -3 3 3
use M3_M2  M3_M2_2348
timestamp 1745462530
transform 1 0 4332 0 1 3485
box -3 -3 3 3
use M3_M2  M3_M2_2349
timestamp 1745462530
transform 1 0 4292 0 1 3485
box -3 -3 3 3
use M3_M2  M3_M2_2350
timestamp 1745462530
transform 1 0 4284 0 1 3155
box -3 -3 3 3
use M3_M2  M3_M2_2351
timestamp 1745462530
transform 1 0 4100 0 1 3245
box -3 -3 3 3
use M3_M2  M3_M2_2352
timestamp 1745462530
transform 1 0 4100 0 1 3155
box -3 -3 3 3
use M3_M2  M3_M2_2353
timestamp 1745462530
transform 1 0 4020 0 1 3155
box -3 -3 3 3
use M3_M2  M3_M2_2354
timestamp 1745462530
transform 1 0 3924 0 1 3245
box -3 -3 3 3
use M3_M2  M3_M2_2355
timestamp 1745462530
transform 1 0 1932 0 1 4155
box -3 -3 3 3
use M3_M2  M3_M2_2356
timestamp 1745462530
transform 1 0 1828 0 1 4015
box -3 -3 3 3
use M3_M2  M3_M2_2357
timestamp 1745462530
transform 1 0 1748 0 1 4145
box -3 -3 3 3
use M3_M2  M3_M2_2358
timestamp 1745462530
transform 1 0 1620 0 1 4145
box -3 -3 3 3
use M3_M2  M3_M2_2359
timestamp 1745462530
transform 1 0 1620 0 1 4015
box -3 -3 3 3
use M3_M2  M3_M2_2360
timestamp 1745462530
transform 1 0 1516 0 1 3945
box -3 -3 3 3
use M3_M2  M3_M2_2361
timestamp 1745462530
transform 1 0 1500 0 1 4015
box -3 -3 3 3
use M3_M2  M3_M2_2362
timestamp 1745462530
transform 1 0 1500 0 1 3945
box -3 -3 3 3
use M3_M2  M3_M2_2363
timestamp 1745462530
transform 1 0 1388 0 1 3945
box -3 -3 3 3
use M3_M2  M3_M2_2364
timestamp 1745462530
transform 1 0 4284 0 1 2745
box -3 -3 3 3
use M3_M2  M3_M2_2365
timestamp 1745462530
transform 1 0 4252 0 1 3105
box -3 -3 3 3
use M3_M2  M3_M2_2366
timestamp 1745462530
transform 1 0 4252 0 1 2955
box -3 -3 3 3
use M3_M2  M3_M2_2367
timestamp 1745462530
transform 1 0 4188 0 1 2955
box -3 -3 3 3
use M3_M2  M3_M2_2368
timestamp 1745462530
transform 1 0 4188 0 1 2745
box -3 -3 3 3
use M3_M2  M3_M2_2369
timestamp 1745462530
transform 1 0 4092 0 1 3455
box -3 -3 3 3
use M3_M2  M3_M2_2370
timestamp 1745462530
transform 1 0 4084 0 1 3105
box -3 -3 3 3
use M3_M2  M3_M2_2371
timestamp 1745462530
transform 1 0 4068 0 1 3605
box -3 -3 3 3
use M3_M2  M3_M2_2372
timestamp 1745462530
transform 1 0 4052 0 1 3455
box -3 -3 3 3
use M3_M2  M3_M2_2373
timestamp 1745462530
transform 1 0 3908 0 1 3625
box -3 -3 3 3
use M3_M2  M3_M2_2374
timestamp 1745462530
transform 1 0 3020 0 1 3795
box -3 -3 3 3
use M3_M2  M3_M2_2375
timestamp 1745462530
transform 1 0 2916 0 1 2955
box -3 -3 3 3
use M3_M2  M3_M2_2376
timestamp 1745462530
transform 1 0 2908 0 1 2915
box -3 -3 3 3
use M3_M2  M3_M2_2377
timestamp 1745462530
transform 1 0 2868 0 1 3715
box -3 -3 3 3
use M3_M2  M3_M2_2378
timestamp 1745462530
transform 1 0 2852 0 1 3405
box -3 -3 3 3
use M3_M2  M3_M2_2379
timestamp 1745462530
transform 1 0 2836 0 1 3795
box -3 -3 3 3
use M3_M2  M3_M2_2380
timestamp 1745462530
transform 1 0 2836 0 1 3725
box -3 -3 3 3
use M3_M2  M3_M2_2381
timestamp 1745462530
transform 1 0 2804 0 1 3405
box -3 -3 3 3
use M3_M2  M3_M2_2382
timestamp 1745462530
transform 1 0 2788 0 1 3815
box -3 -3 3 3
use M3_M2  M3_M2_2383
timestamp 1745462530
transform 1 0 2772 0 1 2915
box -3 -3 3 3
use M3_M2  M3_M2_2384
timestamp 1745462530
transform 1 0 1460 0 1 3815
box -3 -3 3 3
use M3_M2  M3_M2_2385
timestamp 1745462530
transform 1 0 1348 0 1 3815
box -3 -3 3 3
use M3_M2  M3_M2_2386
timestamp 1745462530
transform 1 0 4372 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_2387
timestamp 1745462530
transform 1 0 4372 0 1 1885
box -3 -3 3 3
use M3_M2  M3_M2_2388
timestamp 1745462530
transform 1 0 4284 0 1 2215
box -3 -3 3 3
use M3_M2  M3_M2_2389
timestamp 1745462530
transform 1 0 4284 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_2390
timestamp 1745462530
transform 1 0 4268 0 1 1885
box -3 -3 3 3
use M3_M2  M3_M2_2391
timestamp 1745462530
transform 1 0 4236 0 1 2865
box -3 -3 3 3
use M3_M2  M3_M2_2392
timestamp 1745462530
transform 1 0 4236 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_2393
timestamp 1745462530
transform 1 0 4236 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_2394
timestamp 1745462530
transform 1 0 4236 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_2395
timestamp 1745462530
transform 1 0 4212 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_2396
timestamp 1745462530
transform 1 0 4196 0 1 2215
box -3 -3 3 3
use M3_M2  M3_M2_2397
timestamp 1745462530
transform 1 0 4196 0 1 2045
box -3 -3 3 3
use M3_M2  M3_M2_2398
timestamp 1745462530
transform 1 0 4196 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_2399
timestamp 1745462530
transform 1 0 4188 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_2400
timestamp 1745462530
transform 1 0 4164 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_2401
timestamp 1745462530
transform 1 0 4092 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_2402
timestamp 1745462530
transform 1 0 4012 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_2403
timestamp 1745462530
transform 1 0 3996 0 1 2865
box -3 -3 3 3
use M3_M2  M3_M2_2404
timestamp 1745462530
transform 1 0 3980 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_2405
timestamp 1745462530
transform 1 0 3956 0 1 2215
box -3 -3 3 3
use M3_M2  M3_M2_2406
timestamp 1745462530
transform 1 0 3196 0 1 2215
box -3 -3 3 3
use M3_M2  M3_M2_2407
timestamp 1745462530
transform 1 0 3004 0 1 2215
box -3 -3 3 3
use M3_M2  M3_M2_2408
timestamp 1745462530
transform 1 0 4140 0 1 155
box -3 -3 3 3
use M3_M2  M3_M2_2409
timestamp 1745462530
transform 1 0 4036 0 1 155
box -3 -3 3 3
use M3_M2  M3_M2_2410
timestamp 1745462530
transform 1 0 3916 0 1 155
box -3 -3 3 3
use M3_M2  M3_M2_2411
timestamp 1745462530
transform 1 0 3348 0 1 155
box -3 -3 3 3
use M3_M2  M3_M2_2412
timestamp 1745462530
transform 1 0 3148 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_2413
timestamp 1745462530
transform 1 0 3148 0 1 815
box -3 -3 3 3
use M3_M2  M3_M2_2414
timestamp 1745462530
transform 1 0 3124 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_2415
timestamp 1745462530
transform 1 0 3124 0 1 155
box -3 -3 3 3
use M3_M2  M3_M2_2416
timestamp 1745462530
transform 1 0 3116 0 1 535
box -3 -3 3 3
use M3_M2  M3_M2_2417
timestamp 1745462530
transform 1 0 3004 0 1 535
box -3 -3 3 3
use M3_M2  M3_M2_2418
timestamp 1745462530
transform 1 0 3004 0 1 155
box -3 -3 3 3
use M3_M2  M3_M2_2419
timestamp 1745462530
transform 1 0 2988 0 1 1335
box -3 -3 3 3
use M3_M2  M3_M2_2420
timestamp 1745462530
transform 1 0 2956 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_2421
timestamp 1745462530
transform 1 0 2916 0 1 1335
box -3 -3 3 3
use M3_M2  M3_M2_2422
timestamp 1745462530
transform 1 0 2908 0 1 155
box -3 -3 3 3
use M3_M2  M3_M2_2423
timestamp 1745462530
transform 1 0 2796 0 1 155
box -3 -3 3 3
use M3_M2  M3_M2_2424
timestamp 1745462530
transform 1 0 2148 0 1 1335
box -3 -3 3 3
use M3_M2  M3_M2_2425
timestamp 1745462530
transform 1 0 1852 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_2426
timestamp 1745462530
transform 1 0 1756 0 1 1045
box -3 -3 3 3
use M3_M2  M3_M2_2427
timestamp 1745462530
transform 1 0 1748 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_2428
timestamp 1745462530
transform 1 0 1748 0 1 465
box -3 -3 3 3
use M3_M2  M3_M2_2429
timestamp 1745462530
transform 1 0 1716 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_2430
timestamp 1745462530
transform 1 0 1716 0 1 465
box -3 -3 3 3
use M3_M2  M3_M2_2431
timestamp 1745462530
transform 1 0 1708 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_2432
timestamp 1745462530
transform 1 0 1700 0 1 1045
box -3 -3 3 3
use M3_M2  M3_M2_2433
timestamp 1745462530
transform 1 0 1676 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_2434
timestamp 1745462530
transform 1 0 1620 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_2435
timestamp 1745462530
transform 1 0 1604 0 1 465
box -3 -3 3 3
use M3_M2  M3_M2_2436
timestamp 1745462530
transform 1 0 1524 0 1 465
box -3 -3 3 3
use M3_M2  M3_M2_2437
timestamp 1745462530
transform 1 0 1356 0 1 465
box -3 -3 3 3
use M3_M2  M3_M2_2438
timestamp 1745462530
transform 1 0 732 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_2439
timestamp 1745462530
transform 1 0 732 0 1 465
box -3 -3 3 3
use M3_M2  M3_M2_2440
timestamp 1745462530
transform 1 0 692 0 1 1275
box -3 -3 3 3
use M3_M2  M3_M2_2441
timestamp 1745462530
transform 1 0 692 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_2442
timestamp 1745462530
transform 1 0 588 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_2443
timestamp 1745462530
transform 1 0 588 0 1 1275
box -3 -3 3 3
use M3_M2  M3_M2_2444
timestamp 1745462530
transform 1 0 572 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_2445
timestamp 1745462530
transform 1 0 548 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_2446
timestamp 1745462530
transform 1 0 1828 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_2447
timestamp 1745462530
transform 1 0 1732 0 1 1855
box -3 -3 3 3
use M3_M2  M3_M2_2448
timestamp 1745462530
transform 1 0 1724 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_2449
timestamp 1745462530
transform 1 0 1716 0 1 2355
box -3 -3 3 3
use M3_M2  M3_M2_2450
timestamp 1745462530
transform 1 0 1652 0 1 1855
box -3 -3 3 3
use M3_M2  M3_M2_2451
timestamp 1745462530
transform 1 0 1620 0 1 2355
box -3 -3 3 3
use M3_M2  M3_M2_2452
timestamp 1745462530
transform 1 0 908 0 1 2355
box -3 -3 3 3
use M3_M2  M3_M2_2453
timestamp 1745462530
transform 1 0 540 0 1 2415
box -3 -3 3 3
use M3_M2  M3_M2_2454
timestamp 1745462530
transform 1 0 540 0 1 2355
box -3 -3 3 3
use M3_M2  M3_M2_2455
timestamp 1745462530
transform 1 0 532 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_2456
timestamp 1745462530
transform 1 0 508 0 1 2415
box -3 -3 3 3
use M3_M2  M3_M2_2457
timestamp 1745462530
transform 1 0 324 0 1 2155
box -3 -3 3 3
use M3_M2  M3_M2_2458
timestamp 1745462530
transform 1 0 324 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_2459
timestamp 1745462530
transform 1 0 284 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_2460
timestamp 1745462530
transform 1 0 260 0 1 2555
box -3 -3 3 3
use M3_M2  M3_M2_2461
timestamp 1745462530
transform 1 0 220 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_2462
timestamp 1745462530
transform 1 0 220 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_2463
timestamp 1745462530
transform 1 0 212 0 1 2295
box -3 -3 3 3
use M3_M2  M3_M2_2464
timestamp 1745462530
transform 1 0 212 0 1 2165
box -3 -3 3 3
use M3_M2  M3_M2_2465
timestamp 1745462530
transform 1 0 204 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_2466
timestamp 1745462530
transform 1 0 196 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_2467
timestamp 1745462530
transform 1 0 156 0 1 2555
box -3 -3 3 3
use M3_M2  M3_M2_2468
timestamp 1745462530
transform 1 0 156 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_2469
timestamp 1745462530
transform 1 0 156 0 1 2295
box -3 -3 3 3
use M3_M2  M3_M2_2470
timestamp 1745462530
transform 1 0 140 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_2471
timestamp 1745462530
transform 1 0 132 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_2472
timestamp 1745462530
transform 1 0 100 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_2473
timestamp 1745462530
transform 1 0 92 0 1 2545
box -3 -3 3 3
use M3_M2  M3_M2_2474
timestamp 1745462530
transform 1 0 3716 0 1 2445
box -3 -3 3 3
use M3_M2  M3_M2_2475
timestamp 1745462530
transform 1 0 3708 0 1 2645
box -3 -3 3 3
use M3_M2  M3_M2_2476
timestamp 1745462530
transform 1 0 3692 0 1 2445
box -3 -3 3 3
use M3_M2  M3_M2_2477
timestamp 1745462530
transform 1 0 3676 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_2478
timestamp 1745462530
transform 1 0 3652 0 1 2645
box -3 -3 3 3
use M3_M2  M3_M2_2479
timestamp 1745462530
transform 1 0 3604 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_2480
timestamp 1745462530
transform 1 0 3572 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_2481
timestamp 1745462530
transform 1 0 3476 0 1 2645
box -3 -3 3 3
use M3_M2  M3_M2_2482
timestamp 1745462530
transform 1 0 3476 0 1 2475
box -3 -3 3 3
use M3_M2  M3_M2_2483
timestamp 1745462530
transform 1 0 3468 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_2484
timestamp 1745462530
transform 1 0 2988 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_2485
timestamp 1745462530
transform 1 0 2988 0 1 2475
box -3 -3 3 3
use M3_M2  M3_M2_2486
timestamp 1745462530
transform 1 0 2964 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_2487
timestamp 1745462530
transform 1 0 2836 0 1 2475
box -3 -3 3 3
use M3_M2  M3_M2_2488
timestamp 1745462530
transform 1 0 2836 0 1 2445
box -3 -3 3 3
use M3_M2  M3_M2_2489
timestamp 1745462530
transform 1 0 2524 0 1 2445
box -3 -3 3 3
use M3_M2  M3_M2_2490
timestamp 1745462530
transform 1 0 2204 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_2491
timestamp 1745462530
transform 1 0 2084 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_2492
timestamp 1745462530
transform 1 0 2084 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_2493
timestamp 1745462530
transform 1 0 2068 0 1 2445
box -3 -3 3 3
use M3_M2  M3_M2_2494
timestamp 1745462530
transform 1 0 2052 0 1 2535
box -3 -3 3 3
use M3_M2  M3_M2_2495
timestamp 1745462530
transform 1 0 2044 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_2496
timestamp 1745462530
transform 1 0 2012 0 1 2535
box -3 -3 3 3
use M3_M2  M3_M2_2497
timestamp 1745462530
transform 1 0 1996 0 1 2725
box -3 -3 3 3
use M3_M2  M3_M2_2498
timestamp 1745462530
transform 1 0 1956 0 1 3035
box -3 -3 3 3
use M3_M2  M3_M2_2499
timestamp 1745462530
transform 1 0 1940 0 1 2725
box -3 -3 3 3
use M3_M2  M3_M2_2500
timestamp 1745462530
transform 1 0 1916 0 1 3035
box -3 -3 3 3
use M3_M2  M3_M2_2501
timestamp 1745462530
transform 1 0 4292 0 1 2155
box -3 -3 3 3
use M3_M2  M3_M2_2502
timestamp 1745462530
transform 1 0 4284 0 1 865
box -3 -3 3 3
use M3_M2  M3_M2_2503
timestamp 1745462530
transform 1 0 4092 0 1 865
box -3 -3 3 3
use M3_M2  M3_M2_2504
timestamp 1745462530
transform 1 0 4068 0 1 1215
box -3 -3 3 3
use M3_M2  M3_M2_2505
timestamp 1745462530
transform 1 0 3716 0 1 2155
box -3 -3 3 3
use M3_M2  M3_M2_2506
timestamp 1745462530
transform 1 0 3668 0 1 2545
box -3 -3 3 3
use M3_M2  M3_M2_2507
timestamp 1745462530
transform 1 0 3652 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_2508
timestamp 1745462530
transform 1 0 3652 0 1 1215
box -3 -3 3 3
use M3_M2  M3_M2_2509
timestamp 1745462530
transform 1 0 3652 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_2510
timestamp 1745462530
transform 1 0 3644 0 1 2155
box -3 -3 3 3
use M3_M2  M3_M2_2511
timestamp 1745462530
transform 1 0 3644 0 1 2015
box -3 -3 3 3
use M3_M2  M3_M2_2512
timestamp 1745462530
transform 1 0 3636 0 1 2545
box -3 -3 3 3
use M3_M2  M3_M2_2513
timestamp 1745462530
transform 1 0 3604 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_2514
timestamp 1745462530
transform 1 0 3548 0 1 2015
box -3 -3 3 3
use M3_M2  M3_M2_2515
timestamp 1745462530
transform 1 0 3548 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_2516
timestamp 1745462530
transform 1 0 2820 0 1 2015
box -3 -3 3 3
use M3_M2  M3_M2_2517
timestamp 1745462530
transform 1 0 2788 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_2518
timestamp 1745462530
transform 1 0 2788 0 1 2015
box -3 -3 3 3
use M3_M2  M3_M2_2519
timestamp 1745462530
transform 1 0 2620 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_2520
timestamp 1745462530
transform 1 0 2292 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_2521
timestamp 1745462530
transform 1 0 3684 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_2522
timestamp 1745462530
transform 1 0 3604 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_2523
timestamp 1745462530
transform 1 0 3572 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_2524
timestamp 1745462530
transform 1 0 3236 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_2525
timestamp 1745462530
transform 1 0 3012 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_2526
timestamp 1745462530
transform 1 0 2820 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_2527
timestamp 1745462530
transform 1 0 2780 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_2528
timestamp 1745462530
transform 1 0 2772 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_2529
timestamp 1745462530
transform 1 0 2724 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_2530
timestamp 1745462530
transform 1 0 2724 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_2531
timestamp 1745462530
transform 1 0 2708 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_2532
timestamp 1745462530
transform 1 0 2692 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_2533
timestamp 1745462530
transform 1 0 2692 0 1 125
box -3 -3 3 3
use M3_M2  M3_M2_2534
timestamp 1745462530
transform 1 0 2676 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_2535
timestamp 1745462530
transform 1 0 2676 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_2536
timestamp 1745462530
transform 1 0 2668 0 1 535
box -3 -3 3 3
use M3_M2  M3_M2_2537
timestamp 1745462530
transform 1 0 2556 0 1 125
box -3 -3 3 3
use M3_M2  M3_M2_2538
timestamp 1745462530
transform 1 0 2196 0 1 1575
box -3 -3 3 3
use M3_M2  M3_M2_2539
timestamp 1745462530
transform 1 0 2020 0 1 1575
box -3 -3 3 3
use M3_M2  M3_M2_2540
timestamp 1745462530
transform 1 0 1356 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_2541
timestamp 1745462530
transform 1 0 1284 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_2542
timestamp 1745462530
transform 1 0 1284 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_2543
timestamp 1745462530
transform 1 0 1276 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_2544
timestamp 1745462530
transform 1 0 1268 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_2545
timestamp 1745462530
transform 1 0 1252 0 1 215
box -3 -3 3 3
use M3_M2  M3_M2_2546
timestamp 1745462530
transform 1 0 1236 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_2547
timestamp 1745462530
transform 1 0 1236 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_2548
timestamp 1745462530
transform 1 0 1196 0 1 215
box -3 -3 3 3
use M3_M2  M3_M2_2549
timestamp 1745462530
transform 1 0 1196 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_2550
timestamp 1745462530
transform 1 0 1180 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_2551
timestamp 1745462530
transform 1 0 1116 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_2552
timestamp 1745462530
transform 1 0 1116 0 1 645
box -3 -3 3 3
use M3_M2  M3_M2_2553
timestamp 1745462530
transform 1 0 980 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_2554
timestamp 1745462530
transform 1 0 964 0 1 645
box -3 -3 3 3
use M3_M2  M3_M2_2555
timestamp 1745462530
transform 1 0 956 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_2556
timestamp 1745462530
transform 1 0 748 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_2557
timestamp 1745462530
transform 1 0 724 0 1 215
box -3 -3 3 3
use M3_M2  M3_M2_2558
timestamp 1745462530
transform 1 0 596 0 1 215
box -3 -3 3 3
use M3_M2  M3_M2_2559
timestamp 1745462530
transform 1 0 508 0 1 325
box -3 -3 3 3
use M3_M2  M3_M2_2560
timestamp 1745462530
transform 1 0 460 0 1 325
box -3 -3 3 3
use M3_M2  M3_M2_2561
timestamp 1745462530
transform 1 0 460 0 1 215
box -3 -3 3 3
use M3_M2  M3_M2_2562
timestamp 1745462530
transform 1 0 372 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_2563
timestamp 1745462530
transform 1 0 1380 0 1 2725
box -3 -3 3 3
use M3_M2  M3_M2_2564
timestamp 1745462530
transform 1 0 1380 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_2565
timestamp 1745462530
transform 1 0 1348 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_2566
timestamp 1745462530
transform 1 0 1340 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_2567
timestamp 1745462530
transform 1 0 980 0 1 2725
box -3 -3 3 3
use M3_M2  M3_M2_2568
timestamp 1745462530
transform 1 0 484 0 1 1815
box -3 -3 3 3
use M3_M2  M3_M2_2569
timestamp 1745462530
transform 1 0 476 0 1 2745
box -3 -3 3 3
use M3_M2  M3_M2_2570
timestamp 1745462530
transform 1 0 276 0 1 1415
box -3 -3 3 3
use M3_M2  M3_M2_2571
timestamp 1745462530
transform 1 0 116 0 1 1815
box -3 -3 3 3
use M3_M2  M3_M2_2572
timestamp 1745462530
transform 1 0 108 0 1 2375
box -3 -3 3 3
use M3_M2  M3_M2_2573
timestamp 1745462530
transform 1 0 92 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_2574
timestamp 1745462530
transform 1 0 92 0 1 1415
box -3 -3 3 3
use M3_M2  M3_M2_2575
timestamp 1745462530
transform 1 0 84 0 1 2745
box -3 -3 3 3
use M3_M2  M3_M2_2576
timestamp 1745462530
transform 1 0 84 0 1 2435
box -3 -3 3 3
use M3_M2  M3_M2_2577
timestamp 1745462530
transform 1 0 3268 0 1 2375
box -3 -3 3 3
use M3_M2  M3_M2_2578
timestamp 1745462530
transform 1 0 3236 0 1 2775
box -3 -3 3 3
use M3_M2  M3_M2_2579
timestamp 1745462530
transform 1 0 3164 0 1 2775
box -3 -3 3 3
use M3_M2  M3_M2_2580
timestamp 1745462530
transform 1 0 3148 0 1 2905
box -3 -3 3 3
use M3_M2  M3_M2_2581
timestamp 1745462530
transform 1 0 3132 0 1 2375
box -3 -3 3 3
use M3_M2  M3_M2_2582
timestamp 1745462530
transform 1 0 3132 0 1 2355
box -3 -3 3 3
use M3_M2  M3_M2_2583
timestamp 1745462530
transform 1 0 3060 0 1 2905
box -3 -3 3 3
use M3_M2  M3_M2_2584
timestamp 1745462530
transform 1 0 2884 0 1 2905
box -3 -3 3 3
use M3_M2  M3_M2_2585
timestamp 1745462530
transform 1 0 2884 0 1 2755
box -3 -3 3 3
use M3_M2  M3_M2_2586
timestamp 1745462530
transform 1 0 2748 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_2587
timestamp 1745462530
transform 1 0 2708 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_2588
timestamp 1745462530
transform 1 0 2708 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_2589
timestamp 1745462530
transform 1 0 2684 0 1 2755
box -3 -3 3 3
use M3_M2  M3_M2_2590
timestamp 1745462530
transform 1 0 2684 0 1 2355
box -3 -3 3 3
use M3_M2  M3_M2_2591
timestamp 1745462530
transform 1 0 1540 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_2592
timestamp 1745462530
transform 1 0 1444 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_2593
timestamp 1745462530
transform 1 0 4212 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_2594
timestamp 1745462530
transform 1 0 4204 0 1 675
box -3 -3 3 3
use M3_M2  M3_M2_2595
timestamp 1745462530
transform 1 0 4196 0 1 575
box -3 -3 3 3
use M3_M2  M3_M2_2596
timestamp 1745462530
transform 1 0 4124 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_2597
timestamp 1745462530
transform 1 0 4124 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_2598
timestamp 1745462530
transform 1 0 4116 0 1 575
box -3 -3 3 3
use M3_M2  M3_M2_2599
timestamp 1745462530
transform 1 0 4076 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_2600
timestamp 1745462530
transform 1 0 3988 0 1 675
box -3 -3 3 3
use M3_M2  M3_M2_2601
timestamp 1745462530
transform 1 0 3676 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_2602
timestamp 1745462530
transform 1 0 3668 0 1 1055
box -3 -3 3 3
use M3_M2  M3_M2_2603
timestamp 1745462530
transform 1 0 3644 0 1 1055
box -3 -3 3 3
use M3_M2  M3_M2_2604
timestamp 1745462530
transform 1 0 3636 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_2605
timestamp 1745462530
transform 1 0 3532 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_2606
timestamp 1745462530
transform 1 0 3532 0 1 675
box -3 -3 3 3
use M3_M2  M3_M2_2607
timestamp 1745462530
transform 1 0 3508 0 1 1525
box -3 -3 3 3
use M3_M2  M3_M2_2608
timestamp 1745462530
transform 1 0 3508 0 1 1295
box -3 -3 3 3
use M3_M2  M3_M2_2609
timestamp 1745462530
transform 1 0 3444 0 1 1525
box -3 -3 3 3
use M3_M2  M3_M2_2610
timestamp 1745462530
transform 1 0 3428 0 1 1525
box -3 -3 3 3
use M3_M2  M3_M2_2611
timestamp 1745462530
transform 1 0 3420 0 1 1655
box -3 -3 3 3
use M3_M2  M3_M2_2612
timestamp 1745462530
transform 1 0 3348 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_2613
timestamp 1745462530
transform 1 0 3348 0 1 675
box -3 -3 3 3
use M3_M2  M3_M2_2614
timestamp 1745462530
transform 1 0 3268 0 1 1295
box -3 -3 3 3
use M3_M2  M3_M2_2615
timestamp 1745462530
transform 1 0 3268 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_2616
timestamp 1745462530
transform 1 0 3260 0 1 1655
box -3 -3 3 3
use M3_M2  M3_M2_2617
timestamp 1745462530
transform 1 0 3260 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_2618
timestamp 1745462530
transform 1 0 3236 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_2619
timestamp 1745462530
transform 1 0 2788 0 1 1645
box -3 -3 3 3
use M3_M2  M3_M2_2620
timestamp 1745462530
transform 1 0 2228 0 1 1645
box -3 -3 3 3
use M3_M2  M3_M2_2621
timestamp 1745462530
transform 1 0 3140 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_2622
timestamp 1745462530
transform 1 0 3076 0 1 575
box -3 -3 3 3
use M3_M2  M3_M2_2623
timestamp 1745462530
transform 1 0 3076 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_2624
timestamp 1745462530
transform 1 0 3036 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_2625
timestamp 1745462530
transform 1 0 2980 0 1 845
box -3 -3 3 3
use M3_M2  M3_M2_2626
timestamp 1745462530
transform 1 0 2980 0 1 575
box -3 -3 3 3
use M3_M2  M3_M2_2627
timestamp 1745462530
transform 1 0 2924 0 1 1455
box -3 -3 3 3
use M3_M2  M3_M2_2628
timestamp 1745462530
transform 1 0 2908 0 1 845
box -3 -3 3 3
use M3_M2  M3_M2_2629
timestamp 1745462530
transform 1 0 2852 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_2630
timestamp 1745462530
transform 1 0 2724 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_2631
timestamp 1745462530
transform 1 0 2140 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_2632
timestamp 1745462530
transform 1 0 2140 0 1 1455
box -3 -3 3 3
use M3_M2  M3_M2_2633
timestamp 1745462530
transform 1 0 1716 0 1 1535
box -3 -3 3 3
use M3_M2  M3_M2_2634
timestamp 1745462530
transform 1 0 1700 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_2635
timestamp 1745462530
transform 1 0 1652 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_2636
timestamp 1745462530
transform 1 0 1652 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_2637
timestamp 1745462530
transform 1 0 1580 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_2638
timestamp 1745462530
transform 1 0 1564 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_2639
timestamp 1745462530
transform 1 0 1556 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_2640
timestamp 1745462530
transform 1 0 1524 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_2641
timestamp 1745462530
transform 1 0 1596 0 1 1375
box -3 -3 3 3
use M3_M2  M3_M2_2642
timestamp 1745462530
transform 1 0 1572 0 1 125
box -3 -3 3 3
use M3_M2  M3_M2_2643
timestamp 1745462530
transform 1 0 1556 0 1 375
box -3 -3 3 3
use M3_M2  M3_M2_2644
timestamp 1745462530
transform 1 0 1500 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_2645
timestamp 1745462530
transform 1 0 1500 0 1 375
box -3 -3 3 3
use M3_M2  M3_M2_2646
timestamp 1745462530
transform 1 0 1388 0 1 1375
box -3 -3 3 3
use M3_M2  M3_M2_2647
timestamp 1745462530
transform 1 0 1380 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_2648
timestamp 1745462530
transform 1 0 1380 0 1 125
box -3 -3 3 3
use M3_M2  M3_M2_2649
timestamp 1745462530
transform 1 0 1324 0 1 815
box -3 -3 3 3
use M3_M2  M3_M2_2650
timestamp 1745462530
transform 1 0 1324 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_2651
timestamp 1745462530
transform 1 0 1316 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_2652
timestamp 1745462530
transform 1 0 1292 0 1 815
box -3 -3 3 3
use M3_M2  M3_M2_2653
timestamp 1745462530
transform 1 0 1036 0 1 125
box -3 -3 3 3
use M3_M2  M3_M2_2654
timestamp 1745462530
transform 1 0 924 0 1 125
box -3 -3 3 3
use M3_M2  M3_M2_2655
timestamp 1745462530
transform 1 0 692 0 1 125
box -3 -3 3 3
use M3_M2  M3_M2_2656
timestamp 1745462530
transform 1 0 644 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_2657
timestamp 1745462530
transform 1 0 644 0 1 1375
box -3 -3 3 3
use M3_M2  M3_M2_2658
timestamp 1745462530
transform 1 0 572 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_2659
timestamp 1745462530
transform 1 0 444 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_2660
timestamp 1745462530
transform 1 0 388 0 1 325
box -3 -3 3 3
use M3_M2  M3_M2_2661
timestamp 1745462530
transform 1 0 308 0 1 325
box -3 -3 3 3
use M3_M2  M3_M2_2662
timestamp 1745462530
transform 1 0 308 0 1 125
box -3 -3 3 3
use M3_M2  M3_M2_2663
timestamp 1745462530
transform 1 0 1988 0 1 1865
box -3 -3 3 3
use M3_M2  M3_M2_2664
timestamp 1745462530
transform 1 0 1340 0 1 2905
box -3 -3 3 3
use M3_M2  M3_M2_2665
timestamp 1745462530
transform 1 0 1308 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_2666
timestamp 1745462530
transform 1 0 1300 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_2667
timestamp 1745462530
transform 1 0 1284 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_2668
timestamp 1745462530
transform 1 0 1236 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_2669
timestamp 1745462530
transform 1 0 1236 0 1 1865
box -3 -3 3 3
use M3_M2  M3_M2_2670
timestamp 1745462530
transform 1 0 1228 0 1 2905
box -3 -3 3 3
use M3_M2  M3_M2_2671
timestamp 1745462530
transform 1 0 1212 0 1 2685
box -3 -3 3 3
use M3_M2  M3_M2_2672
timestamp 1745462530
transform 1 0 1140 0 1 2685
box -3 -3 3 3
use M3_M2  M3_M2_2673
timestamp 1745462530
transform 1 0 1132 0 1 2715
box -3 -3 3 3
use M3_M2  M3_M2_2674
timestamp 1745462530
transform 1 0 1044 0 1 2725
box -3 -3 3 3
use M3_M2  M3_M2_2675
timestamp 1745462530
transform 1 0 1028 0 1 2785
box -3 -3 3 3
use M3_M2  M3_M2_2676
timestamp 1745462530
transform 1 0 996 0 1 2905
box -3 -3 3 3
use M3_M2  M3_M2_2677
timestamp 1745462530
transform 1 0 996 0 1 2785
box -3 -3 3 3
use M3_M2  M3_M2_2678
timestamp 1745462530
transform 1 0 972 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_2679
timestamp 1745462530
transform 1 0 972 0 1 1835
box -3 -3 3 3
use M3_M2  M3_M2_2680
timestamp 1745462530
transform 1 0 804 0 1 1835
box -3 -3 3 3
use M3_M2  M3_M2_2681
timestamp 1745462530
transform 1 0 564 0 1 2955
box -3 -3 3 3
use M3_M2  M3_M2_2682
timestamp 1745462530
transform 1 0 564 0 1 2905
box -3 -3 3 3
use M3_M2  M3_M2_2683
timestamp 1745462530
transform 1 0 468 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_2684
timestamp 1745462530
transform 1 0 468 0 1 1835
box -3 -3 3 3
use M3_M2  M3_M2_2685
timestamp 1745462530
transform 1 0 420 0 1 2545
box -3 -3 3 3
use M3_M2  M3_M2_2686
timestamp 1745462530
transform 1 0 412 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_2687
timestamp 1745462530
transform 1 0 348 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_2688
timestamp 1745462530
transform 1 0 332 0 1 2945
box -3 -3 3 3
use M3_M2  M3_M2_2689
timestamp 1745462530
transform 1 0 276 0 1 2545
box -3 -3 3 3
use M3_M2  M3_M2_2690
timestamp 1745462530
transform 1 0 268 0 1 2945
box -3 -3 3 3
use M3_M2  M3_M2_2691
timestamp 1745462530
transform 1 0 188 0 1 2945
box -3 -3 3 3
use M3_M2  M3_M2_2692
timestamp 1745462530
transform 1 0 4292 0 1 2945
box -3 -3 3 3
use M3_M2  M3_M2_2693
timestamp 1745462530
transform 1 0 4292 0 1 2585
box -3 -3 3 3
use M3_M2  M3_M2_2694
timestamp 1745462530
transform 1 0 4276 0 1 2335
box -3 -3 3 3
use M3_M2  M3_M2_2695
timestamp 1745462530
transform 1 0 4268 0 1 2585
box -3 -3 3 3
use M3_M2  M3_M2_2696
timestamp 1745462530
transform 1 0 4252 0 1 2585
box -3 -3 3 3
use M3_M2  M3_M2_2697
timestamp 1745462530
transform 1 0 4164 0 1 2335
box -3 -3 3 3
use M3_M2  M3_M2_2698
timestamp 1745462530
transform 1 0 4164 0 1 2255
box -3 -3 3 3
use M3_M2  M3_M2_2699
timestamp 1745462530
transform 1 0 4116 0 1 2945
box -3 -3 3 3
use M3_M2  M3_M2_2700
timestamp 1745462530
transform 1 0 3964 0 1 2945
box -3 -3 3 3
use M3_M2  M3_M2_2701
timestamp 1745462530
transform 1 0 3308 0 1 2255
box -3 -3 3 3
use M3_M2  M3_M2_2702
timestamp 1745462530
transform 1 0 3108 0 1 2335
box -3 -3 3 3
use M3_M2  M3_M2_2703
timestamp 1745462530
transform 1 0 3108 0 1 2255
box -3 -3 3 3
use M3_M2  M3_M2_2704
timestamp 1745462530
transform 1 0 2860 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_2705
timestamp 1745462530
transform 1 0 2852 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_2706
timestamp 1745462530
transform 1 0 2788 0 1 2475
box -3 -3 3 3
use M3_M2  M3_M2_2707
timestamp 1745462530
transform 1 0 2788 0 1 2325
box -3 -3 3 3
use M3_M2  M3_M2_2708
timestamp 1745462530
transform 1 0 2788 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_2709
timestamp 1745462530
transform 1 0 2788 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_2710
timestamp 1745462530
transform 1 0 2788 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_2711
timestamp 1745462530
transform 1 0 2748 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_2712
timestamp 1745462530
transform 1 0 2748 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_2713
timestamp 1745462530
transform 1 0 2724 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_2714
timestamp 1745462530
transform 1 0 2724 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_2715
timestamp 1745462530
transform 1 0 2700 0 1 2655
box -3 -3 3 3
use M3_M2  M3_M2_2716
timestamp 1745462530
transform 1 0 2700 0 1 2475
box -3 -3 3 3
use M3_M2  M3_M2_2717
timestamp 1745462530
transform 1 0 2620 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_2718
timestamp 1745462530
transform 1 0 2620 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_2719
timestamp 1745462530
transform 1 0 2556 0 1 2755
box -3 -3 3 3
use M3_M2  M3_M2_2720
timestamp 1745462530
transform 1 0 2556 0 1 2655
box -3 -3 3 3
use M3_M2  M3_M2_2721
timestamp 1745462530
transform 1 0 2540 0 1 2905
box -3 -3 3 3
use M3_M2  M3_M2_2722
timestamp 1745462530
transform 1 0 2540 0 1 2755
box -3 -3 3 3
use M3_M2  M3_M2_2723
timestamp 1745462530
transform 1 0 2540 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_2724
timestamp 1745462530
transform 1 0 2508 0 1 2905
box -3 -3 3 3
use M3_M2  M3_M2_2725
timestamp 1745462530
transform 1 0 2308 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_2726
timestamp 1745462530
transform 1 0 1124 0 1 2915
box -3 -3 3 3
use M3_M2  M3_M2_2727
timestamp 1745462530
transform 1 0 4364 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_2728
timestamp 1745462530
transform 1 0 4364 0 1 375
box -3 -3 3 3
use M3_M2  M3_M2_2729
timestamp 1745462530
transform 1 0 4356 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_2730
timestamp 1745462530
transform 1 0 4292 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_2731
timestamp 1745462530
transform 1 0 4292 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_2732
timestamp 1745462530
transform 1 0 4292 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_2733
timestamp 1745462530
transform 1 0 4284 0 1 1675
box -3 -3 3 3
use M3_M2  M3_M2_2734
timestamp 1745462530
transform 1 0 4284 0 1 375
box -3 -3 3 3
use M3_M2  M3_M2_2735
timestamp 1745462530
transform 1 0 4276 0 1 125
box -3 -3 3 3
use M3_M2  M3_M2_2736
timestamp 1745462530
transform 1 0 4068 0 1 125
box -3 -3 3 3
use M3_M2  M3_M2_2737
timestamp 1745462530
transform 1 0 3996 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_2738
timestamp 1745462530
transform 1 0 3804 0 1 125
box -3 -3 3 3
use M3_M2  M3_M2_2739
timestamp 1745462530
transform 1 0 3628 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_2740
timestamp 1745462530
transform 1 0 3604 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_2741
timestamp 1745462530
transform 1 0 3572 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_2742
timestamp 1745462530
transform 1 0 3572 0 1 1675
box -3 -3 3 3
use M3_M2  M3_M2_2743
timestamp 1745462530
transform 1 0 3460 0 1 125
box -3 -3 3 3
use M3_M2  M3_M2_2744
timestamp 1745462530
transform 1 0 2276 0 1 1675
box -3 -3 3 3
use M3_M2  M3_M2_2745
timestamp 1745462530
transform 1 0 2356 0 1 125
box -3 -3 3 3
use M3_M2  M3_M2_2746
timestamp 1745462530
transform 1 0 2228 0 1 1275
box -3 -3 3 3
use M3_M2  M3_M2_2747
timestamp 1745462530
transform 1 0 2228 0 1 125
box -3 -3 3 3
use M3_M2  M3_M2_2748
timestamp 1745462530
transform 1 0 2188 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_2749
timestamp 1745462530
transform 1 0 2188 0 1 1275
box -3 -3 3 3
use M3_M2  M3_M2_2750
timestamp 1745462530
transform 1 0 2172 0 1 865
box -3 -3 3 3
use M3_M2  M3_M2_2751
timestamp 1745462530
transform 1 0 2092 0 1 125
box -3 -3 3 3
use M3_M2  M3_M2_2752
timestamp 1745462530
transform 1 0 2076 0 1 865
box -3 -3 3 3
use M3_M2  M3_M2_2753
timestamp 1745462530
transform 1 0 1988 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_2754
timestamp 1745462530
transform 1 0 1980 0 1 125
box -3 -3 3 3
use M3_M2  M3_M2_2755
timestamp 1745462530
transform 1 0 1948 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_2756
timestamp 1745462530
transform 1 0 1948 0 1 865
box -3 -3 3 3
use M3_M2  M3_M2_2757
timestamp 1745462530
transform 1 0 1900 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_2758
timestamp 1745462530
transform 1 0 1892 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_2759
timestamp 1745462530
transform 1 0 1820 0 1 865
box -3 -3 3 3
use M3_M2  M3_M2_2760
timestamp 1745462530
transform 1 0 1972 0 1 1575
box -3 -3 3 3
use M3_M2  M3_M2_2761
timestamp 1745462530
transform 1 0 1788 0 1 165
box -3 -3 3 3
use M3_M2  M3_M2_2762
timestamp 1745462530
transform 1 0 1676 0 1 165
box -3 -3 3 3
use M3_M2  M3_M2_2763
timestamp 1745462530
transform 1 0 812 0 1 155
box -3 -3 3 3
use M3_M2  M3_M2_2764
timestamp 1745462530
transform 1 0 668 0 1 1575
box -3 -3 3 3
use M3_M2  M3_M2_2765
timestamp 1745462530
transform 1 0 668 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_2766
timestamp 1745462530
transform 1 0 548 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_2767
timestamp 1745462530
transform 1 0 436 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_2768
timestamp 1745462530
transform 1 0 428 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_2769
timestamp 1745462530
transform 1 0 332 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_2770
timestamp 1745462530
transform 1 0 332 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_2771
timestamp 1745462530
transform 1 0 292 0 1 275
box -3 -3 3 3
use M3_M2  M3_M2_2772
timestamp 1745462530
transform 1 0 292 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_2773
timestamp 1745462530
transform 1 0 276 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_2774
timestamp 1745462530
transform 1 0 276 0 1 975
box -3 -3 3 3
use M3_M2  M3_M2_2775
timestamp 1745462530
transform 1 0 268 0 1 275
box -3 -3 3 3
use M3_M2  M3_M2_2776
timestamp 1745462530
transform 1 0 260 0 1 975
box -3 -3 3 3
use M3_M2  M3_M2_2777
timestamp 1745462530
transform 1 0 172 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_2778
timestamp 1745462530
transform 1 0 2380 0 1 2935
box -3 -3 3 3
use M3_M2  M3_M2_2779
timestamp 1745462530
transform 1 0 2060 0 1 2935
box -3 -3 3 3
use M3_M2  M3_M2_2780
timestamp 1745462530
transform 1 0 2060 0 1 2885
box -3 -3 3 3
use M3_M2  M3_M2_2781
timestamp 1745462530
transform 1 0 1972 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_2782
timestamp 1745462530
transform 1 0 1748 0 1 2585
box -3 -3 3 3
use M3_M2  M3_M2_2783
timestamp 1745462530
transform 1 0 1724 0 1 2885
box -3 -3 3 3
use M3_M2  M3_M2_2784
timestamp 1745462530
transform 1 0 1676 0 1 2605
box -3 -3 3 3
use M3_M2  M3_M2_2785
timestamp 1745462530
transform 1 0 1676 0 1 2585
box -3 -3 3 3
use M3_M2  M3_M2_2786
timestamp 1745462530
transform 1 0 1676 0 1 2065
box -3 -3 3 3
use M3_M2  M3_M2_2787
timestamp 1745462530
transform 1 0 1660 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_2788
timestamp 1745462530
transform 1 0 1652 0 1 2065
box -3 -3 3 3
use M3_M2  M3_M2_2789
timestamp 1745462530
transform 1 0 1612 0 1 2445
box -3 -3 3 3
use M3_M2  M3_M2_2790
timestamp 1745462530
transform 1 0 1596 0 1 2605
box -3 -3 3 3
use M3_M2  M3_M2_2791
timestamp 1745462530
transform 1 0 1596 0 1 2445
box -3 -3 3 3
use M3_M2  M3_M2_2792
timestamp 1745462530
transform 1 0 1548 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_2793
timestamp 1745462530
transform 1 0 1012 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_2794
timestamp 1745462530
transform 1 0 428 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_2795
timestamp 1745462530
transform 1 0 404 0 1 2625
box -3 -3 3 3
use M3_M2  M3_M2_2796
timestamp 1745462530
transform 1 0 404 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_2797
timestamp 1745462530
transform 1 0 404 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_2798
timestamp 1745462530
transform 1 0 308 0 1 2625
box -3 -3 3 3
use M3_M2  M3_M2_2799
timestamp 1745462530
transform 1 0 212 0 1 2625
box -3 -3 3 3
use M3_M2  M3_M2_2800
timestamp 1745462530
transform 1 0 4380 0 1 2275
box -3 -3 3 3
use M3_M2  M3_M2_2801
timestamp 1745462530
transform 1 0 4380 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_2802
timestamp 1745462530
transform 1 0 4316 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_2803
timestamp 1745462530
transform 1 0 4316 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_2804
timestamp 1745462530
transform 1 0 3988 0 1 1655
box -3 -3 3 3
use M3_M2  M3_M2_2805
timestamp 1745462530
transform 1 0 3980 0 1 2415
box -3 -3 3 3
use M3_M2  M3_M2_2806
timestamp 1745462530
transform 1 0 3980 0 1 2275
box -3 -3 3 3
use M3_M2  M3_M2_2807
timestamp 1745462530
transform 1 0 3948 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_2808
timestamp 1745462530
transform 1 0 3948 0 1 1655
box -3 -3 3 3
use M3_M2  M3_M2_2809
timestamp 1745462530
transform 1 0 3908 0 1 2845
box -3 -3 3 3
use M3_M2  M3_M2_2810
timestamp 1745462530
transform 1 0 3900 0 1 2415
box -3 -3 3 3
use M3_M2  M3_M2_2811
timestamp 1745462530
transform 1 0 3900 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_2812
timestamp 1745462530
transform 1 0 3900 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_2813
timestamp 1745462530
transform 1 0 3820 0 1 3125
box -3 -3 3 3
use M3_M2  M3_M2_2814
timestamp 1745462530
transform 1 0 3796 0 1 2845
box -3 -3 3 3
use M3_M2  M3_M2_2815
timestamp 1745462530
transform 1 0 3788 0 1 3125
box -3 -3 3 3
use M3_M2  M3_M2_2816
timestamp 1745462530
transform 1 0 3652 0 1 3125
box -3 -3 3 3
use M3_M2  M3_M2_2817
timestamp 1745462530
transform 1 0 3060 0 1 2415
box -3 -3 3 3
use M3_M2  M3_M2_2818
timestamp 1745462530
transform 1 0 3060 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_2819
timestamp 1745462530
transform 1 0 2668 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_2820
timestamp 1745462530
transform 1 0 2668 0 1 1655
box -3 -3 3 3
use M3_M2  M3_M2_2821
timestamp 1745462530
transform 1 0 2572 0 1 1655
box -3 -3 3 3
use M3_M2  M3_M2_2822
timestamp 1745462530
transform 1 0 2540 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_2823
timestamp 1745462530
transform 1 0 4292 0 1 685
box -3 -3 3 3
use M3_M2  M3_M2_2824
timestamp 1745462530
transform 1 0 4284 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_2825
timestamp 1745462530
transform 1 0 4188 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_2826
timestamp 1745462530
transform 1 0 4180 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_2827
timestamp 1745462530
transform 1 0 4132 0 1 685
box -3 -3 3 3
use M3_M2  M3_M2_2828
timestamp 1745462530
transform 1 0 3844 0 1 685
box -3 -3 3 3
use M3_M2  M3_M2_2829
timestamp 1745462530
transform 1 0 3844 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_2830
timestamp 1745462530
transform 1 0 3764 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_2831
timestamp 1745462530
transform 1 0 3764 0 1 1055
box -3 -3 3 3
use M3_M2  M3_M2_2832
timestamp 1745462530
transform 1 0 3764 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_2833
timestamp 1745462530
transform 1 0 3700 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_2834
timestamp 1745462530
transform 1 0 3700 0 1 1205
box -3 -3 3 3
use M3_M2  M3_M2_2835
timestamp 1745462530
transform 1 0 3700 0 1 605
box -3 -3 3 3
use M3_M2  M3_M2_2836
timestamp 1745462530
transform 1 0 3684 0 1 1205
box -3 -3 3 3
use M3_M2  M3_M2_2837
timestamp 1745462530
transform 1 0 3684 0 1 1055
box -3 -3 3 3
use M3_M2  M3_M2_2838
timestamp 1745462530
transform 1 0 3452 0 1 605
box -3 -3 3 3
use M3_M2  M3_M2_2839
timestamp 1745462530
transform 1 0 2604 0 1 1435
box -3 -3 3 3
use M3_M2  M3_M2_2840
timestamp 1745462530
transform 1 0 2572 0 1 1435
box -3 -3 3 3
use M3_M2  M3_M2_2841
timestamp 1745462530
transform 1 0 2564 0 1 1215
box -3 -3 3 3
use M3_M2  M3_M2_2842
timestamp 1745462530
transform 1 0 2468 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_2843
timestamp 1745462530
transform 1 0 2460 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_2844
timestamp 1745462530
transform 1 0 2356 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_2845
timestamp 1745462530
transform 1 0 2356 0 1 285
box -3 -3 3 3
use M3_M2  M3_M2_2846
timestamp 1745462530
transform 1 0 2356 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_2847
timestamp 1745462530
transform 1 0 2340 0 1 775
box -3 -3 3 3
use M3_M2  M3_M2_2848
timestamp 1745462530
transform 1 0 2308 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_2849
timestamp 1745462530
transform 1 0 2308 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_2850
timestamp 1745462530
transform 1 0 2244 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_2851
timestamp 1745462530
transform 1 0 2156 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_2852
timestamp 1745462530
transform 1 0 2156 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_2853
timestamp 1745462530
transform 1 0 2156 0 1 775
box -3 -3 3 3
use M3_M2  M3_M2_2854
timestamp 1745462530
transform 1 0 2076 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_2855
timestamp 1745462530
transform 1 0 2060 0 1 775
box -3 -3 3 3
use M3_M2  M3_M2_2856
timestamp 1745462530
transform 1 0 1988 0 1 285
box -3 -3 3 3
use M3_M2  M3_M2_2857
timestamp 1745462530
transform 1 0 1972 0 1 775
box -3 -3 3 3
use M3_M2  M3_M2_2858
timestamp 1745462530
transform 1 0 1644 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_2859
timestamp 1745462530
transform 1 0 1572 0 1 285
box -3 -3 3 3
use M3_M2  M3_M2_2860
timestamp 1745462530
transform 1 0 1044 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_2861
timestamp 1745462530
transform 1 0 1044 0 1 285
box -3 -3 3 3
use M3_M2  M3_M2_2862
timestamp 1745462530
transform 1 0 892 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_2863
timestamp 1745462530
transform 1 0 804 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_2864
timestamp 1745462530
transform 1 0 772 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_2865
timestamp 1745462530
transform 1 0 764 0 1 1775
box -3 -3 3 3
use M3_M2  M3_M2_2866
timestamp 1745462530
transform 1 0 764 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_2867
timestamp 1745462530
transform 1 0 356 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_2868
timestamp 1745462530
transform 1 0 308 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_2869
timestamp 1745462530
transform 1 0 284 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_2870
timestamp 1745462530
transform 1 0 252 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_2871
timestamp 1745462530
transform 1 0 252 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_2872
timestamp 1745462530
transform 1 0 212 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_2873
timestamp 1745462530
transform 1 0 116 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_2874
timestamp 1745462530
transform 1 0 116 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_2875
timestamp 1745462530
transform 1 0 100 0 1 375
box -3 -3 3 3
use M3_M2  M3_M2_2876
timestamp 1745462530
transform 1 0 76 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_2877
timestamp 1745462530
transform 1 0 2844 0 1 2925
box -3 -3 3 3
use M3_M2  M3_M2_2878
timestamp 1745462530
transform 1 0 2836 0 1 2685
box -3 -3 3 3
use M3_M2  M3_M2_2879
timestamp 1745462530
transform 1 0 2740 0 1 2675
box -3 -3 3 3
use M3_M2  M3_M2_2880
timestamp 1745462530
transform 1 0 2660 0 1 2925
box -3 -3 3 3
use M3_M2  M3_M2_2881
timestamp 1745462530
transform 1 0 2108 0 1 1975
box -3 -3 3 3
use M3_M2  M3_M2_2882
timestamp 1745462530
transform 1 0 1980 0 1 1975
box -3 -3 3 3
use M3_M2  M3_M2_2883
timestamp 1745462530
transform 1 0 1916 0 1 2675
box -3 -3 3 3
use M3_M2  M3_M2_2884
timestamp 1745462530
transform 1 0 1908 0 1 1975
box -3 -3 3 3
use M3_M2  M3_M2_2885
timestamp 1745462530
transform 1 0 1900 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_2886
timestamp 1745462530
transform 1 0 1892 0 1 2675
box -3 -3 3 3
use M3_M2  M3_M2_2887
timestamp 1745462530
transform 1 0 1884 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_2888
timestamp 1745462530
transform 1 0 1884 0 1 1975
box -3 -3 3 3
use M3_M2  M3_M2_2889
timestamp 1745462530
transform 1 0 1876 0 1 2755
box -3 -3 3 3
use M3_M2  M3_M2_2890
timestamp 1745462530
transform 1 0 1836 0 1 2565
box -3 -3 3 3
use M3_M2  M3_M2_2891
timestamp 1745462530
transform 1 0 1836 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_2892
timestamp 1745462530
transform 1 0 1812 0 1 2845
box -3 -3 3 3
use M3_M2  M3_M2_2893
timestamp 1745462530
transform 1 0 1780 0 1 2895
box -3 -3 3 3
use M3_M2  M3_M2_2894
timestamp 1745462530
transform 1 0 1780 0 1 2845
box -3 -3 3 3
use M3_M2  M3_M2_2895
timestamp 1745462530
transform 1 0 1772 0 1 2755
box -3 -3 3 3
use M3_M2  M3_M2_2896
timestamp 1745462530
transform 1 0 1716 0 1 2565
box -3 -3 3 3
use M3_M2  M3_M2_2897
timestamp 1745462530
transform 1 0 1012 0 1 2965
box -3 -3 3 3
use M3_M2  M3_M2_2898
timestamp 1745462530
transform 1 0 1012 0 1 2895
box -3 -3 3 3
use M3_M2  M3_M2_2899
timestamp 1745462530
transform 1 0 756 0 1 2965
box -3 -3 3 3
use M3_M2  M3_M2_2900
timestamp 1745462530
transform 1 0 652 0 1 2965
box -3 -3 3 3
use M3_M2  M3_M2_2901
timestamp 1745462530
transform 1 0 444 0 1 2965
box -3 -3 3 3
use M3_M2  M3_M2_2902
timestamp 1745462530
transform 1 0 4260 0 1 2125
box -3 -3 3 3
use M3_M2  M3_M2_2903
timestamp 1745462530
transform 1 0 4260 0 1 1855
box -3 -3 3 3
use M3_M2  M3_M2_2904
timestamp 1745462530
transform 1 0 4100 0 1 2125
box -3 -3 3 3
use M3_M2  M3_M2_2905
timestamp 1745462530
transform 1 0 4076 0 1 1855
box -3 -3 3 3
use M3_M2  M3_M2_2906
timestamp 1745462530
transform 1 0 4044 0 1 2125
box -3 -3 3 3
use M3_M2  M3_M2_2907
timestamp 1745462530
transform 1 0 4044 0 1 2085
box -3 -3 3 3
use M3_M2  M3_M2_2908
timestamp 1745462530
transform 1 0 3612 0 1 2085
box -3 -3 3 3
use M3_M2  M3_M2_2909
timestamp 1745462530
transform 1 0 3604 0 1 2155
box -3 -3 3 3
use M3_M2  M3_M2_2910
timestamp 1745462530
transform 1 0 3484 0 1 2155
box -3 -3 3 3
use M3_M2  M3_M2_2911
timestamp 1745462530
transform 1 0 3484 0 1 2055
box -3 -3 3 3
use M3_M2  M3_M2_2912
timestamp 1745462530
transform 1 0 3460 0 1 2605
box -3 -3 3 3
use M3_M2  M3_M2_2913
timestamp 1745462530
transform 1 0 3452 0 1 2845
box -3 -3 3 3
use M3_M2  M3_M2_2914
timestamp 1745462530
transform 1 0 3444 0 1 2605
box -3 -3 3 3
use M3_M2  M3_M2_2915
timestamp 1745462530
transform 1 0 3436 0 1 2155
box -3 -3 3 3
use M3_M2  M3_M2_2916
timestamp 1745462530
transform 1 0 3388 0 1 2605
box -3 -3 3 3
use M3_M2  M3_M2_2917
timestamp 1745462530
transform 1 0 3372 0 1 2845
box -3 -3 3 3
use M3_M2  M3_M2_2918
timestamp 1745462530
transform 1 0 3372 0 1 2065
box -3 -3 3 3
use M3_M2  M3_M2_2919
timestamp 1745462530
transform 1 0 3364 0 1 3015
box -3 -3 3 3
use M3_M2  M3_M2_2920
timestamp 1745462530
transform 1 0 3252 0 1 3015
box -3 -3 3 3
use M3_M2  M3_M2_2921
timestamp 1745462530
transform 1 0 2676 0 1 2175
box -3 -3 3 3
use M3_M2  M3_M2_2922
timestamp 1745462530
transform 1 0 2676 0 1 2065
box -3 -3 3 3
use M3_M2  M3_M2_2923
timestamp 1745462530
transform 1 0 2500 0 1 2065
box -3 -3 3 3
use M3_M2  M3_M2_2924
timestamp 1745462530
transform 1 0 2492 0 1 2175
box -3 -3 3 3
use M3_M2  M3_M2_2925
timestamp 1745462530
transform 1 0 2276 0 1 2065
box -3 -3 3 3
use M3_M2  M3_M2_2926
timestamp 1745462530
transform 1 0 3988 0 1 645
box -3 -3 3 3
use M3_M2  M3_M2_2927
timestamp 1745462530
transform 1 0 3988 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_2928
timestamp 1745462530
transform 1 0 3956 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_2929
timestamp 1745462530
transform 1 0 3908 0 1 1015
box -3 -3 3 3
use M3_M2  M3_M2_2930
timestamp 1745462530
transform 1 0 3860 0 1 725
box -3 -3 3 3
use M3_M2  M3_M2_2931
timestamp 1745462530
transform 1 0 3860 0 1 645
box -3 -3 3 3
use M3_M2  M3_M2_2932
timestamp 1745462530
transform 1 0 3476 0 1 1015
box -3 -3 3 3
use M3_M2  M3_M2_2933
timestamp 1745462530
transform 1 0 3476 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_2934
timestamp 1745462530
transform 1 0 3468 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_2935
timestamp 1745462530
transform 1 0 3468 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_2936
timestamp 1745462530
transform 1 0 3436 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_2937
timestamp 1745462530
transform 1 0 3420 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_2938
timestamp 1745462530
transform 1 0 3412 0 1 455
box -3 -3 3 3
use M3_M2  M3_M2_2939
timestamp 1745462530
transform 1 0 3228 0 1 455
box -3 -3 3 3
use M3_M2  M3_M2_2940
timestamp 1745462530
transform 1 0 2668 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_2941
timestamp 1745462530
transform 1 0 2660 0 1 455
box -3 -3 3 3
use M3_M2  M3_M2_2942
timestamp 1745462530
transform 1 0 2612 0 1 865
box -3 -3 3 3
use M3_M2  M3_M2_2943
timestamp 1745462530
transform 1 0 2596 0 1 445
box -3 -3 3 3
use M3_M2  M3_M2_2944
timestamp 1745462530
transform 1 0 2556 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_2945
timestamp 1745462530
transform 1 0 2532 0 1 865
box -3 -3 3 3
use M3_M2  M3_M2_2946
timestamp 1745462530
transform 1 0 2340 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_2947
timestamp 1745462530
transform 1 0 2332 0 1 865
box -3 -3 3 3
use M3_M2  M3_M2_2948
timestamp 1745462530
transform 1 0 2204 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_2949
timestamp 1745462530
transform 1 0 2196 0 1 1435
box -3 -3 3 3
use M3_M2  M3_M2_2950
timestamp 1745462530
transform 1 0 2124 0 1 365
box -3 -3 3 3
use M3_M2  M3_M2_2951
timestamp 1745462530
transform 1 0 2108 0 1 1435
box -3 -3 3 3
use M3_M2  M3_M2_2952
timestamp 1745462530
transform 1 0 2108 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_2953
timestamp 1745462530
transform 1 0 2100 0 1 365
box -3 -3 3 3
use M3_M2  M3_M2_2954
timestamp 1745462530
transform 1 0 1380 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_2955
timestamp 1745462530
transform 1 0 1332 0 1 1085
box -3 -3 3 3
use M3_M2  M3_M2_2956
timestamp 1745462530
transform 1 0 1316 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_2957
timestamp 1745462530
transform 1 0 1308 0 1 1085
box -3 -3 3 3
use M3_M2  M3_M2_2958
timestamp 1745462530
transform 1 0 1292 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_2959
timestamp 1745462530
transform 1 0 1244 0 1 365
box -3 -3 3 3
use M3_M2  M3_M2_2960
timestamp 1745462530
transform 1 0 1212 0 1 495
box -3 -3 3 3
use M3_M2  M3_M2_2961
timestamp 1745462530
transform 1 0 1204 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_2962
timestamp 1745462530
transform 1 0 1196 0 1 495
box -3 -3 3 3
use M3_M2  M3_M2_2963
timestamp 1745462530
transform 1 0 1196 0 1 365
box -3 -3 3 3
use M3_M2  M3_M2_2964
timestamp 1745462530
transform 1 0 1020 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_2965
timestamp 1745462530
transform 1 0 1012 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_2966
timestamp 1745462530
transform 1 0 980 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_2967
timestamp 1745462530
transform 1 0 924 0 1 1495
box -3 -3 3 3
use M3_M2  M3_M2_2968
timestamp 1745462530
transform 1 0 844 0 1 605
box -3 -3 3 3
use M3_M2  M3_M2_2969
timestamp 1745462530
transform 1 0 812 0 1 2525
box -3 -3 3 3
use M3_M2  M3_M2_2970
timestamp 1745462530
transform 1 0 788 0 1 1495
box -3 -3 3 3
use M3_M2  M3_M2_2971
timestamp 1745462530
transform 1 0 652 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_2972
timestamp 1745462530
transform 1 0 132 0 1 2055
box -3 -3 3 3
use M3_M2  M3_M2_2973
timestamp 1745462530
transform 1 0 124 0 1 605
box -3 -3 3 3
use M3_M2  M3_M2_2974
timestamp 1745462530
transform 1 0 92 0 1 2555
box -3 -3 3 3
use M3_M2  M3_M2_2975
timestamp 1745462530
transform 1 0 92 0 1 2525
box -3 -3 3 3
use M3_M2  M3_M2_2976
timestamp 1745462530
transform 1 0 92 0 1 2415
box -3 -3 3 3
use M3_M2  M3_M2_2977
timestamp 1745462530
transform 1 0 92 0 1 2385
box -3 -3 3 3
use M3_M2  M3_M2_2978
timestamp 1745462530
transform 1 0 92 0 1 2055
box -3 -3 3 3
use M3_M2  M3_M2_2979
timestamp 1745462530
transform 1 0 76 0 1 1495
box -3 -3 3 3
use M3_M2  M3_M2_2980
timestamp 1745462530
transform 1 0 1468 0 1 3225
box -3 -3 3 3
use M3_M2  M3_M2_2981
timestamp 1745462530
transform 1 0 1404 0 1 3225
box -3 -3 3 3
use M3_M2  M3_M2_2982
timestamp 1745462530
transform 1 0 1148 0 1 3225
box -3 -3 3 3
use M3_M2  M3_M2_2983
timestamp 1745462530
transform 1 0 1148 0 1 3195
box -3 -3 3 3
use M3_M2  M3_M2_2984
timestamp 1745462530
transform 1 0 1108 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_2985
timestamp 1745462530
transform 1 0 1084 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_2986
timestamp 1745462530
transform 1 0 1084 0 1 2715
box -3 -3 3 3
use M3_M2  M3_M2_2987
timestamp 1745462530
transform 1 0 1052 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_2988
timestamp 1745462530
transform 1 0 1052 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_2989
timestamp 1745462530
transform 1 0 1052 0 1 2525
box -3 -3 3 3
use M3_M2  M3_M2_2990
timestamp 1745462530
transform 1 0 1004 0 1 2165
box -3 -3 3 3
use M3_M2  M3_M2_2991
timestamp 1745462530
transform 1 0 996 0 1 3195
box -3 -3 3 3
use M3_M2  M3_M2_2992
timestamp 1745462530
transform 1 0 988 0 1 2525
box -3 -3 3 3
use M3_M2  M3_M2_2993
timestamp 1745462530
transform 1 0 980 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_2994
timestamp 1745462530
transform 1 0 980 0 1 2715
box -3 -3 3 3
use M3_M2  M3_M2_2995
timestamp 1745462530
transform 1 0 980 0 1 2165
box -3 -3 3 3
use M3_M2  M3_M2_2996
timestamp 1745462530
transform 1 0 980 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_2997
timestamp 1745462530
transform 1 0 868 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_2998
timestamp 1745462530
transform 1 0 852 0 1 3195
box -3 -3 3 3
use M3_M2  M3_M2_2999
timestamp 1745462530
transform 1 0 2364 0 1 2835
box -3 -3 3 3
use M3_M2  M3_M2_3000
timestamp 1745462530
transform 1 0 2308 0 1 3015
box -3 -3 3 3
use M3_M2  M3_M2_3001
timestamp 1745462530
transform 1 0 2292 0 1 2835
box -3 -3 3 3
use M3_M2  M3_M2_3002
timestamp 1745462530
transform 1 0 2268 0 1 3015
box -3 -3 3 3
use M3_M2  M3_M2_3003
timestamp 1745462530
transform 1 0 2260 0 1 3085
box -3 -3 3 3
use M3_M2  M3_M2_3004
timestamp 1745462530
transform 1 0 2196 0 1 2775
box -3 -3 3 3
use M3_M2  M3_M2_3005
timestamp 1745462530
transform 1 0 2132 0 1 2815
box -3 -3 3 3
use M3_M2  M3_M2_3006
timestamp 1745462530
transform 1 0 2132 0 1 2775
box -3 -3 3 3
use M3_M2  M3_M2_3007
timestamp 1745462530
transform 1 0 2100 0 1 2775
box -3 -3 3 3
use M3_M2  M3_M2_3008
timestamp 1745462530
transform 1 0 2012 0 1 3085
box -3 -3 3 3
use M3_M2  M3_M2_3009
timestamp 1745462530
transform 1 0 2012 0 1 2815
box -3 -3 3 3
use M3_M2  M3_M2_3010
timestamp 1745462530
transform 1 0 2012 0 1 2775
box -3 -3 3 3
use M3_M2  M3_M2_3011
timestamp 1745462530
transform 1 0 1996 0 1 2775
box -3 -3 3 3
use M3_M2  M3_M2_3012
timestamp 1745462530
transform 1 0 1044 0 1 3065
box -3 -3 3 3
use M3_M2  M3_M2_3013
timestamp 1745462530
transform 1 0 1036 0 1 3715
box -3 -3 3 3
use M3_M2  M3_M2_3014
timestamp 1745462530
transform 1 0 1028 0 1 3315
box -3 -3 3 3
use M3_M2  M3_M2_3015
timestamp 1745462530
transform 1 0 900 0 1 3715
box -3 -3 3 3
use M3_M2  M3_M2_3016
timestamp 1745462530
transform 1 0 900 0 1 3565
box -3 -3 3 3
use M3_M2  M3_M2_3017
timestamp 1745462530
transform 1 0 764 0 1 3555
box -3 -3 3 3
use M3_M2  M3_M2_3018
timestamp 1745462530
transform 1 0 732 0 1 3315
box -3 -3 3 3
use M3_M2  M3_M2_3019
timestamp 1745462530
transform 1 0 692 0 1 3555
box -3 -3 3 3
use M3_M2  M3_M2_3020
timestamp 1745462530
transform 1 0 1180 0 1 3155
box -3 -3 3 3
use M3_M2  M3_M2_3021
timestamp 1745462530
transform 1 0 964 0 1 3175
box -3 -3 3 3
use M3_M2  M3_M2_3022
timestamp 1745462530
transform 1 0 964 0 1 3155
box -3 -3 3 3
use M3_M2  M3_M2_3023
timestamp 1745462530
transform 1 0 692 0 1 3175
box -3 -3 3 3
use M3_M2  M3_M2_3024
timestamp 1745462530
transform 1 0 620 0 1 3175
box -3 -3 3 3
use M3_M2  M3_M2_3025
timestamp 1745462530
transform 1 0 612 0 1 3305
box -3 -3 3 3
use M3_M2  M3_M2_3026
timestamp 1745462530
transform 1 0 404 0 1 3745
box -3 -3 3 3
use M3_M2  M3_M2_3027
timestamp 1745462530
transform 1 0 356 0 1 3305
box -3 -3 3 3
use M3_M2  M3_M2_3028
timestamp 1745462530
transform 1 0 292 0 1 3745
box -3 -3 3 3
use M3_M2  M3_M2_3029
timestamp 1745462530
transform 1 0 268 0 1 3305
box -3 -3 3 3
use M3_M2  M3_M2_3030
timestamp 1745462530
transform 1 0 156 0 1 3745
box -3 -3 3 3
use M3_M2  M3_M2_3031
timestamp 1745462530
transform 1 0 148 0 1 3345
box -3 -3 3 3
use M3_M2  M3_M2_3032
timestamp 1745462530
transform 1 0 148 0 1 3305
box -3 -3 3 3
use M3_M2  M3_M2_3033
timestamp 1745462530
transform 1 0 92 0 1 3745
box -3 -3 3 3
use M3_M2  M3_M2_3034
timestamp 1745462530
transform 1 0 92 0 1 3345
box -3 -3 3 3
use M3_M2  M3_M2_3035
timestamp 1745462530
transform 1 0 2212 0 1 1535
box -3 -3 3 3
use M3_M2  M3_M2_3036
timestamp 1745462530
transform 1 0 2148 0 1 1535
box -3 -3 3 3
use M3_M2  M3_M2_3037
timestamp 1745462530
transform 1 0 2060 0 1 1655
box -3 -3 3 3
use M3_M2  M3_M2_3038
timestamp 1745462530
transform 1 0 2028 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_3039
timestamp 1745462530
transform 1 0 2028 0 1 1655
box -3 -3 3 3
use M3_M2  M3_M2_3040
timestamp 1745462530
transform 1 0 1988 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_3041
timestamp 1745462530
transform 1 0 2132 0 1 1465
box -3 -3 3 3
use M3_M2  M3_M2_3042
timestamp 1745462530
transform 1 0 2052 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_3043
timestamp 1745462530
transform 1 0 2052 0 1 1465
box -3 -3 3 3
use M3_M2  M3_M2_3044
timestamp 1745462530
transform 1 0 1956 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_3045
timestamp 1745462530
transform 1 0 4372 0 1 3905
box -3 -3 3 3
use M3_M2  M3_M2_3046
timestamp 1745462530
transform 1 0 3964 0 1 3665
box -3 -3 3 3
use M3_M2  M3_M2_3047
timestamp 1745462530
transform 1 0 3964 0 1 3565
box -3 -3 3 3
use M3_M2  M3_M2_3048
timestamp 1745462530
transform 1 0 3940 0 1 3665
box -3 -3 3 3
use M3_M2  M3_M2_3049
timestamp 1745462530
transform 1 0 3932 0 1 3905
box -3 -3 3 3
use M3_M2  M3_M2_3050
timestamp 1745462530
transform 1 0 3916 0 1 3565
box -3 -3 3 3
use M3_M2  M3_M2_3051
timestamp 1745462530
transform 1 0 1860 0 1 3265
box -3 -3 3 3
use M3_M2  M3_M2_3052
timestamp 1745462530
transform 1 0 1780 0 1 3315
box -3 -3 3 3
use M3_M2  M3_M2_3053
timestamp 1745462530
transform 1 0 1780 0 1 3265
box -3 -3 3 3
use M3_M2  M3_M2_3054
timestamp 1745462530
transform 1 0 1740 0 1 3735
box -3 -3 3 3
use M3_M2  M3_M2_3055
timestamp 1745462530
transform 1 0 1740 0 1 3645
box -3 -3 3 3
use M3_M2  M3_M2_3056
timestamp 1745462530
transform 1 0 1716 0 1 3645
box -3 -3 3 3
use M3_M2  M3_M2_3057
timestamp 1745462530
transform 1 0 1716 0 1 3625
box -3 -3 3 3
use M3_M2  M3_M2_3058
timestamp 1745462530
transform 1 0 1676 0 1 3985
box -3 -3 3 3
use M3_M2  M3_M2_3059
timestamp 1745462530
transform 1 0 1668 0 1 3365
box -3 -3 3 3
use M3_M2  M3_M2_3060
timestamp 1745462530
transform 1 0 1668 0 1 3315
box -3 -3 3 3
use M3_M2  M3_M2_3061
timestamp 1745462530
transform 1 0 1620 0 1 3985
box -3 -3 3 3
use M3_M2  M3_M2_3062
timestamp 1745462530
transform 1 0 1620 0 1 3835
box -3 -3 3 3
use M3_M2  M3_M2_3063
timestamp 1745462530
transform 1 0 1524 0 1 3835
box -3 -3 3 3
use M3_M2  M3_M2_3064
timestamp 1745462530
transform 1 0 1524 0 1 3605
box -3 -3 3 3
use M3_M2  M3_M2_3065
timestamp 1745462530
transform 1 0 1524 0 1 3365
box -3 -3 3 3
use M3_M2  M3_M2_3066
timestamp 1745462530
transform 1 0 1516 0 1 3735
box -3 -3 3 3
use M3_M2  M3_M2_3067
timestamp 1745462530
transform 1 0 1572 0 1 2695
box -3 -3 3 3
use M3_M2  M3_M2_3068
timestamp 1745462530
transform 1 0 1556 0 1 2185
box -3 -3 3 3
use M3_M2  M3_M2_3069
timestamp 1745462530
transform 1 0 1548 0 1 2065
box -3 -3 3 3
use M3_M2  M3_M2_3070
timestamp 1745462530
transform 1 0 1540 0 1 2695
box -3 -3 3 3
use M3_M2  M3_M2_3071
timestamp 1745462530
transform 1 0 1524 0 1 2185
box -3 -3 3 3
use M3_M2  M3_M2_3072
timestamp 1745462530
transform 1 0 1524 0 1 2065
box -3 -3 3 3
use M3_M2  M3_M2_3073
timestamp 1745462530
transform 1 0 1380 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_3074
timestamp 1745462530
transform 1 0 1364 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_3075
timestamp 1745462530
transform 1 0 1348 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_3076
timestamp 1745462530
transform 1 0 1348 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_3077
timestamp 1745462530
transform 1 0 1316 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_3078
timestamp 1745462530
transform 1 0 1244 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_3079
timestamp 1745462530
transform 1 0 1244 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_3080
timestamp 1745462530
transform 1 0 924 0 1 2755
box -3 -3 3 3
use M3_M2  M3_M2_3081
timestamp 1745462530
transform 1 0 580 0 1 2755
box -3 -3 3 3
use M3_M2  M3_M2_3082
timestamp 1745462530
transform 1 0 484 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_3083
timestamp 1745462530
transform 1 0 276 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_3084
timestamp 1745462530
transform 1 0 276 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_3085
timestamp 1745462530
transform 1 0 252 0 1 2755
box -3 -3 3 3
use M3_M2  M3_M2_3086
timestamp 1745462530
transform 1 0 252 0 1 2365
box -3 -3 3 3
use M3_M2  M3_M2_3087
timestamp 1745462530
transform 1 0 220 0 1 2755
box -3 -3 3 3
use M3_M2  M3_M2_3088
timestamp 1745462530
transform 1 0 212 0 1 2365
box -3 -3 3 3
use M3_M2  M3_M2_3089
timestamp 1745462530
transform 1 0 204 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_3090
timestamp 1745462530
transform 1 0 172 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_3091
timestamp 1745462530
transform 1 0 172 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_3092
timestamp 1745462530
transform 1 0 1348 0 1 1295
box -3 -3 3 3
use M3_M2  M3_M2_3093
timestamp 1745462530
transform 1 0 1348 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_3094
timestamp 1745462530
transform 1 0 1348 0 1 295
box -3 -3 3 3
use M3_M2  M3_M2_3095
timestamp 1745462530
transform 1 0 1324 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_3096
timestamp 1745462530
transform 1 0 1324 0 1 865
box -3 -3 3 3
use M3_M2  M3_M2_3097
timestamp 1745462530
transform 1 0 1316 0 1 295
box -3 -3 3 3
use M3_M2  M3_M2_3098
timestamp 1745462530
transform 1 0 1292 0 1 1295
box -3 -3 3 3
use M3_M2  M3_M2_3099
timestamp 1745462530
transform 1 0 1268 0 1 295
box -3 -3 3 3
use M3_M2  M3_M2_3100
timestamp 1745462530
transform 1 0 1260 0 1 865
box -3 -3 3 3
use M3_M2  M3_M2_3101
timestamp 1745462530
transform 1 0 1084 0 1 495
box -3 -3 3 3
use M3_M2  M3_M2_3102
timestamp 1745462530
transform 1 0 1084 0 1 295
box -3 -3 3 3
use M3_M2  M3_M2_3103
timestamp 1745462530
transform 1 0 1028 0 1 495
box -3 -3 3 3
use M3_M2  M3_M2_3104
timestamp 1745462530
transform 1 0 844 0 1 1295
box -3 -3 3 3
use M3_M2  M3_M2_3105
timestamp 1745462530
transform 1 0 820 0 1 295
box -3 -3 3 3
use M3_M2  M3_M2_3106
timestamp 1745462530
transform 1 0 612 0 1 295
box -3 -3 3 3
use M3_M2  M3_M2_3107
timestamp 1745462530
transform 1 0 612 0 1 245
box -3 -3 3 3
use M3_M2  M3_M2_3108
timestamp 1745462530
transform 1 0 476 0 1 245
box -3 -3 3 3
use M3_M2  M3_M2_3109
timestamp 1745462530
transform 1 0 428 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_3110
timestamp 1745462530
transform 1 0 412 0 1 1295
box -3 -3 3 3
use M3_M2  M3_M2_3111
timestamp 1745462530
transform 1 0 396 0 1 245
box -3 -3 3 3
use M3_M2  M3_M2_3112
timestamp 1745462530
transform 1 0 372 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_3113
timestamp 1745462530
transform 1 0 3172 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_3114
timestamp 1745462530
transform 1 0 3036 0 1 205
box -3 -3 3 3
use M3_M2  M3_M2_3115
timestamp 1745462530
transform 1 0 2796 0 1 465
box -3 -3 3 3
use M3_M2  M3_M2_3116
timestamp 1745462530
transform 1 0 2796 0 1 205
box -3 -3 3 3
use M3_M2  M3_M2_3117
timestamp 1745462530
transform 1 0 2772 0 1 465
box -3 -3 3 3
use M3_M2  M3_M2_3118
timestamp 1745462530
transform 1 0 2740 0 1 205
box -3 -3 3 3
use M3_M2  M3_M2_3119
timestamp 1745462530
transform 1 0 2724 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_3120
timestamp 1745462530
transform 1 0 2676 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_3121
timestamp 1745462530
transform 1 0 2676 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_3122
timestamp 1745462530
transform 1 0 2652 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_3123
timestamp 1745462530
transform 1 0 2652 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_3124
timestamp 1745462530
transform 1 0 2636 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_3125
timestamp 1745462530
transform 1 0 2612 0 1 205
box -3 -3 3 3
use M3_M2  M3_M2_3126
timestamp 1745462530
transform 1 0 2220 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_3127
timestamp 1745462530
transform 1 0 2180 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_3128
timestamp 1745462530
transform 1 0 2180 0 1 1405
box -3 -3 3 3
use M3_M2  M3_M2_3129
timestamp 1745462530
transform 1 0 2036 0 1 1285
box -3 -3 3 3
use M3_M2  M3_M2_3130
timestamp 1745462530
transform 1 0 2028 0 1 1405
box -3 -3 3 3
use M3_M2  M3_M2_3131
timestamp 1745462530
transform 1 0 1956 0 1 1285
box -3 -3 3 3
use M3_M2  M3_M2_3132
timestamp 1745462530
transform 1 0 1956 0 1 1085
box -3 -3 3 3
use M3_M2  M3_M2_3133
timestamp 1745462530
transform 1 0 1412 0 1 1085
box -3 -3 3 3
use M3_M2  M3_M2_3134
timestamp 1745462530
transform 1 0 4380 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_3135
timestamp 1745462530
transform 1 0 4380 0 1 975
box -3 -3 3 3
use M3_M2  M3_M2_3136
timestamp 1745462530
transform 1 0 4324 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_3137
timestamp 1745462530
transform 1 0 4308 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_3138
timestamp 1745462530
transform 1 0 4252 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_3139
timestamp 1745462530
transform 1 0 4228 0 1 975
box -3 -3 3 3
use M3_M2  M3_M2_3140
timestamp 1745462530
transform 1 0 4228 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_3141
timestamp 1745462530
transform 1 0 4220 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_3142
timestamp 1745462530
transform 1 0 4204 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_3143
timestamp 1745462530
transform 1 0 4156 0 1 975
box -3 -3 3 3
use M3_M2  M3_M2_3144
timestamp 1745462530
transform 1 0 4148 0 1 1085
box -3 -3 3 3
use M3_M2  M3_M2_3145
timestamp 1745462530
transform 1 0 3780 0 1 2005
box -3 -3 3 3
use M3_M2  M3_M2_3146
timestamp 1745462530
transform 1 0 3732 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_3147
timestamp 1745462530
transform 1 0 3716 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_3148
timestamp 1745462530
transform 1 0 3700 0 1 2005
box -3 -3 3 3
use M3_M2  M3_M2_3149
timestamp 1745462530
transform 1 0 3700 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_3150
timestamp 1745462530
transform 1 0 3684 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_3151
timestamp 1745462530
transform 1 0 3660 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_3152
timestamp 1745462530
transform 1 0 3660 0 1 1085
box -3 -3 3 3
use M3_M2  M3_M2_3153
timestamp 1745462530
transform 1 0 3628 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_3154
timestamp 1745462530
transform 1 0 3612 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_3155
timestamp 1745462530
transform 1 0 3540 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_3156
timestamp 1745462530
transform 1 0 2652 0 1 2005
box -3 -3 3 3
use M3_M2  M3_M2_3157
timestamp 1745462530
transform 1 0 3700 0 1 2945
box -3 -3 3 3
use M3_M2  M3_M2_3158
timestamp 1745462530
transform 1 0 3628 0 1 2845
box -3 -3 3 3
use M3_M2  M3_M2_3159
timestamp 1745462530
transform 1 0 3532 0 1 2935
box -3 -3 3 3
use M3_M2  M3_M2_3160
timestamp 1745462530
transform 1 0 3508 0 1 2935
box -3 -3 3 3
use M3_M2  M3_M2_3161
timestamp 1745462530
transform 1 0 3500 0 1 2845
box -3 -3 3 3
use M3_M2  M3_M2_3162
timestamp 1745462530
transform 1 0 3500 0 1 2715
box -3 -3 3 3
use M3_M2  M3_M2_3163
timestamp 1745462530
transform 1 0 3468 0 1 2935
box -3 -3 3 3
use M3_M2  M3_M2_3164
timestamp 1745462530
transform 1 0 2868 0 1 2715
box -3 -3 3 3
use M3_M2  M3_M2_3165
timestamp 1745462530
transform 1 0 2868 0 1 2605
box -3 -3 3 3
use M3_M2  M3_M2_3166
timestamp 1745462530
transform 1 0 2860 0 1 2215
box -3 -3 3 3
use M3_M2  M3_M2_3167
timestamp 1745462530
transform 1 0 2828 0 1 2085
box -3 -3 3 3
use M3_M2  M3_M2_3168
timestamp 1745462530
transform 1 0 2812 0 1 2215
box -3 -3 3 3
use M3_M2  M3_M2_3169
timestamp 1745462530
transform 1 0 2676 0 1 2705
box -3 -3 3 3
use M3_M2  M3_M2_3170
timestamp 1745462530
transform 1 0 2676 0 1 2605
box -3 -3 3 3
use M3_M2  M3_M2_3171
timestamp 1745462530
transform 1 0 2612 0 1 2705
box -3 -3 3 3
use M3_M2  M3_M2_3172
timestamp 1745462530
transform 1 0 2596 0 1 2085
box -3 -3 3 3
use M3_M2  M3_M2_3173
timestamp 1745462530
transform 1 0 2596 0 1 2005
box -3 -3 3 3
use M3_M2  M3_M2_3174
timestamp 1745462530
transform 1 0 2580 0 1 2005
box -3 -3 3 3
use M3_M2  M3_M2_3175
timestamp 1745462530
transform 1 0 1532 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_3176
timestamp 1745462530
transform 1 0 1292 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_3177
timestamp 1745462530
transform 1 0 2556 0 1 2005
box -3 -3 3 3
use M3_M2  M3_M2_3178
timestamp 1745462530
transform 1 0 2220 0 1 2005
box -3 -3 3 3
use M3_M2  M3_M2_3179
timestamp 1745462530
transform 1 0 1236 0 1 2575
box -3 -3 3 3
use M3_M2  M3_M2_3180
timestamp 1745462530
transform 1 0 1228 0 1 2265
box -3 -3 3 3
use M3_M2  M3_M2_3181
timestamp 1745462530
transform 1 0 1180 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_3182
timestamp 1745462530
transform 1 0 1180 0 1 2265
box -3 -3 3 3
use M3_M2  M3_M2_3183
timestamp 1745462530
transform 1 0 1148 0 1 2575
box -3 -3 3 3
use M3_M2  M3_M2_3184
timestamp 1745462530
transform 1 0 1148 0 1 2365
box -3 -3 3 3
use M3_M2  M3_M2_3185
timestamp 1745462530
transform 1 0 1108 0 1 2365
box -3 -3 3 3
use M3_M2  M3_M2_3186
timestamp 1745462530
transform 1 0 1108 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_3187
timestamp 1745462530
transform 1 0 1204 0 1 2285
box -3 -3 3 3
use M3_M2  M3_M2_3188
timestamp 1745462530
transform 1 0 1188 0 1 2465
box -3 -3 3 3
use M3_M2  M3_M2_3189
timestamp 1745462530
transform 1 0 1124 0 1 1645
box -3 -3 3 3
use M3_M2  M3_M2_3190
timestamp 1745462530
transform 1 0 1108 0 1 2465
box -3 -3 3 3
use M3_M2  M3_M2_3191
timestamp 1745462530
transform 1 0 1092 0 1 2285
box -3 -3 3 3
use M3_M2  M3_M2_3192
timestamp 1745462530
transform 1 0 956 0 1 2845
box -3 -3 3 3
use M3_M2  M3_M2_3193
timestamp 1745462530
transform 1 0 860 0 1 2765
box -3 -3 3 3
use M3_M2  M3_M2_3194
timestamp 1745462530
transform 1 0 860 0 1 2715
box -3 -3 3 3
use M3_M2  M3_M2_3195
timestamp 1745462530
transform 1 0 844 0 1 2845
box -3 -3 3 3
use M3_M2  M3_M2_3196
timestamp 1745462530
transform 1 0 844 0 1 2765
box -3 -3 3 3
use M3_M2  M3_M2_3197
timestamp 1745462530
transform 1 0 772 0 1 2715
box -3 -3 3 3
use M3_M2  M3_M2_3198
timestamp 1745462530
transform 1 0 660 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_3199
timestamp 1745462530
transform 1 0 476 0 1 2715
box -3 -3 3 3
use M3_M2  M3_M2_3200
timestamp 1745462530
transform 1 0 476 0 1 2665
box -3 -3 3 3
use M3_M2  M3_M2_3201
timestamp 1745462530
transform 1 0 228 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_3202
timestamp 1745462530
transform 1 0 220 0 1 2665
box -3 -3 3 3
use M3_M2  M3_M2_3203
timestamp 1745462530
transform 1 0 212 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_3204
timestamp 1745462530
transform 1 0 204 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_3205
timestamp 1745462530
transform 1 0 196 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_3206
timestamp 1745462530
transform 1 0 172 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_3207
timestamp 1745462530
transform 1 0 164 0 1 2665
box -3 -3 3 3
use M3_M2  M3_M2_3208
timestamp 1745462530
transform 1 0 164 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_3209
timestamp 1745462530
transform 1 0 164 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_3210
timestamp 1745462530
transform 1 0 1428 0 1 325
box -3 -3 3 3
use M3_M2  M3_M2_3211
timestamp 1745462530
transform 1 0 1356 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_3212
timestamp 1745462530
transform 1 0 1300 0 1 325
box -3 -3 3 3
use M3_M2  M3_M2_3213
timestamp 1745462530
transform 1 0 1292 0 1 375
box -3 -3 3 3
use M3_M2  M3_M2_3214
timestamp 1745462530
transform 1 0 1156 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_3215
timestamp 1745462530
transform 1 0 1156 0 1 375
box -3 -3 3 3
use M3_M2  M3_M2_3216
timestamp 1745462530
transform 1 0 1132 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_3217
timestamp 1745462530
transform 1 0 932 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_3218
timestamp 1745462530
transform 1 0 916 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_3219
timestamp 1745462530
transform 1 0 668 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_3220
timestamp 1745462530
transform 1 0 236 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_3221
timestamp 1745462530
transform 1 0 236 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_3222
timestamp 1745462530
transform 1 0 212 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_3223
timestamp 1745462530
transform 1 0 196 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_3224
timestamp 1745462530
transform 1 0 196 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_3225
timestamp 1745462530
transform 1 0 3308 0 1 255
box -3 -3 3 3
use M3_M2  M3_M2_3226
timestamp 1745462530
transform 1 0 2604 0 1 275
box -3 -3 3 3
use M3_M2  M3_M2_3227
timestamp 1745462530
transform 1 0 2604 0 1 255
box -3 -3 3 3
use M3_M2  M3_M2_3228
timestamp 1745462530
transform 1 0 2556 0 1 1065
box -3 -3 3 3
use M3_M2  M3_M2_3229
timestamp 1745462530
transform 1 0 2444 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_3230
timestamp 1745462530
transform 1 0 2404 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_3231
timestamp 1745462530
transform 1 0 2356 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_3232
timestamp 1745462530
transform 1 0 2356 0 1 1215
box -3 -3 3 3
use M3_M2  M3_M2_3233
timestamp 1745462530
transform 1 0 2356 0 1 1065
box -3 -3 3 3
use M3_M2  M3_M2_3234
timestamp 1745462530
transform 1 0 2316 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_3235
timestamp 1745462530
transform 1 0 2316 0 1 1215
box -3 -3 3 3
use M3_M2  M3_M2_3236
timestamp 1745462530
transform 1 0 2292 0 1 275
box -3 -3 3 3
use M3_M2  M3_M2_3237
timestamp 1745462530
transform 1 0 2284 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_3238
timestamp 1745462530
transform 1 0 2236 0 1 1065
box -3 -3 3 3
use M3_M2  M3_M2_3239
timestamp 1745462530
transform 1 0 2220 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_3240
timestamp 1745462530
transform 1 0 2196 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_3241
timestamp 1745462530
transform 1 0 1916 0 1 1435
box -3 -3 3 3
use M3_M2  M3_M2_3242
timestamp 1745462530
transform 1 0 1900 0 1 1405
box -3 -3 3 3
use M3_M2  M3_M2_3243
timestamp 1745462530
transform 1 0 1852 0 1 1405
box -3 -3 3 3
use M3_M2  M3_M2_3244
timestamp 1745462530
transform 1 0 1852 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_3245
timestamp 1745462530
transform 1 0 1828 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_3246
timestamp 1745462530
transform 1 0 1828 0 1 1275
box -3 -3 3 3
use M3_M2  M3_M2_3247
timestamp 1745462530
transform 1 0 1532 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_3248
timestamp 1745462530
transform 1 0 1532 0 1 1275
box -3 -3 3 3
use M3_M2  M3_M2_3249
timestamp 1745462530
transform 1 0 1516 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_3250
timestamp 1745462530
transform 1 0 1452 0 1 1265
box -3 -3 3 3
use M3_M2  M3_M2_3251
timestamp 1745462530
transform 1 0 1420 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_3252
timestamp 1745462530
transform 1 0 1356 0 1 1265
box -3 -3 3 3
use M3_M2  M3_M2_3253
timestamp 1745462530
transform 1 0 1356 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_3254
timestamp 1745462530
transform 1 0 4196 0 1 2015
box -3 -3 3 3
use M3_M2  M3_M2_3255
timestamp 1745462530
transform 1 0 4196 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_3256
timestamp 1745462530
transform 1 0 4148 0 1 2015
box -3 -3 3 3
use M3_M2  M3_M2_3257
timestamp 1745462530
transform 1 0 4116 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_3258
timestamp 1745462530
transform 1 0 4116 0 1 1775
box -3 -3 3 3
use M3_M2  M3_M2_3259
timestamp 1745462530
transform 1 0 4100 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_3260
timestamp 1745462530
transform 1 0 4076 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_3261
timestamp 1745462530
transform 1 0 4060 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_3262
timestamp 1745462530
transform 1 0 4060 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_3263
timestamp 1745462530
transform 1 0 4020 0 1 1775
box -3 -3 3 3
use M3_M2  M3_M2_3264
timestamp 1745462530
transform 1 0 4020 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_3265
timestamp 1745462530
transform 1 0 4020 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_3266
timestamp 1745462530
transform 1 0 4004 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_3267
timestamp 1745462530
transform 1 0 3956 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_3268
timestamp 1745462530
transform 1 0 3956 0 1 875
box -3 -3 3 3
use M3_M2  M3_M2_3269
timestamp 1745462530
transform 1 0 3956 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_3270
timestamp 1745462530
transform 1 0 3668 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_3271
timestamp 1745462530
transform 1 0 3564 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_3272
timestamp 1745462530
transform 1 0 3564 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_3273
timestamp 1745462530
transform 1 0 3500 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_3274
timestamp 1745462530
transform 1 0 3500 0 1 875
box -3 -3 3 3
use M3_M2  M3_M2_3275
timestamp 1745462530
transform 1 0 3468 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_3276
timestamp 1745462530
transform 1 0 3452 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_3277
timestamp 1745462530
transform 1 0 3324 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_3278
timestamp 1745462530
transform 1 0 3460 0 1 2495
box -3 -3 3 3
use M3_M2  M3_M2_3279
timestamp 1745462530
transform 1 0 3428 0 1 2495
box -3 -3 3 3
use M3_M2  M3_M2_3280
timestamp 1745462530
transform 1 0 3420 0 1 2895
box -3 -3 3 3
use M3_M2  M3_M2_3281
timestamp 1745462530
transform 1 0 3388 0 1 2895
box -3 -3 3 3
use M3_M2  M3_M2_3282
timestamp 1745462530
transform 1 0 3276 0 1 2895
box -3 -3 3 3
use M3_M2  M3_M2_3283
timestamp 1745462530
transform 1 0 3212 0 1 2895
box -3 -3 3 3
use M3_M2  M3_M2_3284
timestamp 1745462530
transform 1 0 2852 0 1 2235
box -3 -3 3 3
use M3_M2  M3_M2_3285
timestamp 1745462530
transform 1 0 2820 0 1 2895
box -3 -3 3 3
use M3_M2  M3_M2_3286
timestamp 1745462530
transform 1 0 2820 0 1 2785
box -3 -3 3 3
use M3_M2  M3_M2_3287
timestamp 1745462530
transform 1 0 2772 0 1 2785
box -3 -3 3 3
use M3_M2  M3_M2_3288
timestamp 1745462530
transform 1 0 2764 0 1 2235
box -3 -3 3 3
use M3_M2  M3_M2_3289
timestamp 1745462530
transform 1 0 2724 0 1 2235
box -3 -3 3 3
use M3_M2  M3_M2_3290
timestamp 1745462530
transform 1 0 2692 0 1 2785
box -3 -3 3 3
use M3_M2  M3_M2_3291
timestamp 1745462530
transform 1 0 2628 0 1 2235
box -3 -3 3 3
use M3_M2  M3_M2_3292
timestamp 1745462530
transform 1 0 1164 0 1 2065
box -3 -3 3 3
use M3_M2  M3_M2_3293
timestamp 1745462530
transform 1 0 1132 0 1 2065
box -3 -3 3 3
use M3_M2  M3_M2_3294
timestamp 1745462530
transform 1 0 3252 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_3295
timestamp 1745462530
transform 1 0 2852 0 1 2095
box -3 -3 3 3
use M3_M2  M3_M2_3296
timestamp 1745462530
transform 1 0 2852 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_3297
timestamp 1745462530
transform 1 0 2836 0 1 2095
box -3 -3 3 3
use M3_M2  M3_M2_3298
timestamp 1745462530
transform 1 0 2764 0 1 2095
box -3 -3 3 3
use M3_M2  M3_M2_3299
timestamp 1745462530
transform 1 0 2764 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_3300
timestamp 1745462530
transform 1 0 2428 0 1 1975
box -3 -3 3 3
use M3_M2  M3_M2_3301
timestamp 1745462530
transform 1 0 2388 0 1 1975
box -3 -3 3 3
use M3_M2  M3_M2_3302
timestamp 1745462530
transform 1 0 1876 0 1 2245
box -3 -3 3 3
use M3_M2  M3_M2_3303
timestamp 1745462530
transform 1 0 1860 0 1 2245
box -3 -3 3 3
use M3_M2  M3_M2_3304
timestamp 1745462530
transform 1 0 1844 0 1 1855
box -3 -3 3 3
use M3_M2  M3_M2_3305
timestamp 1745462530
transform 1 0 1796 0 1 1855
box -3 -3 3 3
use M3_M2  M3_M2_3306
timestamp 1745462530
transform 1 0 1796 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_3307
timestamp 1745462530
transform 1 0 1708 0 1 2545
box -3 -3 3 3
use M3_M2  M3_M2_3308
timestamp 1745462530
transform 1 0 1020 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_3309
timestamp 1745462530
transform 1 0 1020 0 1 1695
box -3 -3 3 3
use M3_M2  M3_M2_3310
timestamp 1745462530
transform 1 0 884 0 1 2915
box -3 -3 3 3
use M3_M2  M3_M2_3311
timestamp 1745462530
transform 1 0 764 0 1 2925
box -3 -3 3 3
use M3_M2  M3_M2_3312
timestamp 1745462530
transform 1 0 660 0 1 2915
box -3 -3 3 3
use M3_M2  M3_M2_3313
timestamp 1745462530
transform 1 0 660 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_3314
timestamp 1745462530
transform 1 0 660 0 1 1695
box -3 -3 3 3
use M3_M2  M3_M2_3315
timestamp 1745462530
transform 1 0 460 0 1 2545
box -3 -3 3 3
use M3_M2  M3_M2_3316
timestamp 1745462530
transform 1 0 460 0 1 2475
box -3 -3 3 3
use M3_M2  M3_M2_3317
timestamp 1745462530
transform 1 0 444 0 1 2915
box -3 -3 3 3
use M3_M2  M3_M2_3318
timestamp 1745462530
transform 1 0 396 0 1 2295
box -3 -3 3 3
use M3_M2  M3_M2_3319
timestamp 1745462530
transform 1 0 388 0 1 2475
box -3 -3 3 3
use M3_M2  M3_M2_3320
timestamp 1745462530
transform 1 0 340 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_3321
timestamp 1745462530
transform 1 0 324 0 1 2295
box -3 -3 3 3
use M3_M2  M3_M2_3322
timestamp 1745462530
transform 1 0 1900 0 1 675
box -3 -3 3 3
use M3_M2  M3_M2_3323
timestamp 1745462530
transform 1 0 1884 0 1 675
box -3 -3 3 3
use M3_M2  M3_M2_3324
timestamp 1745462530
transform 1 0 1884 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_3325
timestamp 1745462530
transform 1 0 1804 0 1 1405
box -3 -3 3 3
use M3_M2  M3_M2_3326
timestamp 1745462530
transform 1 0 1620 0 1 335
box -3 -3 3 3
use M3_M2  M3_M2_3327
timestamp 1745462530
transform 1 0 900 0 1 335
box -3 -3 3 3
use M3_M2  M3_M2_3328
timestamp 1745462530
transform 1 0 844 0 1 1405
box -3 -3 3 3
use M3_M2  M3_M2_3329
timestamp 1745462530
transform 1 0 692 0 1 335
box -3 -3 3 3
use M3_M2  M3_M2_3330
timestamp 1745462530
transform 1 0 404 0 1 1405
box -3 -3 3 3
use M3_M2  M3_M2_3331
timestamp 1745462530
transform 1 0 404 0 1 1205
box -3 -3 3 3
use M3_M2  M3_M2_3332
timestamp 1745462530
transform 1 0 204 0 1 335
box -3 -3 3 3
use M3_M2  M3_M2_3333
timestamp 1745462530
transform 1 0 196 0 1 1205
box -3 -3 3 3
use M3_M2  M3_M2_3334
timestamp 1745462530
transform 1 0 3364 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_3335
timestamp 1745462530
transform 1 0 2604 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_3336
timestamp 1745462530
transform 1 0 2588 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_3337
timestamp 1745462530
transform 1 0 2452 0 1 335
box -3 -3 3 3
use M3_M2  M3_M2_3338
timestamp 1745462530
transform 1 0 2348 0 1 335
box -3 -3 3 3
use M3_M2  M3_M2_3339
timestamp 1745462530
transform 1 0 2340 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_3340
timestamp 1745462530
transform 1 0 2300 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_3341
timestamp 1745462530
transform 1 0 2284 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_3342
timestamp 1745462530
transform 1 0 2284 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_3343
timestamp 1745462530
transform 1 0 2284 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_3344
timestamp 1745462530
transform 1 0 2252 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_3345
timestamp 1745462530
transform 1 0 2252 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_3346
timestamp 1745462530
transform 1 0 2204 0 1 1375
box -3 -3 3 3
use M3_M2  M3_M2_3347
timestamp 1745462530
transform 1 0 2204 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_3348
timestamp 1745462530
transform 1 0 2204 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_3349
timestamp 1745462530
transform 1 0 1996 0 1 1375
box -3 -3 3 3
use M3_M2  M3_M2_3350
timestamp 1745462530
transform 1 0 4188 0 1 455
box -3 -3 3 3
use M3_M2  M3_M2_3351
timestamp 1745462530
transform 1 0 4180 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_3352
timestamp 1745462530
transform 1 0 4172 0 1 1465
box -3 -3 3 3
use M3_M2  M3_M2_3353
timestamp 1745462530
transform 1 0 4148 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_3354
timestamp 1745462530
transform 1 0 4132 0 1 1465
box -3 -3 3 3
use M3_M2  M3_M2_3355
timestamp 1745462530
transform 1 0 3980 0 1 1465
box -3 -3 3 3
use M3_M2  M3_M2_3356
timestamp 1745462530
transform 1 0 3804 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_3357
timestamp 1745462530
transform 1 0 3796 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_3358
timestamp 1745462530
transform 1 0 3780 0 1 1475
box -3 -3 3 3
use M3_M2  M3_M2_3359
timestamp 1745462530
transform 1 0 3780 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_3360
timestamp 1745462530
transform 1 0 3756 0 1 455
box -3 -3 3 3
use M3_M2  M3_M2_3361
timestamp 1745462530
transform 1 0 3756 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_3362
timestamp 1745462530
transform 1 0 3740 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_3363
timestamp 1745462530
transform 1 0 2764 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_3364
timestamp 1745462530
transform 1 0 3948 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_3365
timestamp 1745462530
transform 1 0 3948 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_3366
timestamp 1745462530
transform 1 0 3940 0 1 2455
box -3 -3 3 3
use M3_M2  M3_M2_3367
timestamp 1745462530
transform 1 0 3932 0 1 2245
box -3 -3 3 3
use M3_M2  M3_M2_3368
timestamp 1745462530
transform 1 0 3876 0 1 2245
box -3 -3 3 3
use M3_M2  M3_M2_3369
timestamp 1745462530
transform 1 0 3876 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_3370
timestamp 1745462530
transform 1 0 3876 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_3371
timestamp 1745462530
transform 1 0 3844 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_3372
timestamp 1745462530
transform 1 0 3844 0 1 2935
box -3 -3 3 3
use M3_M2  M3_M2_3373
timestamp 1745462530
transform 1 0 3836 0 1 2455
box -3 -3 3 3
use M3_M2  M3_M2_3374
timestamp 1745462530
transform 1 0 3764 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_3375
timestamp 1745462530
transform 1 0 3732 0 1 2935
box -3 -3 3 3
use M3_M2  M3_M2_3376
timestamp 1745462530
transform 1 0 2996 0 1 2095
box -3 -3 3 3
use M3_M2  M3_M2_3377
timestamp 1745462530
transform 1 0 2996 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_3378
timestamp 1745462530
transform 1 0 2972 0 1 2095
box -3 -3 3 3
use M3_M2  M3_M2_3379
timestamp 1745462530
transform 1 0 2972 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_3380
timestamp 1745462530
transform 1 0 2972 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_3381
timestamp 1745462530
transform 1 0 2940 0 1 2445
box -3 -3 3 3
use M3_M2  M3_M2_3382
timestamp 1745462530
transform 1 0 2924 0 1 2875
box -3 -3 3 3
use M3_M2  M3_M2_3383
timestamp 1745462530
transform 1 0 2716 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_3384
timestamp 1745462530
transform 1 0 2500 0 1 2875
box -3 -3 3 3
use M3_M2  M3_M2_3385
timestamp 1745462530
transform 1 0 1860 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_3386
timestamp 1745462530
transform 1 0 1788 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_3387
timestamp 1745462530
transform 1 0 2700 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_3388
timestamp 1745462530
transform 1 0 2188 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_3389
timestamp 1745462530
transform 1 0 2148 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_3390
timestamp 1745462530
transform 1 0 2148 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_3391
timestamp 1745462530
transform 1 0 1740 0 1 2765
box -3 -3 3 3
use M3_M2  M3_M2_3392
timestamp 1745462530
transform 1 0 1716 0 1 2165
box -3 -3 3 3
use M3_M2  M3_M2_3393
timestamp 1745462530
transform 1 0 1692 0 1 2165
box -3 -3 3 3
use M3_M2  M3_M2_3394
timestamp 1745462530
transform 1 0 1684 0 1 2765
box -3 -3 3 3
use M3_M2  M3_M2_3395
timestamp 1745462530
transform 1 0 1708 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_3396
timestamp 1745462530
transform 1 0 1564 0 1 2055
box -3 -3 3 3
use M3_M2  M3_M2_3397
timestamp 1745462530
transform 1 0 1564 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_3398
timestamp 1745462530
transform 1 0 1540 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_3399
timestamp 1745462530
transform 1 0 1532 0 1 2055
box -3 -3 3 3
use M3_M2  M3_M2_3400
timestamp 1745462530
transform 1 0 1452 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_3401
timestamp 1745462530
transform 1 0 1452 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_3402
timestamp 1745462530
transform 1 0 956 0 1 2565
box -3 -3 3 3
use M3_M2  M3_M2_3403
timestamp 1745462530
transform 1 0 916 0 1 2565
box -3 -3 3 3
use M3_M2  M3_M2_3404
timestamp 1745462530
transform 1 0 900 0 1 2475
box -3 -3 3 3
use M3_M2  M3_M2_3405
timestamp 1745462530
transform 1 0 804 0 1 2475
box -3 -3 3 3
use M3_M2  M3_M2_3406
timestamp 1745462530
transform 1 0 804 0 1 2365
box -3 -3 3 3
use M3_M2  M3_M2_3407
timestamp 1745462530
transform 1 0 556 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_3408
timestamp 1745462530
transform 1 0 548 0 1 2065
box -3 -3 3 3
use M3_M2  M3_M2_3409
timestamp 1745462530
transform 1 0 532 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_3410
timestamp 1745462530
transform 1 0 492 0 1 2565
box -3 -3 3 3
use M3_M2  M3_M2_3411
timestamp 1745462530
transform 1 0 452 0 1 2235
box -3 -3 3 3
use M3_M2  M3_M2_3412
timestamp 1745462530
transform 1 0 452 0 1 2065
box -3 -3 3 3
use M3_M2  M3_M2_3413
timestamp 1745462530
transform 1 0 428 0 1 2565
box -3 -3 3 3
use M3_M2  M3_M2_3414
timestamp 1745462530
transform 1 0 420 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_3415
timestamp 1745462530
transform 1 0 348 0 1 2365
box -3 -3 3 3
use M3_M2  M3_M2_3416
timestamp 1745462530
transform 1 0 348 0 1 2235
box -3 -3 3 3
use M3_M2  M3_M2_3417
timestamp 1745462530
transform 1 0 340 0 1 2565
box -3 -3 3 3
use M3_M2  M3_M2_3418
timestamp 1745462530
transform 1 0 1876 0 1 175
box -3 -3 3 3
use M3_M2  M3_M2_3419
timestamp 1745462530
transform 1 0 1820 0 1 175
box -3 -3 3 3
use M3_M2  M3_M2_3420
timestamp 1745462530
transform 1 0 1780 0 1 175
box -3 -3 3 3
use M3_M2  M3_M2_3421
timestamp 1745462530
transform 1 0 1692 0 1 1485
box -3 -3 3 3
use M3_M2  M3_M2_3422
timestamp 1745462530
transform 1 0 1684 0 1 175
box -3 -3 3 3
use M3_M2  M3_M2_3423
timestamp 1745462530
transform 1 0 812 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_3424
timestamp 1745462530
transform 1 0 740 0 1 1485
box -3 -3 3 3
use M3_M2  M3_M2_3425
timestamp 1745462530
transform 1 0 740 0 1 1455
box -3 -3 3 3
use M3_M2  M3_M2_3426
timestamp 1745462530
transform 1 0 540 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_3427
timestamp 1745462530
transform 1 0 372 0 1 1005
box -3 -3 3 3
use M3_M2  M3_M2_3428
timestamp 1745462530
transform 1 0 372 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_3429
timestamp 1745462530
transform 1 0 316 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_3430
timestamp 1745462530
transform 1 0 308 0 1 1455
box -3 -3 3 3
use M3_M2  M3_M2_3431
timestamp 1745462530
transform 1 0 292 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_3432
timestamp 1745462530
transform 1 0 284 0 1 1005
box -3 -3 3 3
use M3_M2  M3_M2_3433
timestamp 1745462530
transform 1 0 252 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_3434
timestamp 1745462530
transform 1 0 252 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_3435
timestamp 1745462530
transform 1 0 3404 0 1 175
box -3 -3 3 3
use M3_M2  M3_M2_3436
timestamp 1745462530
transform 1 0 2500 0 1 165
box -3 -3 3 3
use M3_M2  M3_M2_3437
timestamp 1745462530
transform 1 0 2364 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_3438
timestamp 1745462530
transform 1 0 2348 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_3439
timestamp 1745462530
transform 1 0 2348 0 1 845
box -3 -3 3 3
use M3_M2  M3_M2_3440
timestamp 1745462530
transform 1 0 2292 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_3441
timestamp 1745462530
transform 1 0 2228 0 1 845
box -3 -3 3 3
use M3_M2  M3_M2_3442
timestamp 1745462530
transform 1 0 2228 0 1 165
box -3 -3 3 3
use M3_M2  M3_M2_3443
timestamp 1745462530
transform 1 0 2220 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_3444
timestamp 1745462530
transform 1 0 2220 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_3445
timestamp 1745462530
transform 1 0 2020 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_3446
timestamp 1745462530
transform 1 0 1996 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_3447
timestamp 1745462530
transform 1 0 1996 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_3448
timestamp 1745462530
transform 1 0 1996 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_3449
timestamp 1745462530
transform 1 0 1980 0 1 1405
box -3 -3 3 3
use M3_M2  M3_M2_3450
timestamp 1745462530
transform 1 0 1980 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_3451
timestamp 1745462530
transform 1 0 1924 0 1 1405
box -3 -3 3 3
use M3_M2  M3_M2_3452
timestamp 1745462530
transform 1 0 4356 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_3453
timestamp 1745462530
transform 1 0 4356 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_3454
timestamp 1745462530
transform 1 0 4316 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_3455
timestamp 1745462530
transform 1 0 4308 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_3456
timestamp 1745462530
transform 1 0 4308 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_3457
timestamp 1745462530
transform 1 0 4252 0 1 1295
box -3 -3 3 3
use M3_M2  M3_M2_3458
timestamp 1745462530
transform 1 0 4244 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_3459
timestamp 1745462530
transform 1 0 4244 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_3460
timestamp 1745462530
transform 1 0 4220 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_3461
timestamp 1745462530
transform 1 0 4220 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_3462
timestamp 1745462530
transform 1 0 4220 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_3463
timestamp 1745462530
transform 1 0 4180 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_3464
timestamp 1745462530
transform 1 0 3964 0 1 215
box -3 -3 3 3
use M3_M2  M3_M2_3465
timestamp 1745462530
transform 1 0 3916 0 1 1295
box -3 -3 3 3
use M3_M2  M3_M2_3466
timestamp 1745462530
transform 1 0 3820 0 1 215
box -3 -3 3 3
use M3_M2  M3_M2_3467
timestamp 1745462530
transform 1 0 3668 0 1 1295
box -3 -3 3 3
use M3_M2  M3_M2_3468
timestamp 1745462530
transform 1 0 3636 0 1 1645
box -3 -3 3 3
use M3_M2  M3_M2_3469
timestamp 1745462530
transform 1 0 2860 0 1 1645
box -3 -3 3 3
use M3_M2  M3_M2_3470
timestamp 1745462530
transform 1 0 2860 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_3471
timestamp 1745462530
transform 1 0 2724 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_3472
timestamp 1745462530
transform 1 0 4276 0 1 2905
box -3 -3 3 3
use M3_M2  M3_M2_3473
timestamp 1745462530
transform 1 0 4276 0 1 2715
box -3 -3 3 3
use M3_M2  M3_M2_3474
timestamp 1745462530
transform 1 0 4220 0 1 2905
box -3 -3 3 3
use M3_M2  M3_M2_3475
timestamp 1745462530
transform 1 0 4220 0 1 2525
box -3 -3 3 3
use M3_M2  M3_M2_3476
timestamp 1745462530
transform 1 0 4220 0 1 2405
box -3 -3 3 3
use M3_M2  M3_M2_3477
timestamp 1745462530
transform 1 0 4196 0 1 2715
box -3 -3 3 3
use M3_M2  M3_M2_3478
timestamp 1745462530
transform 1 0 4196 0 1 2655
box -3 -3 3 3
use M3_M2  M3_M2_3479
timestamp 1745462530
transform 1 0 4196 0 1 2545
box -3 -3 3 3
use M3_M2  M3_M2_3480
timestamp 1745462530
transform 1 0 4180 0 1 2405
box -3 -3 3 3
use M3_M2  M3_M2_3481
timestamp 1745462530
transform 1 0 4140 0 1 2905
box -3 -3 3 3
use M3_M2  M3_M2_3482
timestamp 1745462530
transform 1 0 4052 0 1 2895
box -3 -3 3 3
use M3_M2  M3_M2_3483
timestamp 1745462530
transform 1 0 3900 0 1 2895
box -3 -3 3 3
use M3_M2  M3_M2_3484
timestamp 1745462530
transform 1 0 3244 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_3485
timestamp 1745462530
transform 1 0 2868 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_3486
timestamp 1745462530
transform 1 0 2852 0 1 2255
box -3 -3 3 3
use M3_M2  M3_M2_3487
timestamp 1745462530
transform 1 0 2828 0 1 2545
box -3 -3 3 3
use M3_M2  M3_M2_3488
timestamp 1745462530
transform 1 0 2828 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_3489
timestamp 1745462530
transform 1 0 2828 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_3490
timestamp 1745462530
transform 1 0 2804 0 1 2655
box -3 -3 3 3
use M3_M2  M3_M2_3491
timestamp 1745462530
transform 1 0 2804 0 1 2545
box -3 -3 3 3
use M3_M2  M3_M2_3492
timestamp 1745462530
transform 1 0 2756 0 1 2845
box -3 -3 3 3
use M3_M2  M3_M2_3493
timestamp 1745462530
transform 1 0 2756 0 1 2655
box -3 -3 3 3
use M3_M2  M3_M2_3494
timestamp 1745462530
transform 1 0 2748 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_3495
timestamp 1745462530
transform 1 0 2740 0 1 2255
box -3 -3 3 3
use M3_M2  M3_M2_3496
timestamp 1745462530
transform 1 0 2732 0 1 1875
box -3 -3 3 3
use M3_M2  M3_M2_3497
timestamp 1745462530
transform 1 0 2668 0 1 1875
box -3 -3 3 3
use M3_M2  M3_M2_3498
timestamp 1745462530
transform 1 0 2612 0 1 2845
box -3 -3 3 3
use M3_M2  M3_M2_3499
timestamp 1745462530
transform 1 0 1708 0 1 1665
box -3 -3 3 3
use M3_M2  M3_M2_3500
timestamp 1745462530
transform 1 0 1684 0 1 1665
box -3 -3 3 3
use M3_M2  M3_M2_3501
timestamp 1745462530
transform 1 0 2724 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_3502
timestamp 1745462530
transform 1 0 2692 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_3503
timestamp 1745462530
transform 1 0 2324 0 1 1615
box -3 -3 3 3
use M3_M2  M3_M2_3504
timestamp 1745462530
transform 1 0 2324 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_3505
timestamp 1745462530
transform 1 0 2292 0 1 1655
box -3 -3 3 3
use M3_M2  M3_M2_3506
timestamp 1745462530
transform 1 0 2292 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_3507
timestamp 1745462530
transform 1 0 2188 0 1 1655
box -3 -3 3 3
use M3_M2  M3_M2_3508
timestamp 1745462530
transform 1 0 1324 0 1 2185
box -3 -3 3 3
use M3_M2  M3_M2_3509
timestamp 1745462530
transform 1 0 1324 0 1 2075
box -3 -3 3 3
use M3_M2  M3_M2_3510
timestamp 1745462530
transform 1 0 1292 0 1 2185
box -3 -3 3 3
use M3_M2  M3_M2_3511
timestamp 1745462530
transform 1 0 1284 0 1 2075
box -3 -3 3 3
use M3_M2  M3_M2_3512
timestamp 1745462530
transform 1 0 1236 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_3513
timestamp 1745462530
transform 1 0 1204 0 1 1865
box -3 -3 3 3
use M3_M2  M3_M2_3514
timestamp 1745462530
transform 1 0 1204 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_3515
timestamp 1745462530
transform 1 0 1196 0 1 2675
box -3 -3 3 3
use M3_M2  M3_M2_3516
timestamp 1745462530
transform 1 0 1108 0 1 2675
box -3 -3 3 3
use M3_M2  M3_M2_3517
timestamp 1745462530
transform 1 0 1092 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_3518
timestamp 1745462530
transform 1 0 1028 0 1 1875
box -3 -3 3 3
use M3_M2  M3_M2_3519
timestamp 1745462530
transform 1 0 1028 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_3520
timestamp 1745462530
transform 1 0 956 0 1 2975
box -3 -3 3 3
use M3_M2  M3_M2_3521
timestamp 1745462530
transform 1 0 956 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_3522
timestamp 1745462530
transform 1 0 684 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_3523
timestamp 1745462530
transform 1 0 532 0 1 2975
box -3 -3 3 3
use M3_M2  M3_M2_3524
timestamp 1745462530
transform 1 0 532 0 1 2805
box -3 -3 3 3
use M3_M2  M3_M2_3525
timestamp 1745462530
transform 1 0 468 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_3526
timestamp 1745462530
transform 1 0 420 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_3527
timestamp 1745462530
transform 1 0 404 0 1 2155
box -3 -3 3 3
use M3_M2  M3_M2_3528
timestamp 1745462530
transform 1 0 388 0 1 2805
box -3 -3 3 3
use M3_M2  M3_M2_3529
timestamp 1745462530
transform 1 0 388 0 1 2705
box -3 -3 3 3
use M3_M2  M3_M2_3530
timestamp 1745462530
transform 1 0 372 0 1 2705
box -3 -3 3 3
use M3_M2  M3_M2_3531
timestamp 1745462530
transform 1 0 372 0 1 2605
box -3 -3 3 3
use M3_M2  M3_M2_3532
timestamp 1745462530
transform 1 0 356 0 1 2605
box -3 -3 3 3
use M3_M2  M3_M2_3533
timestamp 1745462530
transform 1 0 356 0 1 2155
box -3 -3 3 3
use M3_M2  M3_M2_3534
timestamp 1745462530
transform 1 0 292 0 1 2805
box -3 -3 3 3
use M3_M2  M3_M2_3535
timestamp 1745462530
transform 1 0 1452 0 1 245
box -3 -3 3 3
use M3_M2  M3_M2_3536
timestamp 1745462530
transform 1 0 1412 0 1 1415
box -3 -3 3 3
use M3_M2  M3_M2_3537
timestamp 1745462530
transform 1 0 1396 0 1 245
box -3 -3 3 3
use M3_M2  M3_M2_3538
timestamp 1745462530
transform 1 0 1292 0 1 1415
box -3 -3 3 3
use M3_M2  M3_M2_3539
timestamp 1745462530
transform 1 0 1140 0 1 235
box -3 -3 3 3
use M3_M2  M3_M2_3540
timestamp 1745462530
transform 1 0 900 0 1 235
box -3 -3 3 3
use M3_M2  M3_M2_3541
timestamp 1745462530
transform 1 0 900 0 1 205
box -3 -3 3 3
use M3_M2  M3_M2_3542
timestamp 1745462530
transform 1 0 700 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_3543
timestamp 1745462530
transform 1 0 636 0 1 205
box -3 -3 3 3
use M3_M2  M3_M2_3544
timestamp 1745462530
transform 1 0 404 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_3545
timestamp 1745462530
transform 1 0 404 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_3546
timestamp 1745462530
transform 1 0 396 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_3547
timestamp 1745462530
transform 1 0 396 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_3548
timestamp 1745462530
transform 1 0 396 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_3549
timestamp 1745462530
transform 1 0 380 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_3550
timestamp 1745462530
transform 1 0 380 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_3551
timestamp 1745462530
transform 1 0 380 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_3552
timestamp 1745462530
transform 1 0 332 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_3553
timestamp 1745462530
transform 1 0 324 0 1 205
box -3 -3 3 3
use M3_M2  M3_M2_3554
timestamp 1745462530
transform 1 0 3252 0 1 415
box -3 -3 3 3
use M3_M2  M3_M2_3555
timestamp 1745462530
transform 1 0 3068 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_3556
timestamp 1745462530
transform 1 0 3060 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_3557
timestamp 1745462530
transform 1 0 3012 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_3558
timestamp 1745462530
transform 1 0 3012 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_3559
timestamp 1745462530
transform 1 0 2980 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_3560
timestamp 1745462530
transform 1 0 2980 0 1 415
box -3 -3 3 3
use M3_M2  M3_M2_3561
timestamp 1745462530
transform 1 0 2956 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_3562
timestamp 1745462530
transform 1 0 2956 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_3563
timestamp 1745462530
transform 1 0 2900 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_3564
timestamp 1745462530
transform 1 0 2836 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_3565
timestamp 1745462530
transform 1 0 2820 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_3566
timestamp 1745462530
transform 1 0 2636 0 1 415
box -3 -3 3 3
use M3_M2  M3_M2_3567
timestamp 1745462530
transform 1 0 2596 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_3568
timestamp 1745462530
transform 1 0 1668 0 1 1415
box -3 -3 3 3
use M3_M2  M3_M2_3569
timestamp 1745462530
transform 1 0 1636 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_3570
timestamp 1745462530
transform 1 0 1604 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_3571
timestamp 1745462530
transform 1 0 1604 0 1 1075
box -3 -3 3 3
use M3_M2  M3_M2_3572
timestamp 1745462530
transform 1 0 1588 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_3573
timestamp 1745462530
transform 1 0 1588 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_3574
timestamp 1745462530
transform 1 0 1588 0 1 1075
box -3 -3 3 3
use M3_M2  M3_M2_3575
timestamp 1745462530
transform 1 0 4164 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_3576
timestamp 1745462530
transform 1 0 4140 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_3577
timestamp 1745462530
transform 1 0 4140 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_3578
timestamp 1745462530
transform 1 0 4124 0 1 645
box -3 -3 3 3
use M3_M2  M3_M2_3579
timestamp 1745462530
transform 1 0 4124 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_3580
timestamp 1745462530
transform 1 0 4100 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_3581
timestamp 1745462530
transform 1 0 4100 0 1 975
box -3 -3 3 3
use M3_M2  M3_M2_3582
timestamp 1745462530
transform 1 0 4076 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_3583
timestamp 1745462530
transform 1 0 4068 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_3584
timestamp 1745462530
transform 1 0 4060 0 1 645
box -3 -3 3 3
use M3_M2  M3_M2_3585
timestamp 1745462530
transform 1 0 4060 0 1 405
box -3 -3 3 3
use M3_M2  M3_M2_3586
timestamp 1745462530
transform 1 0 4052 0 1 975
box -3 -3 3 3
use M3_M2  M3_M2_3587
timestamp 1745462530
transform 1 0 3540 0 1 1525
box -3 -3 3 3
use M3_M2  M3_M2_3588
timestamp 1745462530
transform 1 0 3540 0 1 1465
box -3 -3 3 3
use M3_M2  M3_M2_3589
timestamp 1745462530
transform 1 0 3492 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_3590
timestamp 1745462530
transform 1 0 3484 0 1 1465
box -3 -3 3 3
use M3_M2  M3_M2_3591
timestamp 1745462530
transform 1 0 3372 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_3592
timestamp 1745462530
transform 1 0 3356 0 1 405
box -3 -3 3 3
use M3_M2  M3_M2_3593
timestamp 1745462530
transform 1 0 2908 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_3594
timestamp 1745462530
transform 1 0 3284 0 1 2435
box -3 -3 3 3
use M3_M2  M3_M2_3595
timestamp 1745462530
transform 1 0 3276 0 1 2275
box -3 -3 3 3
use M3_M2  M3_M2_3596
timestamp 1745462530
transform 1 0 3276 0 1 1665
box -3 -3 3 3
use M3_M2  M3_M2_3597
timestamp 1745462530
transform 1 0 3236 0 1 2275
box -3 -3 3 3
use M3_M2  M3_M2_3598
timestamp 1745462530
transform 1 0 3228 0 1 2925
box -3 -3 3 3
use M3_M2  M3_M2_3599
timestamp 1745462530
transform 1 0 3212 0 1 3015
box -3 -3 3 3
use M3_M2  M3_M2_3600
timestamp 1745462530
transform 1 0 3196 0 1 2435
box -3 -3 3 3
use M3_M2  M3_M2_3601
timestamp 1745462530
transform 1 0 3188 0 1 2925
box -3 -3 3 3
use M3_M2  M3_M2_3602
timestamp 1745462530
transform 1 0 3172 0 1 1665
box -3 -3 3 3
use M3_M2  M3_M2_3603
timestamp 1745462530
transform 1 0 3172 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_3604
timestamp 1745462530
transform 1 0 3156 0 1 3015
box -3 -3 3 3
use M3_M2  M3_M2_3605
timestamp 1745462530
transform 1 0 3156 0 1 2925
box -3 -3 3 3
use M3_M2  M3_M2_3606
timestamp 1745462530
transform 1 0 3012 0 1 2925
box -3 -3 3 3
use M3_M2  M3_M2_3607
timestamp 1745462530
transform 1 0 2884 0 1 1615
box -3 -3 3 3
use M3_M2  M3_M2_3608
timestamp 1745462530
transform 1 0 2884 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_3609
timestamp 1745462530
transform 1 0 2788 0 1 2545
box -3 -3 3 3
use M3_M2  M3_M2_3610
timestamp 1745462530
transform 1 0 2780 0 1 2435
box -3 -3 3 3
use M3_M2  M3_M2_3611
timestamp 1745462530
transform 1 0 2772 0 1 2405
box -3 -3 3 3
use M3_M2  M3_M2_3612
timestamp 1745462530
transform 1 0 2772 0 1 1615
box -3 -3 3 3
use M3_M2  M3_M2_3613
timestamp 1745462530
transform 1 0 2764 0 1 2545
box -3 -3 3 3
use M3_M2  M3_M2_3614
timestamp 1745462530
transform 1 0 2756 0 1 2405
box -3 -3 3 3
use M3_M2  M3_M2_3615
timestamp 1745462530
transform 1 0 1644 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_3616
timestamp 1745462530
transform 1 0 1292 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_3617
timestamp 1745462530
transform 1 0 1284 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_3618
timestamp 1745462530
transform 1 0 1220 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_3619
timestamp 1745462530
transform 1 0 2844 0 1 1465
box -3 -3 3 3
use M3_M2  M3_M2_3620
timestamp 1745462530
transform 1 0 2580 0 1 1465
box -3 -3 3 3
use M3_M2  M3_M2_3621
timestamp 1745462530
transform 1 0 1948 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_3622
timestamp 1745462530
transform 1 0 1884 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_3623
timestamp 1745462530
transform 1 0 1788 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_3624
timestamp 1745462530
transform 1 0 1788 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_3625
timestamp 1745462530
transform 1 0 1772 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_3626
timestamp 1745462530
transform 1 0 1764 0 1 2415
box -3 -3 3 3
use M3_M2  M3_M2_3627
timestamp 1745462530
transform 1 0 1724 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_3628
timestamp 1745462530
transform 1 0 972 0 1 2415
box -3 -3 3 3
use M3_M2  M3_M2_3629
timestamp 1745462530
transform 1 0 588 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_3630
timestamp 1745462530
transform 1 0 580 0 1 2445
box -3 -3 3 3
use M3_M2  M3_M2_3631
timestamp 1745462530
transform 1 0 580 0 1 2415
box -3 -3 3 3
use M3_M2  M3_M2_3632
timestamp 1745462530
transform 1 0 508 0 1 2495
box -3 -3 3 3
use M3_M2  M3_M2_3633
timestamp 1745462530
transform 1 0 508 0 1 2445
box -3 -3 3 3
use M3_M2  M3_M2_3634
timestamp 1745462530
transform 1 0 372 0 1 2495
box -3 -3 3 3
use M3_M2  M3_M2_3635
timestamp 1745462530
transform 1 0 332 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_3636
timestamp 1745462530
transform 1 0 260 0 1 2495
box -3 -3 3 3
use M3_M2  M3_M2_3637
timestamp 1745462530
transform 1 0 260 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_3638
timestamp 1745462530
transform 1 0 212 0 1 2495
box -3 -3 3 3
use M3_M2  M3_M2_3639
timestamp 1745462530
transform 1 0 1780 0 1 1015
box -3 -3 3 3
use M3_M2  M3_M2_3640
timestamp 1745462530
transform 1 0 1764 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_3641
timestamp 1745462530
transform 1 0 1748 0 1 1035
box -3 -3 3 3
use M3_M2  M3_M2_3642
timestamp 1745462530
transform 1 0 1748 0 1 1015
box -3 -3 3 3
use M3_M2  M3_M2_3643
timestamp 1745462530
transform 1 0 1732 0 1 445
box -3 -3 3 3
use M3_M2  M3_M2_3644
timestamp 1745462530
transform 1 0 1716 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_3645
timestamp 1745462530
transform 1 0 1708 0 1 1035
box -3 -3 3 3
use M3_M2  M3_M2_3646
timestamp 1745462530
transform 1 0 1684 0 1 445
box -3 -3 3 3
use M3_M2  M3_M2_3647
timestamp 1745462530
transform 1 0 1660 0 1 445
box -3 -3 3 3
use M3_M2  M3_M2_3648
timestamp 1745462530
transform 1 0 1492 0 1 445
box -3 -3 3 3
use M3_M2  M3_M2_3649
timestamp 1745462530
transform 1 0 844 0 1 445
box -3 -3 3 3
use M3_M2  M3_M2_3650
timestamp 1745462530
transform 1 0 708 0 1 445
box -3 -3 3 3
use M3_M2  M3_M2_3651
timestamp 1745462530
transform 1 0 684 0 1 1335
box -3 -3 3 3
use M3_M2  M3_M2_3652
timestamp 1745462530
transform 1 0 484 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_3653
timestamp 1745462530
transform 1 0 484 0 1 1085
box -3 -3 3 3
use M3_M2  M3_M2_3654
timestamp 1745462530
transform 1 0 468 0 1 445
box -3 -3 3 3
use M3_M2  M3_M2_3655
timestamp 1745462530
transform 1 0 436 0 1 665
box -3 -3 3 3
use M3_M2  M3_M2_3656
timestamp 1745462530
transform 1 0 268 0 1 1085
box -3 -3 3 3
use M3_M2  M3_M2_3657
timestamp 1745462530
transform 1 0 244 0 1 665
box -3 -3 3 3
use M3_M2  M3_M2_3658
timestamp 1745462530
transform 1 0 3308 0 1 235
box -3 -3 3 3
use M3_M2  M3_M2_3659
timestamp 1745462530
transform 1 0 3076 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_3660
timestamp 1745462530
transform 1 0 3036 0 1 465
box -3 -3 3 3
use M3_M2  M3_M2_3661
timestamp 1745462530
transform 1 0 2932 0 1 465
box -3 -3 3 3
use M3_M2  M3_M2_3662
timestamp 1745462530
transform 1 0 2924 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_3663
timestamp 1745462530
transform 1 0 2908 0 1 465
box -3 -3 3 3
use M3_M2  M3_M2_3664
timestamp 1745462530
transform 1 0 2900 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_3665
timestamp 1745462530
transform 1 0 2844 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_3666
timestamp 1745462530
transform 1 0 2836 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_3667
timestamp 1745462530
transform 1 0 2812 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_3668
timestamp 1745462530
transform 1 0 2796 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_3669
timestamp 1745462530
transform 1 0 2580 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_3670
timestamp 1745462530
transform 1 0 1836 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_3671
timestamp 1745462530
transform 1 0 1788 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_3672
timestamp 1745462530
transform 1 0 4316 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_3673
timestamp 1745462530
transform 1 0 4308 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_3674
timestamp 1745462530
transform 1 0 4220 0 1 1975
box -3 -3 3 3
use M3_M2  M3_M2_3675
timestamp 1745462530
transform 1 0 4180 0 1 1975
box -3 -3 3 3
use M3_M2  M3_M2_3676
timestamp 1745462530
transform 1 0 4156 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_3677
timestamp 1745462530
transform 1 0 4148 0 1 1845
box -3 -3 3 3
use M3_M2  M3_M2_3678
timestamp 1745462530
transform 1 0 4148 0 1 1275
box -3 -3 3 3
use M3_M2  M3_M2_3679
timestamp 1745462530
transform 1 0 4140 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_3680
timestamp 1745462530
transform 1 0 4132 0 1 1275
box -3 -3 3 3
use M3_M2  M3_M2_3681
timestamp 1745462530
transform 1 0 4132 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_3682
timestamp 1745462530
transform 1 0 4124 0 1 255
box -3 -3 3 3
use M3_M2  M3_M2_3683
timestamp 1745462530
transform 1 0 4108 0 1 1845
box -3 -3 3 3
use M3_M2  M3_M2_3684
timestamp 1745462530
transform 1 0 4108 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_3685
timestamp 1745462530
transform 1 0 3956 0 1 255
box -3 -3 3 3
use M3_M2  M3_M2_3686
timestamp 1745462530
transform 1 0 3884 0 1 255
box -3 -3 3 3
use M3_M2  M3_M2_3687
timestamp 1745462530
transform 1 0 3876 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_3688
timestamp 1745462530
transform 1 0 3820 0 1 1975
box -3 -3 3 3
use M3_M2  M3_M2_3689
timestamp 1745462530
transform 1 0 3804 0 1 1975
box -3 -3 3 3
use M3_M2  M3_M2_3690
timestamp 1745462530
transform 1 0 4228 0 1 2665
box -3 -3 3 3
use M3_M2  M3_M2_3691
timestamp 1745462530
transform 1 0 4212 0 1 2265
box -3 -3 3 3
use M3_M2  M3_M2_3692
timestamp 1745462530
transform 1 0 4188 0 1 2735
box -3 -3 3 3
use M3_M2  M3_M2_3693
timestamp 1745462530
transform 1 0 4188 0 1 2665
box -3 -3 3 3
use M3_M2  M3_M2_3694
timestamp 1745462530
transform 1 0 4140 0 1 3015
box -3 -3 3 3
use M3_M2  M3_M2_3695
timestamp 1745462530
transform 1 0 4140 0 1 2735
box -3 -3 3 3
use M3_M2  M3_M2_3696
timestamp 1745462530
transform 1 0 4124 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_3697
timestamp 1745462530
transform 1 0 4084 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_3698
timestamp 1745462530
transform 1 0 4068 0 1 3015
box -3 -3 3 3
use M3_M2  M3_M2_3699
timestamp 1745462530
transform 1 0 3908 0 1 3025
box -3 -3 3 3
use M3_M2  M3_M2_3700
timestamp 1745462530
transform 1 0 3852 0 1 2265
box -3 -3 3 3
use M3_M2  M3_M2_3701
timestamp 1745462530
transform 1 0 3124 0 1 3025
box -3 -3 3 3
use M3_M2  M3_M2_3702
timestamp 1745462530
transform 1 0 3124 0 1 2875
box -3 -3 3 3
use M3_M2  M3_M2_3703
timestamp 1745462530
transform 1 0 3100 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_3704
timestamp 1745462530
transform 1 0 2940 0 1 2875
box -3 -3 3 3
use M3_M2  M3_M2_3705
timestamp 1745462530
transform 1 0 2940 0 1 2805
box -3 -3 3 3
use M3_M2  M3_M2_3706
timestamp 1745462530
transform 1 0 2924 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_3707
timestamp 1745462530
transform 1 0 2916 0 1 2215
box -3 -3 3 3
use M3_M2  M3_M2_3708
timestamp 1745462530
transform 1 0 2876 0 1 2805
box -3 -3 3 3
use M3_M2  M3_M2_3709
timestamp 1745462530
transform 1 0 2876 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_3710
timestamp 1745462530
transform 1 0 2772 0 1 2805
box -3 -3 3 3
use M3_M2  M3_M2_3711
timestamp 1745462530
transform 1 0 1868 0 1 2125
box -3 -3 3 3
use M3_M2  M3_M2_3712
timestamp 1745462530
transform 1 0 1852 0 1 2125
box -3 -3 3 3
use M3_M2  M3_M2_3713
timestamp 1745462530
transform 1 0 1852 0 1 2065
box -3 -3 3 3
use M3_M2  M3_M2_3714
timestamp 1745462530
transform 1 0 1772 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_3715
timestamp 1745462530
transform 1 0 1740 0 1 2065
box -3 -3 3 3
use M3_M2  M3_M2_3716
timestamp 1745462530
transform 1 0 1732 0 1 1975
box -3 -3 3 3
use M3_M2  M3_M2_3717
timestamp 1745462530
transform 1 0 3804 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_3718
timestamp 1745462530
transform 1 0 3780 0 1 1975
box -3 -3 3 3
use M3_M2  M3_M2_3719
timestamp 1745462530
transform 1 0 3764 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_3720
timestamp 1745462530
transform 1 0 3764 0 1 1975
box -3 -3 3 3
use M3_M2  M3_M2_3721
timestamp 1745462530
transform 1 0 2580 0 1 1975
box -3 -3 3 3
use M3_M2  M3_M2_3722
timestamp 1745462530
transform 1 0 2572 0 1 1875
box -3 -3 3 3
use M3_M2  M3_M2_3723
timestamp 1745462530
transform 1 0 2572 0 1 1695
box -3 -3 3 3
use M3_M2  M3_M2_3724
timestamp 1745462530
transform 1 0 2556 0 1 1435
box -3 -3 3 3
use M3_M2  M3_M2_3725
timestamp 1745462530
transform 1 0 2540 0 1 2085
box -3 -3 3 3
use M3_M2  M3_M2_3726
timestamp 1745462530
transform 1 0 2540 0 1 1875
box -3 -3 3 3
use M3_M2  M3_M2_3727
timestamp 1745462530
transform 1 0 2540 0 1 1695
box -3 -3 3 3
use M3_M2  M3_M2_3728
timestamp 1745462530
transform 1 0 2540 0 1 1435
box -3 -3 3 3
use M3_M2  M3_M2_3729
timestamp 1745462530
transform 1 0 2468 0 1 2085
box -3 -3 3 3
use M3_M2  M3_M2_3730
timestamp 1745462530
transform 1 0 3860 0 1 1055
box -3 -3 3 3
use M3_M2  M3_M2_3731
timestamp 1745462530
transform 1 0 3860 0 1 975
box -3 -3 3 3
use M3_M2  M3_M2_3732
timestamp 1745462530
transform 1 0 3836 0 1 975
box -3 -3 3 3
use M3_M2  M3_M2_3733
timestamp 1745462530
transform 1 0 3828 0 1 2245
box -3 -3 3 3
use M3_M2  M3_M2_3734
timestamp 1745462530
transform 1 0 3828 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_3735
timestamp 1745462530
transform 1 0 3828 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_3736
timestamp 1745462530
transform 1 0 3812 0 1 1615
box -3 -3 3 3
use M3_M2  M3_M2_3737
timestamp 1745462530
transform 1 0 3796 0 1 1055
box -3 -3 3 3
use M3_M2  M3_M2_3738
timestamp 1745462530
transform 1 0 3788 0 1 1645
box -3 -3 3 3
use M3_M2  M3_M2_3739
timestamp 1745462530
transform 1 0 3740 0 1 1645
box -3 -3 3 3
use M3_M2  M3_M2_3740
timestamp 1745462530
transform 1 0 3740 0 1 1615
box -3 -3 3 3
use M3_M2  M3_M2_3741
timestamp 1745462530
transform 1 0 3732 0 1 1895
box -3 -3 3 3
use M3_M2  M3_M2_3742
timestamp 1745462530
transform 1 0 3716 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_3743
timestamp 1745462530
transform 1 0 3676 0 1 2235
box -3 -3 3 3
use M3_M2  M3_M2_3744
timestamp 1745462530
transform 1 0 3652 0 1 2045
box -3 -3 3 3
use M3_M2  M3_M2_3745
timestamp 1745462530
transform 1 0 3628 0 1 2045
box -3 -3 3 3
use M3_M2  M3_M2_3746
timestamp 1745462530
transform 1 0 3628 0 1 1895
box -3 -3 3 3
use M3_M2  M3_M2_3747
timestamp 1745462530
transform 1 0 3572 0 1 2235
box -3 -3 3 3
use M3_M2  M3_M2_3748
timestamp 1745462530
transform 1 0 2428 0 1 2015
box -3 -3 3 3
use M3_M2  M3_M2_3749
timestamp 1745462530
transform 1 0 2412 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_3750
timestamp 1745462530
transform 1 0 2116 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_3751
timestamp 1745462530
transform 1 0 1932 0 1 2015
box -3 -3 3 3
use M3_M2  M3_M2_3752
timestamp 1745462530
transform 1 0 1932 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_3753
timestamp 1745462530
transform 1 0 1932 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_3754
timestamp 1745462530
transform 1 0 1932 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_3755
timestamp 1745462530
transform 1 0 1924 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_3756
timestamp 1745462530
transform 1 0 1860 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_3757
timestamp 1745462530
transform 1 0 1836 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_3758
timestamp 1745462530
transform 1 0 1532 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_3759
timestamp 1745462530
transform 1 0 1532 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_3760
timestamp 1745462530
transform 1 0 1140 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_3761
timestamp 1745462530
transform 1 0 1140 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_3762
timestamp 1745462530
transform 1 0 1028 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_3763
timestamp 1745462530
transform 1 0 996 0 1 2055
box -3 -3 3 3
use M3_M2  M3_M2_3764
timestamp 1745462530
transform 1 0 996 0 1 2015
box -3 -3 3 3
use M3_M2  M3_M2_3765
timestamp 1745462530
transform 1 0 948 0 1 2055
box -3 -3 3 3
use M3_M2  M3_M2_3766
timestamp 1745462530
transform 1 0 3388 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_3767
timestamp 1745462530
transform 1 0 3388 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_3768
timestamp 1745462530
transform 1 0 3348 0 1 2265
box -3 -3 3 3
use M3_M2  M3_M2_3769
timestamp 1745462530
transform 1 0 3340 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_3770
timestamp 1745462530
transform 1 0 3324 0 1 2265
box -3 -3 3 3
use M3_M2  M3_M2_3771
timestamp 1745462530
transform 1 0 3324 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_3772
timestamp 1745462530
transform 1 0 2812 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_3773
timestamp 1745462530
transform 1 0 2588 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_3774
timestamp 1745462530
transform 1 0 2588 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_3775
timestamp 1745462530
transform 1 0 2564 0 1 2265
box -3 -3 3 3
use M3_M2  M3_M2_3776
timestamp 1745462530
transform 1 0 2564 0 1 2205
box -3 -3 3 3
use M3_M2  M3_M2_3777
timestamp 1745462530
transform 1 0 2460 0 1 1275
box -3 -3 3 3
use M3_M2  M3_M2_3778
timestamp 1745462530
transform 1 0 2452 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_3779
timestamp 1745462530
transform 1 0 2452 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_3780
timestamp 1745462530
transform 1 0 2428 0 1 1275
box -3 -3 3 3
use M3_M2  M3_M2_3781
timestamp 1745462530
transform 1 0 2412 0 1 2205
box -3 -3 3 3
use M3_M2  M3_M2_3782
timestamp 1745462530
transform 1 0 2412 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_3783
timestamp 1745462530
transform 1 0 2348 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_3784
timestamp 1745462530
transform 1 0 2348 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_3785
timestamp 1745462530
transform 1 0 1476 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_3786
timestamp 1745462530
transform 1 0 1404 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_3787
timestamp 1745462530
transform 1 0 1404 0 1 1645
box -3 -3 3 3
use M3_M2  M3_M2_3788
timestamp 1745462530
transform 1 0 1212 0 1 1645
box -3 -3 3 3
use M3_M2  M3_M2_3789
timestamp 1745462530
transform 1 0 1204 0 1 2055
box -3 -3 3 3
use M3_M2  M3_M2_3790
timestamp 1745462530
transform 1 0 1180 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_3791
timestamp 1745462530
transform 1 0 1108 0 1 2055
box -3 -3 3 3
use M3_M2  M3_M2_3792
timestamp 1745462530
transform 1 0 1100 0 1 2185
box -3 -3 3 3
use M3_M2  M3_M2_3793
timestamp 1745462530
transform 1 0 1036 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_3794
timestamp 1745462530
transform 1 0 1028 0 1 2185
box -3 -3 3 3
use M3_M2  M3_M2_3795
timestamp 1745462530
transform 1 0 972 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_3796
timestamp 1745462530
transform 1 0 4356 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_3797
timestamp 1745462530
transform 1 0 4348 0 1 1835
box -3 -3 3 3
use M3_M2  M3_M2_3798
timestamp 1745462530
transform 1 0 4348 0 1 1005
box -3 -3 3 3
use M3_M2  M3_M2_3799
timestamp 1745462530
transform 1 0 4340 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_3800
timestamp 1745462530
transform 1 0 4116 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_3801
timestamp 1745462530
transform 1 0 4068 0 1 1005
box -3 -3 3 3
use M3_M2  M3_M2_3802
timestamp 1745462530
transform 1 0 4004 0 1 1035
box -3 -3 3 3
use M3_M2  M3_M2_3803
timestamp 1745462530
transform 1 0 4004 0 1 1005
box -3 -3 3 3
use M3_M2  M3_M2_3804
timestamp 1745462530
transform 1 0 3964 0 1 2135
box -3 -3 3 3
use M3_M2  M3_M2_3805
timestamp 1745462530
transform 1 0 3068 0 1 1035
box -3 -3 3 3
use M3_M2  M3_M2_3806
timestamp 1745462530
transform 1 0 2404 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_3807
timestamp 1745462530
transform 1 0 2076 0 1 2205
box -3 -3 3 3
use M3_M2  M3_M2_3808
timestamp 1745462530
transform 1 0 2060 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_3809
timestamp 1745462530
transform 1 0 1868 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_3810
timestamp 1745462530
transform 1 0 1868 0 1 1035
box -3 -3 3 3
use M3_M2  M3_M2_3811
timestamp 1745462530
transform 1 0 1724 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_3812
timestamp 1745462530
transform 1 0 1628 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_3813
timestamp 1745462530
transform 1 0 1628 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_3814
timestamp 1745462530
transform 1 0 932 0 1 2205
box -3 -3 3 3
use M3_M2  M3_M2_3815
timestamp 1745462530
transform 1 0 908 0 1 2205
box -3 -3 3 3
use M3_M2  M3_M2_3816
timestamp 1745462530
transform 1 0 908 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_3817
timestamp 1745462530
transform 1 0 892 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_3818
timestamp 1745462530
transform 1 0 3228 0 1 1775
box -3 -3 3 3
use M3_M2  M3_M2_3819
timestamp 1745462530
transform 1 0 3212 0 1 845
box -3 -3 3 3
use M3_M2  M3_M2_3820
timestamp 1745462530
transform 1 0 3204 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_3821
timestamp 1745462530
transform 1 0 3140 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_3822
timestamp 1745462530
transform 1 0 3132 0 1 815
box -3 -3 3 3
use M3_M2  M3_M2_3823
timestamp 1745462530
transform 1 0 3124 0 1 845
box -3 -3 3 3
use M3_M2  M3_M2_3824
timestamp 1745462530
transform 1 0 2660 0 1 1775
box -3 -3 3 3
use M3_M2  M3_M2_3825
timestamp 1745462530
transform 1 0 2660 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_3826
timestamp 1745462530
transform 1 0 2612 0 1 815
box -3 -3 3 3
use M3_M2  M3_M2_3827
timestamp 1745462530
transform 1 0 2604 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_3828
timestamp 1745462530
transform 1 0 2436 0 1 1885
box -3 -3 3 3
use M3_M2  M3_M2_3829
timestamp 1745462530
transform 1 0 2396 0 1 1885
box -3 -3 3 3
use M3_M2  M3_M2_3830
timestamp 1745462530
transform 1 0 2396 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_3831
timestamp 1745462530
transform 1 0 2340 0 1 815
box -3 -3 3 3
use M3_M2  M3_M2_3832
timestamp 1745462530
transform 1 0 1660 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_3833
timestamp 1745462530
transform 1 0 1660 0 1 1885
box -3 -3 3 3
use M3_M2  M3_M2_3834
timestamp 1745462530
transform 1 0 1428 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_3835
timestamp 1745462530
transform 1 0 1420 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_3836
timestamp 1745462530
transform 1 0 1420 0 1 1975
box -3 -3 3 3
use M3_M2  M3_M2_3837
timestamp 1745462530
transform 1 0 1372 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_3838
timestamp 1745462530
transform 1 0 1372 0 1 775
box -3 -3 3 3
use M3_M2  M3_M2_3839
timestamp 1745462530
transform 1 0 1332 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_3840
timestamp 1745462530
transform 1 0 1196 0 1 775
box -3 -3 3 3
use M3_M2  M3_M2_3841
timestamp 1745462530
transform 1 0 1196 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_3842
timestamp 1745462530
transform 1 0 1180 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_3843
timestamp 1745462530
transform 1 0 1180 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_3844
timestamp 1745462530
transform 1 0 1068 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_3845
timestamp 1745462530
transform 1 0 1068 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_3846
timestamp 1745462530
transform 1 0 1004 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_3847
timestamp 1745462530
transform 1 0 3860 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_3848
timestamp 1745462530
transform 1 0 3844 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_3849
timestamp 1745462530
transform 1 0 3836 0 1 1275
box -3 -3 3 3
use M3_M2  M3_M2_3850
timestamp 1745462530
transform 1 0 3836 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_3851
timestamp 1745462530
transform 1 0 3820 0 1 2325
box -3 -3 3 3
use M3_M2  M3_M2_3852
timestamp 1745462530
transform 1 0 3804 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_3853
timestamp 1745462530
transform 1 0 3796 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_3854
timestamp 1745462530
transform 1 0 3700 0 1 1275
box -3 -3 3 3
use M3_M2  M3_M2_3855
timestamp 1745462530
transform 1 0 3700 0 1 885
box -3 -3 3 3
use M3_M2  M3_M2_3856
timestamp 1745462530
transform 1 0 3700 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_3857
timestamp 1745462530
transform 1 0 3684 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_3858
timestamp 1745462530
transform 1 0 3564 0 1 2325
box -3 -3 3 3
use M3_M2  M3_M2_3859
timestamp 1745462530
transform 1 0 3548 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_3860
timestamp 1745462530
transform 1 0 3468 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_3861
timestamp 1745462530
transform 1 0 3468 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_3862
timestamp 1745462530
transform 1 0 2380 0 1 2045
box -3 -3 3 3
use M3_M2  M3_M2_3863
timestamp 1745462530
transform 1 0 2380 0 1 1405
box -3 -3 3 3
use M3_M2  M3_M2_3864
timestamp 1745462530
transform 1 0 2380 0 1 1265
box -3 -3 3 3
use M3_M2  M3_M2_3865
timestamp 1745462530
transform 1 0 2380 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_3866
timestamp 1745462530
transform 1 0 2364 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_3867
timestamp 1745462530
transform 1 0 2364 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_3868
timestamp 1745462530
transform 1 0 2364 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_3869
timestamp 1745462530
transform 1 0 2348 0 1 2045
box -3 -3 3 3
use M3_M2  M3_M2_3870
timestamp 1745462530
transform 1 0 2332 0 1 1405
box -3 -3 3 3
use M3_M2  M3_M2_3871
timestamp 1745462530
transform 1 0 2332 0 1 1265
box -3 -3 3 3
use M3_M2  M3_M2_3872
timestamp 1745462530
transform 1 0 2100 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_3873
timestamp 1745462530
transform 1 0 2092 0 1 845
box -3 -3 3 3
use M3_M2  M3_M2_3874
timestamp 1745462530
transform 1 0 1924 0 1 2045
box -3 -3 3 3
use M3_M2  M3_M2_3875
timestamp 1745462530
transform 1 0 1124 0 1 845
box -3 -3 3 3
use M3_M2  M3_M2_3876
timestamp 1745462530
transform 1 0 1124 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_3877
timestamp 1745462530
transform 1 0 1012 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_3878
timestamp 1745462530
transform 1 0 988 0 1 2045
box -3 -3 3 3
use M3_M2  M3_M2_3879
timestamp 1745462530
transform 1 0 980 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_3880
timestamp 1745462530
transform 1 0 940 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_3881
timestamp 1745462530
transform 1 0 3372 0 1 2205
box -3 -3 3 3
use M3_M2  M3_M2_3882
timestamp 1745462530
transform 1 0 3356 0 1 875
box -3 -3 3 3
use M3_M2  M3_M2_3883
timestamp 1745462530
transform 1 0 3300 0 1 2205
box -3 -3 3 3
use M3_M2  M3_M2_3884
timestamp 1745462530
transform 1 0 3300 0 1 2125
box -3 -3 3 3
use M3_M2  M3_M2_3885
timestamp 1745462530
transform 1 0 2788 0 1 885
box -3 -3 3 3
use M3_M2  M3_M2_3886
timestamp 1745462530
transform 1 0 2436 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_3887
timestamp 1745462530
transform 1 0 2412 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_3888
timestamp 1745462530
transform 1 0 2412 0 1 885
box -3 -3 3 3
use M3_M2  M3_M2_3889
timestamp 1745462530
transform 1 0 2372 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_3890
timestamp 1745462530
transform 1 0 1492 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_3891
timestamp 1745462530
transform 1 0 1492 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_3892
timestamp 1745462530
transform 1 0 1468 0 1 2135
box -3 -3 3 3
use M3_M2  M3_M2_3893
timestamp 1745462530
transform 1 0 1468 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_3894
timestamp 1745462530
transform 1 0 1468 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_3895
timestamp 1745462530
transform 1 0 1468 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_3896
timestamp 1745462530
transform 1 0 1468 0 1 865
box -3 -3 3 3
use M3_M2  M3_M2_3897
timestamp 1745462530
transform 1 0 1156 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_3898
timestamp 1745462530
transform 1 0 1156 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_3899
timestamp 1745462530
transform 1 0 1092 0 1 2135
box -3 -3 3 3
use M3_M2  M3_M2_3900
timestamp 1745462530
transform 1 0 1044 0 1 2205
box -3 -3 3 3
use M3_M2  M3_M2_3901
timestamp 1745462530
transform 1 0 1044 0 1 2135
box -3 -3 3 3
use M3_M2  M3_M2_3902
timestamp 1745462530
transform 1 0 1028 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_3903
timestamp 1745462530
transform 1 0 1028 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_3904
timestamp 1745462530
transform 1 0 1012 0 1 2205
box -3 -3 3 3
use M3_M2  M3_M2_3905
timestamp 1745462530
transform 1 0 924 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_3906
timestamp 1745462530
transform 1 0 4100 0 1 2185
box -3 -3 3 3
use M3_M2  M3_M2_3907
timestamp 1745462530
transform 1 0 4028 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_3908
timestamp 1745462530
transform 1 0 3988 0 1 1045
box -3 -3 3 3
use M3_M2  M3_M2_3909
timestamp 1745462530
transform 1 0 3988 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_3910
timestamp 1745462530
transform 1 0 3956 0 1 2185
box -3 -3 3 3
use M3_M2  M3_M2_3911
timestamp 1745462530
transform 1 0 3036 0 1 1045
box -3 -3 3 3
use M3_M2  M3_M2_3912
timestamp 1745462530
transform 1 0 2332 0 1 2185
box -3 -3 3 3
use M3_M2  M3_M2_3913
timestamp 1745462530
transform 1 0 2028 0 1 2185
box -3 -3 3 3
use M3_M2  M3_M2_3914
timestamp 1745462530
transform 1 0 1828 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_3915
timestamp 1745462530
transform 1 0 1676 0 1 1015
box -3 -3 3 3
use M3_M2  M3_M2_3916
timestamp 1745462530
transform 1 0 892 0 1 2175
box -3 -3 3 3
use M3_M2  M3_M2_3917
timestamp 1745462530
transform 1 0 884 0 1 1015
box -3 -3 3 3
use M3_M2  M3_M2_3918
timestamp 1745462530
transform 1 0 876 0 1 2065
box -3 -3 3 3
use M3_M2  M3_M2_3919
timestamp 1745462530
transform 1 0 876 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_3920
timestamp 1745462530
transform 1 0 868 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_3921
timestamp 1745462530
transform 1 0 844 0 1 2065
box -3 -3 3 3
use M3_M2  M3_M2_3922
timestamp 1745462530
transform 1 0 812 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_3923
timestamp 1745462530
transform 1 0 812 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_3924
timestamp 1745462530
transform 1 0 3220 0 1 1935
box -3 -3 3 3
use M3_M2  M3_M2_3925
timestamp 1745462530
transform 1 0 3172 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_3926
timestamp 1745462530
transform 1 0 3108 0 1 1875
box -3 -3 3 3
use M3_M2  M3_M2_3927
timestamp 1745462530
transform 1 0 3108 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_3928
timestamp 1745462530
transform 1 0 3084 0 1 1935
box -3 -3 3 3
use M3_M2  M3_M2_3929
timestamp 1745462530
transform 1 0 3084 0 1 1875
box -3 -3 3 3
use M3_M2  M3_M2_3930
timestamp 1745462530
transform 1 0 2332 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_3931
timestamp 1745462530
transform 1 0 2332 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_3932
timestamp 1745462530
transform 1 0 2316 0 1 1935
box -3 -3 3 3
use M3_M2  M3_M2_3933
timestamp 1745462530
transform 1 0 1692 0 1 1935
box -3 -3 3 3
use M3_M2  M3_M2_3934
timestamp 1745462530
transform 1 0 1684 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_3935
timestamp 1745462530
transform 1 0 1644 0 1 1935
box -3 -3 3 3
use M3_M2  M3_M2_3936
timestamp 1745462530
transform 1 0 1524 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_3937
timestamp 1745462530
transform 1 0 1524 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_3938
timestamp 1745462530
transform 1 0 1420 0 1 815
box -3 -3 3 3
use M3_M2  M3_M2_3939
timestamp 1745462530
transform 1 0 1364 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_3940
timestamp 1745462530
transform 1 0 1364 0 1 815
box -3 -3 3 3
use M3_M2  M3_M2_3941
timestamp 1745462530
transform 1 0 1364 0 1 675
box -3 -3 3 3
use M3_M2  M3_M2_3942
timestamp 1745462530
transform 1 0 1348 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_3943
timestamp 1745462530
transform 1 0 1316 0 1 1975
box -3 -3 3 3
use M3_M2  M3_M2_3944
timestamp 1745462530
transform 1 0 1316 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_3945
timestamp 1745462530
transform 1 0 1252 0 1 2125
box -3 -3 3 3
use M3_M2  M3_M2_3946
timestamp 1745462530
transform 1 0 1252 0 1 1975
box -3 -3 3 3
use M3_M2  M3_M2_3947
timestamp 1745462530
transform 1 0 1060 0 1 2125
box -3 -3 3 3
use M3_M2  M3_M2_3948
timestamp 1745462530
transform 1 0 1020 0 1 675
box -3 -3 3 3
use M3_M2  M3_M2_3949
timestamp 1745462530
transform 1 0 988 0 1 675
box -3 -3 3 3
use M3_M2  M3_M2_3950
timestamp 1745462530
transform 1 0 3660 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_3951
timestamp 1745462530
transform 1 0 3548 0 1 1265
box -3 -3 3 3
use M3_M2  M3_M2_3952
timestamp 1745462530
transform 1 0 3548 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_3953
timestamp 1745462530
transform 1 0 3068 0 1 2255
box -3 -3 3 3
use M3_M2  M3_M2_3954
timestamp 1745462530
transform 1 0 2636 0 1 1685
box -3 -3 3 3
use M3_M2  M3_M2_3955
timestamp 1745462530
transform 1 0 2524 0 1 2245
box -3 -3 3 3
use M3_M2  M3_M2_3956
timestamp 1745462530
transform 1 0 2524 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_3957
timestamp 1745462530
transform 1 0 2524 0 1 1685
box -3 -3 3 3
use M3_M2  M3_M2_3958
timestamp 1745462530
transform 1 0 2516 0 1 1285
box -3 -3 3 3
use M3_M2  M3_M2_3959
timestamp 1745462530
transform 1 0 2092 0 1 1285
box -3 -3 3 3
use M3_M2  M3_M2_3960
timestamp 1745462530
transform 1 0 2068 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_3961
timestamp 1745462530
transform 1 0 2068 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_3962
timestamp 1745462530
transform 1 0 1940 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_3963
timestamp 1745462530
transform 1 0 1220 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_3964
timestamp 1745462530
transform 1 0 1036 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_3965
timestamp 1745462530
transform 1 0 1028 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_3966
timestamp 1745462530
transform 1 0 1028 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_3967
timestamp 1745462530
transform 1 0 924 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_3968
timestamp 1745462530
transform 1 0 924 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_3969
timestamp 1745462530
transform 1 0 876 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_3970
timestamp 1745462530
transform 1 0 3308 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_3971
timestamp 1745462530
transform 1 0 2892 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_3972
timestamp 1745462530
transform 1 0 2836 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_3973
timestamp 1745462530
transform 1 0 2836 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_3974
timestamp 1745462530
transform 1 0 2756 0 1 2065
box -3 -3 3 3
use M3_M2  M3_M2_3975
timestamp 1745462530
transform 1 0 2756 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_3976
timestamp 1745462530
transform 1 0 2732 0 1 2165
box -3 -3 3 3
use M3_M2  M3_M2_3977
timestamp 1745462530
transform 1 0 2732 0 1 2065
box -3 -3 3 3
use M3_M2  M3_M2_3978
timestamp 1745462530
transform 1 0 2716 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_3979
timestamp 1745462530
transform 1 0 2516 0 1 2165
box -3 -3 3 3
use M3_M2  M3_M2_3980
timestamp 1745462530
transform 1 0 2476 0 1 1695
box -3 -3 3 3
use M3_M2  M3_M2_3981
timestamp 1745462530
transform 1 0 2460 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_3982
timestamp 1745462530
transform 1 0 1332 0 1 1695
box -3 -3 3 3
use M3_M2  M3_M2_3983
timestamp 1745462530
transform 1 0 1316 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_3984
timestamp 1745462530
transform 1 0 1260 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_3985
timestamp 1745462530
transform 1 0 1260 0 1 1495
box -3 -3 3 3
use M3_M2  M3_M2_3986
timestamp 1745462530
transform 1 0 1220 0 1 1495
box -3 -3 3 3
use M3_M2  M3_M2_3987
timestamp 1745462530
transform 1 0 1220 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_3988
timestamp 1745462530
transform 1 0 1164 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_3989
timestamp 1745462530
transform 1 0 1164 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_3990
timestamp 1745462530
transform 1 0 1116 0 1 1495
box -3 -3 3 3
use M3_M2  M3_M2_3991
timestamp 1745462530
transform 1 0 1084 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_3992
timestamp 1745462530
transform 1 0 1084 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_3993
timestamp 1745462530
transform 1 0 1084 0 1 1495
box -3 -3 3 3
use M3_M2  M3_M2_3994
timestamp 1745462530
transform 1 0 996 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_3995
timestamp 1745462530
transform 1 0 3860 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_3996
timestamp 1745462530
transform 1 0 3116 0 1 1465
box -3 -3 3 3
use M3_M2  M3_M2_3997
timestamp 1745462530
transform 1 0 3108 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_3998
timestamp 1745462530
transform 1 0 3108 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_3999
timestamp 1745462530
transform 1 0 3100 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_4000
timestamp 1745462530
transform 1 0 3100 0 1 1465
box -3 -3 3 3
use M3_M2  M3_M2_4001
timestamp 1745462530
transform 1 0 3076 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_4002
timestamp 1745462530
transform 1 0 3028 0 1 2275
box -3 -3 3 3
use M3_M2  M3_M2_4003
timestamp 1745462530
transform 1 0 2980 0 1 2275
box -3 -3 3 3
use M3_M2  M3_M2_4004
timestamp 1745462530
transform 1 0 2884 0 1 1415
box -3 -3 3 3
use M3_M2  M3_M2_4005
timestamp 1745462530
transform 1 0 2884 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_4006
timestamp 1745462530
transform 1 0 2484 0 1 2095
box -3 -3 3 3
use M3_M2  M3_M2_4007
timestamp 1745462530
transform 1 0 2332 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_4008
timestamp 1745462530
transform 1 0 2324 0 1 1435
box -3 -3 3 3
use M3_M2  M3_M2_4009
timestamp 1745462530
transform 1 0 2268 0 1 2095
box -3 -3 3 3
use M3_M2  M3_M2_4010
timestamp 1745462530
transform 1 0 2268 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_4011
timestamp 1745462530
transform 1 0 2220 0 1 1895
box -3 -3 3 3
use M3_M2  M3_M2_4012
timestamp 1745462530
transform 1 0 2220 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_4013
timestamp 1745462530
transform 1 0 2180 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_4014
timestamp 1745462530
transform 1 0 2180 0 1 1895
box -3 -3 3 3
use M3_M2  M3_M2_4015
timestamp 1745462530
transform 1 0 2012 0 1 1895
box -3 -3 3 3
use M3_M2  M3_M2_4016
timestamp 1745462530
transform 1 0 2012 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_4017
timestamp 1745462530
transform 1 0 1940 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_4018
timestamp 1745462530
transform 1 0 1900 0 1 1435
box -3 -3 3 3
use M3_M2  M3_M2_4019
timestamp 1745462530
transform 1 0 1692 0 1 1435
box -3 -3 3 3
use M3_M2  M3_M2_4020
timestamp 1745462530
transform 1 0 988 0 1 1885
box -3 -3 3 3
use M3_M2  M3_M2_4021
timestamp 1745462530
transform 1 0 932 0 1 1435
box -3 -3 3 3
use M3_M2  M3_M2_4022
timestamp 1745462530
transform 1 0 924 0 1 1885
box -3 -3 3 3
use M3_M2  M3_M2_4023
timestamp 1745462530
transform 1 0 924 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_4024
timestamp 1745462530
transform 1 0 924 0 1 1655
box -3 -3 3 3
use M3_M2  M3_M2_4025
timestamp 1745462530
transform 1 0 868 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_4026
timestamp 1745462530
transform 1 0 868 0 1 1655
box -3 -3 3 3
use M3_M2  M3_M2_4027
timestamp 1745462530
transform 1 0 3092 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_4028
timestamp 1745462530
transform 1 0 2980 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_4029
timestamp 1745462530
transform 1 0 2940 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_4030
timestamp 1745462530
transform 1 0 2876 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_4031
timestamp 1745462530
transform 1 0 2732 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_4032
timestamp 1745462530
transform 1 0 2620 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_4033
timestamp 1745462530
transform 1 0 2612 0 1 1615
box -3 -3 3 3
use M3_M2  M3_M2_4034
timestamp 1745462530
transform 1 0 2580 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_4035
timestamp 1745462530
transform 1 0 2580 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_4036
timestamp 1745462530
transform 1 0 2508 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_4037
timestamp 1745462530
transform 1 0 2508 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_4038
timestamp 1745462530
transform 1 0 2420 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_4039
timestamp 1745462530
transform 1 0 2420 0 1 1475
box -3 -3 3 3
use M3_M2  M3_M2_4040
timestamp 1745462530
transform 1 0 2332 0 1 1475
box -3 -3 3 3
use M3_M2  M3_M2_4041
timestamp 1745462530
transform 1 0 1516 0 1 1475
box -3 -3 3 3
use M3_M2  M3_M2_4042
timestamp 1745462530
transform 1 0 1492 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_4043
timestamp 1745462530
transform 1 0 1252 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_4044
timestamp 1745462530
transform 1 0 1044 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_4045
timestamp 1745462530
transform 1 0 1044 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_4046
timestamp 1745462530
transform 1 0 1028 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_4047
timestamp 1745462530
transform 1 0 996 0 1 1495
box -3 -3 3 3
use M3_M2  M3_M2_4048
timestamp 1745462530
transform 1 0 964 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_4049
timestamp 1745462530
transform 1 0 956 0 1 1495
box -3 -3 3 3
use M3_M2  M3_M2_4050
timestamp 1745462530
transform 1 0 4372 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_4051
timestamp 1745462530
transform 1 0 4364 0 1 2645
box -3 -3 3 3
use M3_M2  M3_M2_4052
timestamp 1745462530
transform 1 0 4364 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_4053
timestamp 1745462530
transform 1 0 4356 0 1 1375
box -3 -3 3 3
use M3_M2  M3_M2_4054
timestamp 1745462530
transform 1 0 3972 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_4055
timestamp 1745462530
transform 1 0 3964 0 1 1375
box -3 -3 3 3
use M3_M2  M3_M2_4056
timestamp 1745462530
transform 1 0 3916 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_4057
timestamp 1745462530
transform 1 0 3916 0 1 1075
box -3 -3 3 3
use M3_M2  M3_M2_4058
timestamp 1745462530
transform 1 0 3900 0 1 1075
box -3 -3 3 3
use M3_M2  M3_M2_4059
timestamp 1745462530
transform 1 0 3900 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_4060
timestamp 1745462530
transform 1 0 3868 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_4061
timestamp 1745462530
transform 1 0 3868 0 1 775
box -3 -3 3 3
use M3_M2  M3_M2_4062
timestamp 1745462530
transform 1 0 3812 0 1 2645
box -3 -3 3 3
use M3_M2  M3_M2_4063
timestamp 1745462530
transform 1 0 3796 0 1 2715
box -3 -3 3 3
use M3_M2  M3_M2_4064
timestamp 1745462530
transform 1 0 3772 0 1 1375
box -3 -3 3 3
use M3_M2  M3_M2_4065
timestamp 1745462530
transform 1 0 3708 0 1 775
box -3 -3 3 3
use M3_M2  M3_M2_4066
timestamp 1745462530
transform 1 0 3708 0 1 685
box -3 -3 3 3
use M3_M2  M3_M2_4067
timestamp 1745462530
transform 1 0 3668 0 1 2765
box -3 -3 3 3
use M3_M2  M3_M2_4068
timestamp 1745462530
transform 1 0 3668 0 1 2715
box -3 -3 3 3
use M3_M2  M3_M2_4069
timestamp 1745462530
transform 1 0 3668 0 1 2665
box -3 -3 3 3
use M3_M2  M3_M2_4070
timestamp 1745462530
transform 1 0 3652 0 1 685
box -3 -3 3 3
use M3_M2  M3_M2_4071
timestamp 1745462530
transform 1 0 3612 0 1 2665
box -3 -3 3 3
use M3_M2  M3_M2_4072
timestamp 1745462530
transform 1 0 3492 0 1 685
box -3 -3 3 3
use M3_M2  M3_M2_4073
timestamp 1745462530
transform 1 0 3484 0 1 265
box -3 -3 3 3
use M3_M2  M3_M2_4074
timestamp 1745462530
transform 1 0 2564 0 1 2765
box -3 -3 3 3
use M3_M2  M3_M2_4075
timestamp 1745462530
transform 1 0 2556 0 1 445
box -3 -3 3 3
use M3_M2  M3_M2_4076
timestamp 1745462530
transform 1 0 2540 0 1 265
box -3 -3 3 3
use M3_M2  M3_M2_4077
timestamp 1745462530
transform 1 0 2540 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_4078
timestamp 1745462530
transform 1 0 2532 0 1 445
box -3 -3 3 3
use M3_M2  M3_M2_4079
timestamp 1745462530
transform 1 0 2028 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_4080
timestamp 1745462530
transform 1 0 2028 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_4081
timestamp 1745462530
transform 1 0 1852 0 1 2765
box -3 -3 3 3
use M3_M2  M3_M2_4082
timestamp 1745462530
transform 1 0 1092 0 1 605
box -3 -3 3 3
use M3_M2  M3_M2_4083
timestamp 1745462530
transform 1 0 1028 0 1 2765
box -3 -3 3 3
use M3_M2  M3_M2_4084
timestamp 1745462530
transform 1 0 1028 0 1 2645
box -3 -3 3 3
use M3_M2  M3_M2_4085
timestamp 1745462530
transform 1 0 932 0 1 675
box -3 -3 3 3
use M3_M2  M3_M2_4086
timestamp 1745462530
transform 1 0 932 0 1 605
box -3 -3 3 3
use M3_M2  M3_M2_4087
timestamp 1745462530
transform 1 0 820 0 1 2685
box -3 -3 3 3
use M3_M2  M3_M2_4088
timestamp 1745462530
transform 1 0 820 0 1 2655
box -3 -3 3 3
use M3_M2  M3_M2_4089
timestamp 1745462530
transform 1 0 804 0 1 675
box -3 -3 3 3
use M3_M2  M3_M2_4090
timestamp 1745462530
transform 1 0 788 0 1 2685
box -3 -3 3 3
use M3_M2  M3_M2_4091
timestamp 1745462530
transform 1 0 3596 0 1 2665
box -3 -3 3 3
use M3_M2  M3_M2_4092
timestamp 1745462530
transform 1 0 3580 0 1 655
box -3 -3 3 3
use M3_M2  M3_M2_4093
timestamp 1745462530
transform 1 0 3548 0 1 2665
box -3 -3 3 3
use M3_M2  M3_M2_4094
timestamp 1745462530
transform 1 0 3476 0 1 655
box -3 -3 3 3
use M3_M2  M3_M2_4095
timestamp 1745462530
transform 1 0 3476 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_4096
timestamp 1745462530
transform 1 0 3460 0 1 655
box -3 -3 3 3
use M3_M2  M3_M2_4097
timestamp 1745462530
transform 1 0 2708 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_4098
timestamp 1745462530
transform 1 0 2588 0 1 2685
box -3 -3 3 3
use M3_M2  M3_M2_4099
timestamp 1745462530
transform 1 0 2588 0 1 2665
box -3 -3 3 3
use M3_M2  M3_M2_4100
timestamp 1745462530
transform 1 0 2428 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_4101
timestamp 1745462530
transform 1 0 2404 0 1 675
box -3 -3 3 3
use M3_M2  M3_M2_4102
timestamp 1745462530
transform 1 0 2244 0 1 675
box -3 -3 3 3
use M3_M2  M3_M2_4103
timestamp 1745462530
transform 1 0 2244 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_4104
timestamp 1745462530
transform 1 0 2180 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_4105
timestamp 1745462530
transform 1 0 2180 0 1 65
box -3 -3 3 3
use M3_M2  M3_M2_4106
timestamp 1745462530
transform 1 0 1604 0 1 455
box -3 -3 3 3
use M3_M2  M3_M2_4107
timestamp 1745462530
transform 1 0 1604 0 1 65
box -3 -3 3 3
use M3_M2  M3_M2_4108
timestamp 1745462530
transform 1 0 1556 0 1 2685
box -3 -3 3 3
use M3_M2  M3_M2_4109
timestamp 1745462530
transform 1 0 1548 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_4110
timestamp 1745462530
transform 1 0 1444 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_4111
timestamp 1745462530
transform 1 0 1444 0 1 2785
box -3 -3 3 3
use M3_M2  M3_M2_4112
timestamp 1745462530
transform 1 0 1236 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_4113
timestamp 1745462530
transform 1 0 1236 0 1 455
box -3 -3 3 3
use M3_M2  M3_M2_4114
timestamp 1745462530
transform 1 0 1212 0 1 2785
box -3 -3 3 3
use M3_M2  M3_M2_4115
timestamp 1745462530
transform 1 0 1180 0 1 775
box -3 -3 3 3
use M3_M2  M3_M2_4116
timestamp 1745462530
transform 1 0 1172 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_4117
timestamp 1745462530
transform 1 0 1156 0 1 815
box -3 -3 3 3
use M3_M2  M3_M2_4118
timestamp 1745462530
transform 1 0 1156 0 1 775
box -3 -3 3 3
use M3_M2  M3_M2_4119
timestamp 1745462530
transform 1 0 1124 0 1 2785
box -3 -3 3 3
use M3_M2  M3_M2_4120
timestamp 1745462530
transform 1 0 1124 0 1 2685
box -3 -3 3 3
use M3_M2  M3_M2_4121
timestamp 1745462530
transform 1 0 876 0 1 2685
box -3 -3 3 3
use M3_M2  M3_M2_4122
timestamp 1745462530
transform 1 0 756 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_4123
timestamp 1745462530
transform 1 0 756 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_4124
timestamp 1745462530
transform 1 0 644 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_4125
timestamp 1745462530
transform 1 0 580 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_4126
timestamp 1745462530
transform 1 0 4148 0 1 2555
box -3 -3 3 3
use M3_M2  M3_M2_4127
timestamp 1745462530
transform 1 0 4036 0 1 2585
box -3 -3 3 3
use M3_M2  M3_M2_4128
timestamp 1745462530
transform 1 0 4036 0 1 2555
box -3 -3 3 3
use M3_M2  M3_M2_4129
timestamp 1745462530
transform 1 0 3940 0 1 535
box -3 -3 3 3
use M3_M2  M3_M2_4130
timestamp 1745462530
transform 1 0 3876 0 1 665
box -3 -3 3 3
use M3_M2  M3_M2_4131
timestamp 1745462530
transform 1 0 3876 0 1 535
box -3 -3 3 3
use M3_M2  M3_M2_4132
timestamp 1745462530
transform 1 0 3100 0 1 295
box -3 -3 3 3
use M3_M2  M3_M2_4133
timestamp 1745462530
transform 1 0 3084 0 1 655
box -3 -3 3 3
use M3_M2  M3_M2_4134
timestamp 1745462530
transform 1 0 2988 0 1 655
box -3 -3 3 3
use M3_M2  M3_M2_4135
timestamp 1745462530
transform 1 0 2652 0 1 2585
box -3 -3 3 3
use M3_M2  M3_M2_4136
timestamp 1745462530
transform 1 0 2004 0 1 2585
box -3 -3 3 3
use M3_M2  M3_M2_4137
timestamp 1745462530
transform 1 0 1996 0 1 2665
box -3 -3 3 3
use M3_M2  M3_M2_4138
timestamp 1745462530
transform 1 0 1812 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_4139
timestamp 1745462530
transform 1 0 1812 0 1 295
box -3 -3 3 3
use M3_M2  M3_M2_4140
timestamp 1745462530
transform 1 0 1796 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_4141
timestamp 1745462530
transform 1 0 1796 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_4142
timestamp 1745462530
transform 1 0 1772 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_4143
timestamp 1745462530
transform 1 0 1652 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_4144
timestamp 1745462530
transform 1 0 1420 0 1 575
box -3 -3 3 3
use M3_M2  M3_M2_4145
timestamp 1745462530
transform 1 0 1420 0 1 415
box -3 -3 3 3
use M3_M2  M3_M2_4146
timestamp 1745462530
transform 1 0 684 0 1 665
box -3 -3 3 3
use M3_M2  M3_M2_4147
timestamp 1745462530
transform 1 0 684 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_4148
timestamp 1745462530
transform 1 0 668 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_4149
timestamp 1745462530
transform 1 0 668 0 1 665
box -3 -3 3 3
use M3_M2  M3_M2_4150
timestamp 1745462530
transform 1 0 652 0 1 2565
box -3 -3 3 3
use M3_M2  M3_M2_4151
timestamp 1745462530
transform 1 0 620 0 1 2565
box -3 -3 3 3
use M3_M2  M3_M2_4152
timestamp 1745462530
transform 1 0 612 0 1 2655
box -3 -3 3 3
use M3_M2  M3_M2_4153
timestamp 1745462530
transform 1 0 604 0 1 875
box -3 -3 3 3
use M3_M2  M3_M2_4154
timestamp 1745462530
transform 1 0 604 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_4155
timestamp 1745462530
transform 1 0 188 0 1 2655
box -3 -3 3 3
use M3_M2  M3_M2_4156
timestamp 1745462530
transform 1 0 188 0 1 1835
box -3 -3 3 3
use M3_M2  M3_M2_4157
timestamp 1745462530
transform 1 0 188 0 1 1775
box -3 -3 3 3
use M3_M2  M3_M2_4158
timestamp 1745462530
transform 1 0 188 0 1 875
box -3 -3 3 3
use M3_M2  M3_M2_4159
timestamp 1745462530
transform 1 0 148 0 1 1835
box -3 -3 3 3
use M3_M2  M3_M2_4160
timestamp 1745462530
transform 1 0 148 0 1 1775
box -3 -3 3 3
use M3_M2  M3_M2_4161
timestamp 1745462530
transform 1 0 3460 0 1 1415
box -3 -3 3 3
use M3_M2  M3_M2_4162
timestamp 1745462530
transform 1 0 3372 0 1 1415
box -3 -3 3 3
use M3_M2  M3_M2_4163
timestamp 1745462530
transform 1 0 3372 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_4164
timestamp 1745462530
transform 1 0 3372 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_4165
timestamp 1745462530
transform 1 0 3364 0 1 2605
box -3 -3 3 3
use M3_M2  M3_M2_4166
timestamp 1745462530
transform 1 0 3364 0 1 1875
box -3 -3 3 3
use M3_M2  M3_M2_4167
timestamp 1745462530
transform 1 0 3356 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_4168
timestamp 1745462530
transform 1 0 3356 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_4169
timestamp 1745462530
transform 1 0 3348 0 1 1875
box -3 -3 3 3
use M3_M2  M3_M2_4170
timestamp 1745462530
transform 1 0 3340 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_4171
timestamp 1745462530
transform 1 0 3252 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_4172
timestamp 1745462530
transform 1 0 3244 0 1 2625
box -3 -3 3 3
use M3_M2  M3_M2_4173
timestamp 1745462530
transform 1 0 3244 0 1 2605
box -3 -3 3 3
use M3_M2  M3_M2_4174
timestamp 1745462530
transform 1 0 3236 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_4175
timestamp 1745462530
transform 1 0 2924 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_4176
timestamp 1745462530
transform 1 0 2924 0 1 495
box -3 -3 3 3
use M3_M2  M3_M2_4177
timestamp 1745462530
transform 1 0 2628 0 1 2625
box -3 -3 3 3
use M3_M2  M3_M2_4178
timestamp 1745462530
transform 1 0 2508 0 1 2785
box -3 -3 3 3
use M3_M2  M3_M2_4179
timestamp 1745462530
transform 1 0 2508 0 1 2625
box -3 -3 3 3
use M3_M2  M3_M2_4180
timestamp 1745462530
transform 1 0 2252 0 1 575
box -3 -3 3 3
use M3_M2  M3_M2_4181
timestamp 1745462530
transform 1 0 1700 0 1 2815
box -3 -3 3 3
use M3_M2  M3_M2_4182
timestamp 1745462530
transform 1 0 1700 0 1 2785
box -3 -3 3 3
use M3_M2  M3_M2_4183
timestamp 1745462530
transform 1 0 1396 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_4184
timestamp 1745462530
transform 1 0 1364 0 1 2815
box -3 -3 3 3
use M3_M2  M3_M2_4185
timestamp 1745462530
transform 1 0 628 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_4186
timestamp 1745462530
transform 1 0 612 0 1 2805
box -3 -3 3 3
use M3_M2  M3_M2_4187
timestamp 1745462530
transform 1 0 612 0 1 725
box -3 -3 3 3
use M3_M2  M3_M2_4188
timestamp 1745462530
transform 1 0 532 0 1 725
box -3 -3 3 3
use M3_M2  M3_M2_4189
timestamp 1745462530
transform 1 0 3796 0 1 2645
box -3 -3 3 3
use M3_M2  M3_M2_4190
timestamp 1745462530
transform 1 0 3756 0 1 2745
box -3 -3 3 3
use M3_M2  M3_M2_4191
timestamp 1745462530
transform 1 0 3756 0 1 2645
box -3 -3 3 3
use M3_M2  M3_M2_4192
timestamp 1745462530
transform 1 0 3756 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_4193
timestamp 1745462530
transform 1 0 3692 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_4194
timestamp 1745462530
transform 1 0 3676 0 1 645
box -3 -3 3 3
use M3_M2  M3_M2_4195
timestamp 1745462530
transform 1 0 3404 0 1 645
box -3 -3 3 3
use M3_M2  M3_M2_4196
timestamp 1745462530
transform 1 0 3404 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_4197
timestamp 1745462530
transform 1 0 3324 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_4198
timestamp 1745462530
transform 1 0 3324 0 1 405
box -3 -3 3 3
use M3_M2  M3_M2_4199
timestamp 1745462530
transform 1 0 2876 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_4200
timestamp 1745462530
transform 1 0 2876 0 1 405
box -3 -3 3 3
use M3_M2  M3_M2_4201
timestamp 1745462530
transform 1 0 2812 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_4202
timestamp 1745462530
transform 1 0 2812 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_4203
timestamp 1745462530
transform 1 0 2596 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_4204
timestamp 1745462530
transform 1 0 2596 0 1 535
box -3 -3 3 3
use M3_M2  M3_M2_4205
timestamp 1745462530
transform 1 0 2524 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_4206
timestamp 1745462530
transform 1 0 2500 0 1 2745
box -3 -3 3 3
use M3_M2  M3_M2_4207
timestamp 1745462530
transform 1 0 2156 0 1 655
box -3 -3 3 3
use M3_M2  M3_M2_4208
timestamp 1745462530
transform 1 0 2156 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_4209
timestamp 1745462530
transform 1 0 1988 0 1 655
box -3 -3 3 3
use M3_M2  M3_M2_4210
timestamp 1745462530
transform 1 0 1820 0 1 2745
box -3 -3 3 3
use M3_M2  M3_M2_4211
timestamp 1745462530
transform 1 0 1060 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_4212
timestamp 1745462530
transform 1 0 852 0 1 685
box -3 -3 3 3
use M3_M2  M3_M2_4213
timestamp 1745462530
transform 1 0 852 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_4214
timestamp 1745462530
transform 1 0 788 0 1 2745
box -3 -3 3 3
use M3_M2  M3_M2_4215
timestamp 1745462530
transform 1 0 772 0 1 685
box -3 -3 3 3
use M3_M2  M3_M2_4216
timestamp 1745462530
transform 1 0 3628 0 1 1885
box -3 -3 3 3
use M3_M2  M3_M2_4217
timestamp 1745462530
transform 1 0 3628 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_4218
timestamp 1745462530
transform 1 0 3628 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_4219
timestamp 1745462530
transform 1 0 3596 0 1 1085
box -3 -3 3 3
use M3_M2  M3_M2_4220
timestamp 1745462530
transform 1 0 3596 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_4221
timestamp 1745462530
transform 1 0 3588 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_4222
timestamp 1745462530
transform 1 0 3580 0 1 1885
box -3 -3 3 3
use M3_M2  M3_M2_4223
timestamp 1745462530
transform 1 0 3548 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_4224
timestamp 1745462530
transform 1 0 3548 0 1 1085
box -3 -3 3 3
use M3_M2  M3_M2_4225
timestamp 1745462530
transform 1 0 3524 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_4226
timestamp 1745462530
transform 1 0 3516 0 1 2685
box -3 -3 3 3
use M3_M2  M3_M2_4227
timestamp 1745462530
transform 1 0 3476 0 1 2815
box -3 -3 3 3
use M3_M2  M3_M2_4228
timestamp 1745462530
transform 1 0 3476 0 1 2685
box -3 -3 3 3
use M3_M2  M3_M2_4229
timestamp 1745462530
transform 1 0 3428 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_4230
timestamp 1745462530
transform 1 0 2724 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_4231
timestamp 1745462530
transform 1 0 2692 0 1 465
box -3 -3 3 3
use M3_M2  M3_M2_4232
timestamp 1745462530
transform 1 0 2476 0 1 2805
box -3 -3 3 3
use M3_M2  M3_M2_4233
timestamp 1745462530
transform 1 0 1500 0 1 2875
box -3 -3 3 3
use M3_M2  M3_M2_4234
timestamp 1745462530
transform 1 0 1500 0 1 2805
box -3 -3 3 3
use M3_M2  M3_M2_4235
timestamp 1745462530
transform 1 0 1300 0 1 2875
box -3 -3 3 3
use M3_M2  M3_M2_4236
timestamp 1745462530
transform 1 0 1276 0 1 2845
box -3 -3 3 3
use M3_M2  M3_M2_4237
timestamp 1745462530
transform 1 0 1180 0 1 2845
box -3 -3 3 3
use M3_M2  M3_M2_4238
timestamp 1745462530
transform 1 0 1180 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_4239
timestamp 1745462530
transform 1 0 1132 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_4240
timestamp 1745462530
transform 1 0 1108 0 1 655
box -3 -3 3 3
use M3_M2  M3_M2_4241
timestamp 1745462530
transform 1 0 972 0 1 865
box -3 -3 3 3
use M3_M2  M3_M2_4242
timestamp 1745462530
transform 1 0 972 0 1 655
box -3 -3 3 3
use M3_M2  M3_M2_4243
timestamp 1745462530
transform 1 0 836 0 1 2775
box -3 -3 3 3
use M3_M2  M3_M2_4244
timestamp 1745462530
transform 1 0 748 0 1 2775
box -3 -3 3 3
use M3_M2  M3_M2_4245
timestamp 1745462530
transform 1 0 612 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_4246
timestamp 1745462530
transform 1 0 548 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_4247
timestamp 1745462530
transform 1 0 548 0 1 865
box -3 -3 3 3
use M3_M2  M3_M2_4248
timestamp 1745462530
transform 1 0 4108 0 1 2635
box -3 -3 3 3
use M3_M2  M3_M2_4249
timestamp 1745462530
transform 1 0 4100 0 1 2585
box -3 -3 3 3
use M3_M2  M3_M2_4250
timestamp 1745462530
transform 1 0 4036 0 1 2385
box -3 -3 3 3
use M3_M2  M3_M2_4251
timestamp 1745462530
transform 1 0 4028 0 1 2575
box -3 -3 3 3
use M3_M2  M3_M2_4252
timestamp 1745462530
transform 1 0 4020 0 1 2385
box -3 -3 3 3
use M3_M2  M3_M2_4253
timestamp 1745462530
transform 1 0 4020 0 1 2055
box -3 -3 3 3
use M3_M2  M3_M2_4254
timestamp 1745462530
transform 1 0 3908 0 1 475
box -3 -3 3 3
use M3_M2  M3_M2_4255
timestamp 1745462530
transform 1 0 3572 0 1 2055
box -3 -3 3 3
use M3_M2  M3_M2_4256
timestamp 1745462530
transform 1 0 2956 0 1 685
box -3 -3 3 3
use M3_M2  M3_M2_4257
timestamp 1745462530
transform 1 0 2868 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_4258
timestamp 1745462530
transform 1 0 2868 0 1 475
box -3 -3 3 3
use M3_M2  M3_M2_4259
timestamp 1745462530
transform 1 0 2828 0 1 685
box -3 -3 3 3
use M3_M2  M3_M2_4260
timestamp 1745462530
transform 1 0 2828 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_4261
timestamp 1745462530
transform 1 0 2780 0 1 685
box -3 -3 3 3
use M3_M2  M3_M2_4262
timestamp 1745462530
transform 1 0 2748 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_4263
timestamp 1745462530
transform 1 0 2580 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_4264
timestamp 1745462530
transform 1 0 2580 0 1 645
box -3 -3 3 3
use M3_M2  M3_M2_4265
timestamp 1745462530
transform 1 0 2532 0 1 2635
box -3 -3 3 3
use M3_M2  M3_M2_4266
timestamp 1745462530
transform 1 0 2356 0 1 645
box -3 -3 3 3
use M3_M2  M3_M2_4267
timestamp 1745462530
transform 1 0 1956 0 1 2615
box -3 -3 3 3
use M3_M2  M3_M2_4268
timestamp 1745462530
transform 1 0 1820 0 1 675
box -3 -3 3 3
use M3_M2  M3_M2_4269
timestamp 1745462530
transform 1 0 1820 0 1 645
box -3 -3 3 3
use M3_M2  M3_M2_4270
timestamp 1745462530
transform 1 0 1748 0 1 675
box -3 -3 3 3
use M3_M2  M3_M2_4271
timestamp 1745462530
transform 1 0 1748 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_4272
timestamp 1745462530
transform 1 0 1628 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_4273
timestamp 1745462530
transform 1 0 1596 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_4274
timestamp 1745462530
transform 1 0 796 0 1 655
box -3 -3 3 3
use M3_M2  M3_M2_4275
timestamp 1745462530
transform 1 0 796 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_4276
timestamp 1745462530
transform 1 0 780 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_4277
timestamp 1745462530
transform 1 0 780 0 1 655
box -3 -3 3 3
use M3_M2  M3_M2_4278
timestamp 1745462530
transform 1 0 604 0 1 2615
box -3 -3 3 3
use M3_M2  M3_M2_4279
timestamp 1745462530
transform 1 0 604 0 1 2565
box -3 -3 3 3
use M3_M2  M3_M2_4280
timestamp 1745462530
transform 1 0 588 0 1 2615
box -3 -3 3 3
use M3_M2  M3_M2_4281
timestamp 1745462530
transform 1 0 588 0 1 2565
box -3 -3 3 3
use M3_M2  M3_M2_4282
timestamp 1745462530
transform 1 0 580 0 1 2685
box -3 -3 3 3
use M3_M2  M3_M2_4283
timestamp 1745462530
transform 1 0 572 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_4284
timestamp 1745462530
transform 1 0 68 0 1 2685
box -3 -3 3 3
use M3_M2  M3_M2_4285
timestamp 1745462530
transform 1 0 68 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_4286
timestamp 1745462530
transform 1 0 3860 0 1 375
box -3 -3 3 3
use M3_M2  M3_M2_4287
timestamp 1745462530
transform 1 0 3492 0 1 1215
box -3 -3 3 3
use M3_M2  M3_M2_4288
timestamp 1745462530
transform 1 0 3492 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_4289
timestamp 1745462530
transform 1 0 3444 0 1 1275
box -3 -3 3 3
use M3_M2  M3_M2_4290
timestamp 1745462530
transform 1 0 3444 0 1 1215
box -3 -3 3 3
use M3_M2  M3_M2_4291
timestamp 1745462530
transform 1 0 3444 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_4292
timestamp 1745462530
transform 1 0 3444 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_4293
timestamp 1745462530
transform 1 0 3388 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_4294
timestamp 1745462530
transform 1 0 3388 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_4295
timestamp 1745462530
transform 1 0 3380 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_4296
timestamp 1745462530
transform 1 0 3348 0 1 1275
box -3 -3 3 3
use M3_M2  M3_M2_4297
timestamp 1745462530
transform 1 0 3332 0 1 2565
box -3 -3 3 3
use M3_M2  M3_M2_4298
timestamp 1745462530
transform 1 0 3332 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_4299
timestamp 1745462530
transform 1 0 3300 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_4300
timestamp 1745462530
transform 1 0 3212 0 1 2685
box -3 -3 3 3
use M3_M2  M3_M2_4301
timestamp 1745462530
transform 1 0 3212 0 1 2555
box -3 -3 3 3
use M3_M2  M3_M2_4302
timestamp 1745462530
transform 1 0 3204 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_4303
timestamp 1745462530
transform 1 0 3204 0 1 375
box -3 -3 3 3
use M3_M2  M3_M2_4304
timestamp 1745462530
transform 1 0 3116 0 1 2685
box -3 -3 3 3
use M3_M2  M3_M2_4305
timestamp 1745462530
transform 1 0 3108 0 1 2855
box -3 -3 3 3
use M3_M2  M3_M2_4306
timestamp 1745462530
transform 1 0 2924 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_4307
timestamp 1745462530
transform 1 0 2924 0 1 375
box -3 -3 3 3
use M3_M2  M3_M2_4308
timestamp 1745462530
transform 1 0 2868 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_4309
timestamp 1745462530
transform 1 0 2868 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_4310
timestamp 1745462530
transform 1 0 2460 0 1 2855
box -3 -3 3 3
use M3_M2  M3_M2_4311
timestamp 1745462530
transform 1 0 2308 0 1 475
box -3 -3 3 3
use M3_M2  M3_M2_4312
timestamp 1745462530
transform 1 0 2308 0 1 415
box -3 -3 3 3
use M3_M2  M3_M2_4313
timestamp 1745462530
transform 1 0 2220 0 1 475
box -3 -3 3 3
use M3_M2  M3_M2_4314
timestamp 1745462530
transform 1 0 1660 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_4315
timestamp 1745462530
transform 1 0 1644 0 1 2855
box -3 -3 3 3
use M3_M2  M3_M2_4316
timestamp 1745462530
transform 1 0 1644 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_4317
timestamp 1745462530
transform 1 0 1372 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_4318
timestamp 1745462530
transform 1 0 1332 0 1 2855
box -3 -3 3 3
use M3_M2  M3_M2_4319
timestamp 1745462530
transform 1 0 1292 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_4320
timestamp 1745462530
transform 1 0 1292 0 1 475
box -3 -3 3 3
use M3_M2  M3_M2_4321
timestamp 1745462530
transform 1 0 716 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_4322
timestamp 1745462530
transform 1 0 716 0 1 475
box -3 -3 3 3
use M3_M2  M3_M2_4323
timestamp 1745462530
transform 1 0 580 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_4324
timestamp 1745462530
transform 1 0 572 0 1 2855
box -3 -3 3 3
use M3_M2  M3_M2_4325
timestamp 1745462530
transform 1 0 508 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_4326
timestamp 1745462530
transform 1 0 3740 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_4327
timestamp 1745462530
transform 1 0 3732 0 1 2525
box -3 -3 3 3
use M3_M2  M3_M2_4328
timestamp 1745462530
transform 1 0 3724 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_4329
timestamp 1745462530
transform 1 0 3724 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_4330
timestamp 1745462530
transform 1 0 3708 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_4331
timestamp 1745462530
transform 1 0 3708 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_4332
timestamp 1745462530
transform 1 0 3628 0 1 2525
box -3 -3 3 3
use M3_M2  M3_M2_4333
timestamp 1745462530
transform 1 0 3620 0 1 2465
box -3 -3 3 3
use M3_M2  M3_M2_4334
timestamp 1745462530
transform 1 0 3620 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_4335
timestamp 1745462530
transform 1 0 2540 0 1 2465
box -3 -3 3 3
use M3_M2  M3_M2_4336
timestamp 1745462530
transform 1 0 2508 0 1 725
box -3 -3 3 3
use M3_M2  M3_M2_4337
timestamp 1745462530
transform 1 0 2492 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_4338
timestamp 1745462530
transform 1 0 2468 0 1 2495
box -3 -3 3 3
use M3_M2  M3_M2_4339
timestamp 1745462530
transform 1 0 2468 0 1 2465
box -3 -3 3 3
use M3_M2  M3_M2_4340
timestamp 1745462530
transform 1 0 2036 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_4341
timestamp 1745462530
transform 1 0 1852 0 1 2495
box -3 -3 3 3
use M3_M2  M3_M2_4342
timestamp 1745462530
transform 1 0 1068 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_4343
timestamp 1745462530
transform 1 0 876 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_4344
timestamp 1745462530
transform 1 0 876 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_4345
timestamp 1745462530
transform 1 0 812 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_4346
timestamp 1745462530
transform 1 0 788 0 1 2495
box -3 -3 3 3
use M3_M2  M3_M2_4347
timestamp 1745462530
transform 1 0 772 0 1 2495
box -3 -3 3 3
use M3_M2  M3_M2_4348
timestamp 1745462530
transform 1 0 3452 0 1 2245
box -3 -3 3 3
use M3_M2  M3_M2_4349
timestamp 1745462530
transform 1 0 3436 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_4350
timestamp 1745462530
transform 1 0 3420 0 1 2245
box -3 -3 3 3
use M3_M2  M3_M2_4351
timestamp 1745462530
transform 1 0 3412 0 1 2615
box -3 -3 3 3
use M3_M2  M3_M2_4352
timestamp 1745462530
transform 1 0 3412 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_4353
timestamp 1745462530
transform 1 0 3396 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_4354
timestamp 1745462530
transform 1 0 3380 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_4355
timestamp 1745462530
transform 1 0 2788 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_4356
timestamp 1745462530
transform 1 0 2508 0 1 2535
box -3 -3 3 3
use M3_M2  M3_M2_4357
timestamp 1745462530
transform 1 0 2500 0 1 2725
box -3 -3 3 3
use M3_M2  M3_M2_4358
timestamp 1745462530
transform 1 0 2500 0 1 2615
box -3 -3 3 3
use M3_M2  M3_M2_4359
timestamp 1745462530
transform 1 0 2460 0 1 2535
box -3 -3 3 3
use M3_M2  M3_M2_4360
timestamp 1745462530
transform 1 0 2452 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_4361
timestamp 1745462530
transform 1 0 2388 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_4362
timestamp 1745462530
transform 1 0 2388 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_4363
timestamp 1745462530
transform 1 0 1484 0 1 2735
box -3 -3 3 3
use M3_M2  M3_M2_4364
timestamp 1745462530
transform 1 0 1484 0 1 2705
box -3 -3 3 3
use M3_M2  M3_M2_4365
timestamp 1745462530
transform 1 0 1244 0 1 2705
box -3 -3 3 3
use M3_M2  M3_M2_4366
timestamp 1745462530
transform 1 0 1244 0 1 2645
box -3 -3 3 3
use M3_M2  M3_M2_4367
timestamp 1745462530
transform 1 0 1180 0 1 2645
box -3 -3 3 3
use M3_M2  M3_M2_4368
timestamp 1745462530
transform 1 0 1124 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_4369
timestamp 1745462530
transform 1 0 1124 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_4370
timestamp 1745462530
transform 1 0 1084 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_4371
timestamp 1745462530
transform 1 0 1076 0 1 2645
box -3 -3 3 3
use M3_M2  M3_M2_4372
timestamp 1745462530
transform 1 0 1076 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_4373
timestamp 1745462530
transform 1 0 1012 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_4374
timestamp 1745462530
transform 1 0 1012 0 1 2385
box -3 -3 3 3
use M3_M2  M3_M2_4375
timestamp 1745462530
transform 1 0 932 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_4376
timestamp 1745462530
transform 1 0 932 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_4377
timestamp 1745462530
transform 1 0 860 0 1 2385
box -3 -3 3 3
use M3_M2  M3_M2_4378
timestamp 1745462530
transform 1 0 844 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_4379
timestamp 1745462530
transform 1 0 796 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_4380
timestamp 1745462530
transform 1 0 4332 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_4381
timestamp 1745462530
transform 1 0 4332 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_4382
timestamp 1745462530
transform 1 0 4332 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_4383
timestamp 1745462530
transform 1 0 4324 0 1 2055
box -3 -3 3 3
use M3_M2  M3_M2_4384
timestamp 1745462530
transform 1 0 4092 0 1 2405
box -3 -3 3 3
use M3_M2  M3_M2_4385
timestamp 1745462530
transform 1 0 4012 0 1 2405
box -3 -3 3 3
use M3_M2  M3_M2_4386
timestamp 1745462530
transform 1 0 4004 0 1 2045
box -3 -3 3 3
use M3_M2  M3_M2_4387
timestamp 1745462530
transform 1 0 3964 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_4388
timestamp 1745462530
transform 1 0 3124 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_4389
timestamp 1745462530
transform 1 0 2428 0 1 2385
box -3 -3 3 3
use M3_M2  M3_M2_4390
timestamp 1745462530
transform 1 0 2236 0 1 2385
box -3 -3 3 3
use M3_M2  M3_M2_4391
timestamp 1745462530
transform 1 0 2236 0 1 2335
box -3 -3 3 3
use M3_M2  M3_M2_4392
timestamp 1745462530
transform 1 0 2036 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_4393
timestamp 1745462530
transform 1 0 1996 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_4394
timestamp 1745462530
transform 1 0 1996 0 1 2335
box -3 -3 3 3
use M3_M2  M3_M2_4395
timestamp 1745462530
transform 1 0 1788 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_4396
timestamp 1745462530
transform 1 0 1788 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_4397
timestamp 1745462530
transform 1 0 1612 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_4398
timestamp 1745462530
transform 1 0 636 0 1 2325
box -3 -3 3 3
use M3_M2  M3_M2_4399
timestamp 1745462530
transform 1 0 636 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_4400
timestamp 1745462530
transform 1 0 636 0 1 1205
box -3 -3 3 3
use M3_M2  M3_M2_4401
timestamp 1745462530
transform 1 0 636 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_4402
timestamp 1745462530
transform 1 0 604 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_4403
timestamp 1745462530
transform 1 0 604 0 1 1205
box -3 -3 3 3
use M3_M2  M3_M2_4404
timestamp 1745462530
transform 1 0 556 0 1 2325
box -3 -3 3 3
use M3_M2  M3_M2_4405
timestamp 1745462530
transform 1 0 3268 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_4406
timestamp 1745462530
transform 1 0 3260 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_4407
timestamp 1745462530
transform 1 0 3220 0 1 2495
box -3 -3 3 3
use M3_M2  M3_M2_4408
timestamp 1745462530
transform 1 0 3220 0 1 1495
box -3 -3 3 3
use M3_M2  M3_M2_4409
timestamp 1745462530
transform 1 0 3172 0 1 1495
box -3 -3 3 3
use M3_M2  M3_M2_4410
timestamp 1745462530
transform 1 0 3164 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_4411
timestamp 1745462530
transform 1 0 3028 0 1 665
box -3 -3 3 3
use M3_M2  M3_M2_4412
timestamp 1745462530
transform 1 0 3020 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_4413
timestamp 1745462530
transform 1 0 2500 0 1 2575
box -3 -3 3 3
use M3_M2  M3_M2_4414
timestamp 1745462530
transform 1 0 2500 0 1 2495
box -3 -3 3 3
use M3_M2  M3_M2_4415
timestamp 1745462530
transform 1 0 2252 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_4416
timestamp 1745462530
transform 1 0 2252 0 1 665
box -3 -3 3 3
use M3_M2  M3_M2_4417
timestamp 1745462530
transform 1 0 1604 0 1 2575
box -3 -3 3 3
use M3_M2  M3_M2_4418
timestamp 1745462530
transform 1 0 1516 0 1 725
box -3 -3 3 3
use M3_M2  M3_M2_4419
timestamp 1745462530
transform 1 0 1396 0 1 2575
box -3 -3 3 3
use M3_M2  M3_M2_4420
timestamp 1745462530
transform 1 0 1372 0 1 2635
box -3 -3 3 3
use M3_M2  M3_M2_4421
timestamp 1745462530
transform 1 0 1332 0 1 2635
box -3 -3 3 3
use M3_M2  M3_M2_4422
timestamp 1745462530
transform 1 0 1100 0 1 2635
box -3 -3 3 3
use M3_M2  M3_M2_4423
timestamp 1745462530
transform 1 0 1092 0 1 2475
box -3 -3 3 3
use M3_M2  M3_M2_4424
timestamp 1745462530
transform 1 0 892 0 1 2485
box -3 -3 3 3
use M3_M2  M3_M2_4425
timestamp 1745462530
transform 1 0 892 0 1 2465
box -3 -3 3 3
use M3_M2  M3_M2_4426
timestamp 1745462530
transform 1 0 620 0 1 2485
box -3 -3 3 3
use M3_M2  M3_M2_4427
timestamp 1745462530
transform 1 0 604 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_4428
timestamp 1745462530
transform 1 0 580 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_4429
timestamp 1745462530
transform 1 0 3692 0 1 2475
box -3 -3 3 3
use M3_M2  M3_M2_4430
timestamp 1745462530
transform 1 0 3668 0 1 975
box -3 -3 3 3
use M3_M2  M3_M2_4431
timestamp 1745462530
transform 1 0 3604 0 1 975
box -3 -3 3 3
use M3_M2  M3_M2_4432
timestamp 1745462530
transform 1 0 3588 0 1 2475
box -3 -3 3 3
use M3_M2  M3_M2_4433
timestamp 1745462530
transform 1 0 3588 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_4434
timestamp 1745462530
transform 1 0 3588 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_4435
timestamp 1745462530
transform 1 0 3588 0 1 975
box -3 -3 3 3
use M3_M2  M3_M2_4436
timestamp 1745462530
transform 1 0 3508 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_4437
timestamp 1745462530
transform 1 0 3300 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_4438
timestamp 1745462530
transform 1 0 3300 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_4439
timestamp 1745462530
transform 1 0 3276 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_4440
timestamp 1745462530
transform 1 0 3276 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_4441
timestamp 1745462530
transform 1 0 3220 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_4442
timestamp 1745462530
transform 1 0 2684 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_4443
timestamp 1745462530
transform 1 0 2684 0 1 1005
box -3 -3 3 3
use M3_M2  M3_M2_4444
timestamp 1745462530
transform 1 0 2532 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_4445
timestamp 1745462530
transform 1 0 2524 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_4446
timestamp 1745462530
transform 1 0 2524 0 1 1005
box -3 -3 3 3
use M3_M2  M3_M2_4447
timestamp 1745462530
transform 1 0 2148 0 1 1055
box -3 -3 3 3
use M3_M2  M3_M2_4448
timestamp 1745462530
transform 1 0 2148 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_4449
timestamp 1745462530
transform 1 0 1972 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_4450
timestamp 1745462530
transform 1 0 1940 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_4451
timestamp 1745462530
transform 1 0 1940 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_4452
timestamp 1745462530
transform 1 0 1220 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_4453
timestamp 1745462530
transform 1 0 1204 0 1 1055
box -3 -3 3 3
use M3_M2  M3_M2_4454
timestamp 1745462530
transform 1 0 1036 0 1 1055
box -3 -3 3 3
use M3_M2  M3_M2_4455
timestamp 1745462530
transform 1 0 772 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_4456
timestamp 1745462530
transform 1 0 772 0 1 2325
box -3 -3 3 3
use M3_M2  M3_M2_4457
timestamp 1745462530
transform 1 0 748 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_4458
timestamp 1745462530
transform 1 0 740 0 1 2315
box -3 -3 3 3
use M3_M2  M3_M2_4459
timestamp 1745462530
transform 1 0 732 0 1 2065
box -3 -3 3 3
use M3_M2  M3_M2_4460
timestamp 1745462530
transform 1 0 732 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_4461
timestamp 1745462530
transform 1 0 732 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_4462
timestamp 1745462530
transform 1 0 716 0 1 2065
box -3 -3 3 3
use M3_M2  M3_M2_4463
timestamp 1745462530
transform 1 0 3308 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_4464
timestamp 1745462530
transform 1 0 3292 0 1 2575
box -3 -3 3 3
use M3_M2  M3_M2_4465
timestamp 1745462530
transform 1 0 3252 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_4466
timestamp 1745462530
transform 1 0 3252 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_4467
timestamp 1745462530
transform 1 0 3212 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_4468
timestamp 1745462530
transform 1 0 3100 0 1 2575
box -3 -3 3 3
use M3_M2  M3_M2_4469
timestamp 1745462530
transform 1 0 3100 0 1 2375
box -3 -3 3 3
use M3_M2  M3_M2_4470
timestamp 1745462530
transform 1 0 3060 0 1 2375
box -3 -3 3 3
use M3_M2  M3_M2_4471
timestamp 1745462530
transform 1 0 3060 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_4472
timestamp 1745462530
transform 1 0 2764 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_4473
timestamp 1745462530
transform 1 0 2516 0 1 2655
box -3 -3 3 3
use M3_M2  M3_M2_4474
timestamp 1745462530
transform 1 0 2516 0 1 2575
box -3 -3 3 3
use M3_M2  M3_M2_4475
timestamp 1745462530
transform 1 0 2396 0 1 1205
box -3 -3 3 3
use M3_M2  M3_M2_4476
timestamp 1745462530
transform 1 0 2396 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_4477
timestamp 1745462530
transform 1 0 1492 0 1 2695
box -3 -3 3 3
use M3_M2  M3_M2_4478
timestamp 1745462530
transform 1 0 1492 0 1 2655
box -3 -3 3 3
use M3_M2  M3_M2_4479
timestamp 1745462530
transform 1 0 1164 0 1 2695
box -3 -3 3 3
use M3_M2  M3_M2_4480
timestamp 1745462530
transform 1 0 1092 0 1 1205
box -3 -3 3 3
use M3_M2  M3_M2_4481
timestamp 1745462530
transform 1 0 1052 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_4482
timestamp 1745462530
transform 1 0 1052 0 1 1205
box -3 -3 3 3
use M3_M2  M3_M2_4483
timestamp 1745462530
transform 1 0 964 0 1 1285
box -3 -3 3 3
use M3_M2  M3_M2_4484
timestamp 1745462530
transform 1 0 964 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_4485
timestamp 1745462530
transform 1 0 892 0 1 1875
box -3 -3 3 3
use M3_M2  M3_M2_4486
timestamp 1745462530
transform 1 0 892 0 1 1285
box -3 -3 3 3
use M3_M2  M3_M2_4487
timestamp 1745462530
transform 1 0 868 0 1 1875
box -3 -3 3 3
use M3_M2  M3_M2_4488
timestamp 1745462530
transform 1 0 284 0 1 2695
box -3 -3 3 3
use M3_M2  M3_M2_4489
timestamp 1745462530
transform 1 0 284 0 1 1875
box -3 -3 3 3
use M3_M2  M3_M2_4490
timestamp 1745462530
transform 1 0 4324 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_4491
timestamp 1745462530
transform 1 0 4324 0 1 1045
box -3 -3 3 3
use M3_M2  M3_M2_4492
timestamp 1745462530
transform 1 0 4284 0 1 2065
box -3 -3 3 3
use M3_M2  M3_M2_4493
timestamp 1745462530
transform 1 0 4284 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_4494
timestamp 1745462530
transform 1 0 4220 0 1 2065
box -3 -3 3 3
use M3_M2  M3_M2_4495
timestamp 1745462530
transform 1 0 4212 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_4496
timestamp 1745462530
transform 1 0 4148 0 1 2095
box -3 -3 3 3
use M3_M2  M3_M2_4497
timestamp 1745462530
transform 1 0 4148 0 1 2065
box -3 -3 3 3
use M3_M2  M3_M2_4498
timestamp 1745462530
transform 1 0 4028 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_4499
timestamp 1745462530
transform 1 0 4004 0 1 1055
box -3 -3 3 3
use M3_M2  M3_M2_4500
timestamp 1745462530
transform 1 0 3956 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_4501
timestamp 1745462530
transform 1 0 3948 0 1 1055
box -3 -3 3 3
use M3_M2  M3_M2_4502
timestamp 1745462530
transform 1 0 3932 0 1 2095
box -3 -3 3 3
use M3_M2  M3_M2_4503
timestamp 1745462530
transform 1 0 3156 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_4504
timestamp 1745462530
transform 1 0 2540 0 1 2265
box -3 -3 3 3
use M3_M2  M3_M2_4505
timestamp 1745462530
transform 1 0 2212 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_4506
timestamp 1745462530
transform 1 0 2212 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_4507
timestamp 1745462530
transform 1 0 2180 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_4508
timestamp 1745462530
transform 1 0 2180 0 1 1675
box -3 -3 3 3
use M3_M2  M3_M2_4509
timestamp 1745462530
transform 1 0 2156 0 1 1675
box -3 -3 3 3
use M3_M2  M3_M2_4510
timestamp 1745462530
transform 1 0 2156 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_4511
timestamp 1745462530
transform 1 0 2140 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_4512
timestamp 1745462530
transform 1 0 2124 0 1 2245
box -3 -3 3 3
use M3_M2  M3_M2_4513
timestamp 1745462530
transform 1 0 2044 0 1 2245
box -3 -3 3 3
use M3_M2  M3_M2_4514
timestamp 1745462530
transform 1 0 1844 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_4515
timestamp 1745462530
transform 1 0 1740 0 1 1215
box -3 -3 3 3
use M3_M2  M3_M2_4516
timestamp 1745462530
transform 1 0 1740 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_4517
timestamp 1745462530
transform 1 0 596 0 1 2085
box -3 -3 3 3
use M3_M2  M3_M2_4518
timestamp 1745462530
transform 1 0 572 0 1 1265
box -3 -3 3 3
use M3_M2  M3_M2_4519
timestamp 1745462530
transform 1 0 572 0 1 1215
box -3 -3 3 3
use M3_M2  M3_M2_4520
timestamp 1745462530
transform 1 0 532 0 1 1265
box -3 -3 3 3
use M3_M2  M3_M2_4521
timestamp 1745462530
transform 1 0 516 0 1 2085
box -3 -3 3 3
use M3_M2  M3_M2_4522
timestamp 1745462530
transform 1 0 3108 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_4523
timestamp 1745462530
transform 1 0 3092 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_4524
timestamp 1745462530
transform 1 0 3092 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_4525
timestamp 1745462530
transform 1 0 3060 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_4526
timestamp 1745462530
transform 1 0 3060 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_4527
timestamp 1745462530
transform 1 0 3036 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_4528
timestamp 1745462530
transform 1 0 3036 0 1 2375
box -3 -3 3 3
use M3_M2  M3_M2_4529
timestamp 1745462530
transform 1 0 3028 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_4530
timestamp 1745462530
transform 1 0 2964 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_4531
timestamp 1745462530
transform 1 0 2964 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_4532
timestamp 1745462530
transform 1 0 2892 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_4533
timestamp 1745462530
transform 1 0 2892 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_4534
timestamp 1745462530
transform 1 0 2700 0 1 2055
box -3 -3 3 3
use M3_M2  M3_M2_4535
timestamp 1745462530
transform 1 0 2700 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_4536
timestamp 1745462530
transform 1 0 2636 0 1 2385
box -3 -3 3 3
use M3_M2  M3_M2_4537
timestamp 1745462530
transform 1 0 2620 0 1 2065
box -3 -3 3 3
use M3_M2  M3_M2_4538
timestamp 1745462530
transform 1 0 2564 0 1 2385
box -3 -3 3 3
use M3_M2  M3_M2_4539
timestamp 1745462530
transform 1 0 2220 0 1 1065
box -3 -3 3 3
use M3_M2  M3_M2_4540
timestamp 1745462530
transform 1 0 2220 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_4541
timestamp 1745462530
transform 1 0 1652 0 1 2585
box -3 -3 3 3
use M3_M2  M3_M2_4542
timestamp 1745462530
transform 1 0 1548 0 1 1065
box -3 -3 3 3
use M3_M2  M3_M2_4543
timestamp 1745462530
transform 1 0 1548 0 1 1035
box -3 -3 3 3
use M3_M2  M3_M2_4544
timestamp 1745462530
transform 1 0 1364 0 1 2585
box -3 -3 3 3
use M3_M2  M3_M2_4545
timestamp 1745462530
transform 1 0 652 0 1 2285
box -3 -3 3 3
use M3_M2  M3_M2_4546
timestamp 1745462530
transform 1 0 596 0 1 1035
box -3 -3 3 3
use M3_M2  M3_M2_4547
timestamp 1745462530
transform 1 0 588 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_4548
timestamp 1745462530
transform 1 0 468 0 1 2285
box -3 -3 3 3
use M3_M2  M3_M2_4549
timestamp 1745462530
transform 1 0 452 0 1 2585
box -3 -3 3 3
use M3_M2  M3_M2_4550
timestamp 1745462530
transform 1 0 156 0 1 2285
box -3 -3 3 3
use M3_M2  M3_M2_4551
timestamp 1745462530
transform 1 0 156 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_4552
timestamp 1745462530
transform 1 0 3652 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_4553
timestamp 1745462530
transform 1 0 3644 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_4554
timestamp 1745462530
transform 1 0 3636 0 1 2535
box -3 -3 3 3
use M3_M2  M3_M2_4555
timestamp 1745462530
transform 1 0 3588 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_4556
timestamp 1745462530
transform 1 0 3508 0 1 2535
box -3 -3 3 3
use M3_M2  M3_M2_4557
timestamp 1745462530
transform 1 0 3300 0 1 1275
box -3 -3 3 3
use M3_M2  M3_M2_4558
timestamp 1745462530
transform 1 0 3300 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_4559
timestamp 1745462530
transform 1 0 3236 0 1 1335
box -3 -3 3 3
use M3_M2  M3_M2_4560
timestamp 1745462530
transform 1 0 3236 0 1 1275
box -3 -3 3 3
use M3_M2  M3_M2_4561
timestamp 1745462530
transform 1 0 3204 0 1 1335
box -3 -3 3 3
use M3_M2  M3_M2_4562
timestamp 1745462530
transform 1 0 2548 0 1 2535
box -3 -3 3 3
use M3_M2  M3_M2_4563
timestamp 1745462530
transform 1 0 2540 0 1 1275
box -3 -3 3 3
use M3_M2  M3_M2_4564
timestamp 1745462530
transform 1 0 2540 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_4565
timestamp 1745462530
transform 1 0 2516 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_4566
timestamp 1745462530
transform 1 0 2340 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_4567
timestamp 1745462530
transform 1 0 2340 0 1 1015
box -3 -3 3 3
use M3_M2  M3_M2_4568
timestamp 1745462530
transform 1 0 2132 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_4569
timestamp 1745462530
transform 1 0 1940 0 1 2525
box -3 -3 3 3
use M3_M2  M3_M2_4570
timestamp 1745462530
transform 1 0 1932 0 1 2455
box -3 -3 3 3
use M3_M2  M3_M2_4571
timestamp 1745462530
transform 1 0 1012 0 1 1005
box -3 -3 3 3
use M3_M2  M3_M2_4572
timestamp 1745462530
transform 1 0 1012 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_4573
timestamp 1745462530
transform 1 0 876 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_4574
timestamp 1745462530
transform 1 0 876 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_4575
timestamp 1745462530
transform 1 0 756 0 1 2455
box -3 -3 3 3
use M3_M2  M3_M2_4576
timestamp 1745462530
transform 1 0 724 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_4577
timestamp 1745462530
transform 1 0 3292 0 1 1065
box -3 -3 3 3
use M3_M2  M3_M2_4578
timestamp 1745462530
transform 1 0 3276 0 1 2565
box -3 -3 3 3
use M3_M2  M3_M2_4579
timestamp 1745462530
transform 1 0 3188 0 1 2175
box -3 -3 3 3
use M3_M2  M3_M2_4580
timestamp 1745462530
transform 1 0 3156 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_4581
timestamp 1745462530
transform 1 0 3156 0 1 1065
box -3 -3 3 3
use M3_M2  M3_M2_4582
timestamp 1745462530
transform 1 0 3140 0 1 2175
box -3 -3 3 3
use M3_M2  M3_M2_4583
timestamp 1745462530
transform 1 0 3140 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_4584
timestamp 1745462530
transform 1 0 3108 0 1 2555
box -3 -3 3 3
use M3_M2  M3_M2_4585
timestamp 1745462530
transform 1 0 3036 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_4586
timestamp 1745462530
transform 1 0 3036 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_4587
timestamp 1745462530
transform 1 0 2748 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_4588
timestamp 1745462530
transform 1 0 2588 0 1 2555
box -3 -3 3 3
use M3_M2  M3_M2_4589
timestamp 1745462530
transform 1 0 2372 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_4590
timestamp 1745462530
transform 1 0 1468 0 1 2655
box -3 -3 3 3
use M3_M2  M3_M2_4591
timestamp 1745462530
transform 1 0 1468 0 1 2555
box -3 -3 3 3
use M3_M2  M3_M2_4592
timestamp 1745462530
transform 1 0 1156 0 1 2655
box -3 -3 3 3
use M3_M2  M3_M2_4593
timestamp 1745462530
transform 1 0 1044 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_4594
timestamp 1745462530
transform 1 0 932 0 1 1135
box -3 -3 3 3
use M3_M2  M3_M2_4595
timestamp 1745462530
transform 1 0 884 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_4596
timestamp 1745462530
transform 1 0 860 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_4597
timestamp 1745462530
transform 1 0 3980 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_4598
timestamp 1745462530
transform 1 0 3972 0 1 2425
box -3 -3 3 3
use M3_M2  M3_M2_4599
timestamp 1745462530
transform 1 0 3972 0 1 2385
box -3 -3 3 3
use M3_M2  M3_M2_4600
timestamp 1745462530
transform 1 0 3940 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_4601
timestamp 1745462530
transform 1 0 3908 0 1 2385
box -3 -3 3 3
use M3_M2  M3_M2_4602
timestamp 1745462530
transform 1 0 3900 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_4603
timestamp 1745462530
transform 1 0 3140 0 1 1135
box -3 -3 3 3
use M3_M2  M3_M2_4604
timestamp 1745462530
transform 1 0 2612 0 1 2415
box -3 -3 3 3
use M3_M2  M3_M2_4605
timestamp 1745462530
transform 1 0 2044 0 1 2415
box -3 -3 3 3
use M3_M2  M3_M2_4606
timestamp 1745462530
transform 1 0 1828 0 1 1135
box -3 -3 3 3
use M3_M2  M3_M2_4607
timestamp 1745462530
transform 1 0 1732 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_4608
timestamp 1745462530
transform 1 0 1724 0 1 1135
box -3 -3 3 3
use M3_M2  M3_M2_4609
timestamp 1745462530
transform 1 0 588 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_4610
timestamp 1745462530
transform 1 0 540 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_4611
timestamp 1745462530
transform 1 0 516 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_4612
timestamp 1745462530
transform 1 0 476 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_4613
timestamp 1745462530
transform 1 0 3076 0 1 1085
box -3 -3 3 3
use M3_M2  M3_M2_4614
timestamp 1745462530
transform 1 0 3060 0 1 2535
box -3 -3 3 3
use M3_M2  M3_M2_4615
timestamp 1745462530
transform 1 0 3060 0 1 1465
box -3 -3 3 3
use M3_M2  M3_M2_4616
timestamp 1745462530
transform 1 0 3012 0 1 1465
box -3 -3 3 3
use M3_M2  M3_M2_4617
timestamp 1745462530
transform 1 0 2956 0 1 1465
box -3 -3 3 3
use M3_M2  M3_M2_4618
timestamp 1745462530
transform 1 0 2932 0 1 1085
box -3 -3 3 3
use M3_M2  M3_M2_4619
timestamp 1745462530
transform 1 0 2636 0 1 2605
box -3 -3 3 3
use M3_M2  M3_M2_4620
timestamp 1745462530
transform 1 0 2612 0 1 2605
box -3 -3 3 3
use M3_M2  M3_M2_4621
timestamp 1745462530
transform 1 0 2612 0 1 2535
box -3 -3 3 3
use M3_M2  M3_M2_4622
timestamp 1745462530
transform 1 0 2204 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_4623
timestamp 1745462530
transform 1 0 2204 0 1 1085
box -3 -3 3 3
use M3_M2  M3_M2_4624
timestamp 1745462530
transform 1 0 1692 0 1 2625
box -3 -3 3 3
use M3_M2  M3_M2_4625
timestamp 1745462530
transform 1 0 1692 0 1 2605
box -3 -3 3 3
use M3_M2  M3_M2_4626
timestamp 1745462530
transform 1 0 1636 0 1 2625
box -3 -3 3 3
use M3_M2  M3_M2_4627
timestamp 1745462530
transform 1 0 1524 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_4628
timestamp 1745462530
transform 1 0 1524 0 1 1075
box -3 -3 3 3
use M3_M2  M3_M2_4629
timestamp 1745462530
transform 1 0 1348 0 1 2625
box -3 -3 3 3
use M3_M2  M3_M2_4630
timestamp 1745462530
transform 1 0 628 0 1 2055
box -3 -3 3 3
use M3_M2  M3_M2_4631
timestamp 1745462530
transform 1 0 612 0 1 2315
box -3 -3 3 3
use M3_M2  M3_M2_4632
timestamp 1745462530
transform 1 0 612 0 1 2055
box -3 -3 3 3
use M3_M2  M3_M2_4633
timestamp 1745462530
transform 1 0 612 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_4634
timestamp 1745462530
transform 1 0 572 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_4635
timestamp 1745462530
transform 1 0 572 0 1 1075
box -3 -3 3 3
use M3_M2  M3_M2_4636
timestamp 1745462530
transform 1 0 436 0 1 2625
box -3 -3 3 3
use M3_M2  M3_M2_4637
timestamp 1745462530
transform 1 0 436 0 1 2585
box -3 -3 3 3
use M3_M2  M3_M2_4638
timestamp 1745462530
transform 1 0 340 0 1 2315
box -3 -3 3 3
use M3_M2  M3_M2_4639
timestamp 1745462530
transform 1 0 332 0 1 2585
box -3 -3 3 3
use M3_M2  M3_M2_4640
timestamp 1745462530
transform 1 0 3124 0 1 3495
box -3 -3 3 3
use M3_M2  M3_M2_4641
timestamp 1745462530
transform 1 0 2804 0 1 3505
box -3 -3 3 3
use M3_M2  M3_M2_4642
timestamp 1745462530
transform 1 0 2804 0 1 3435
box -3 -3 3 3
use M3_M2  M3_M2_4643
timestamp 1745462530
transform 1 0 2332 0 1 3435
box -3 -3 3 3
use M3_M2  M3_M2_4644
timestamp 1745462530
transform 1 0 2332 0 1 3245
box -3 -3 3 3
use M3_M2  M3_M2_4645
timestamp 1745462530
transform 1 0 2212 0 1 3245
box -3 -3 3 3
use M3_M2  M3_M2_4646
timestamp 1745462530
transform 1 0 2164 0 1 3245
box -3 -3 3 3
use M3_M2  M3_M2_4647
timestamp 1745462530
transform 1 0 3852 0 1 3245
box -3 -3 3 3
use M3_M2  M3_M2_4648
timestamp 1745462530
transform 1 0 3836 0 1 3245
box -3 -3 3 3
use M3_M2  M3_M2_4649
timestamp 1745462530
transform 1 0 3820 0 1 3245
box -3 -3 3 3
use M3_M2  M3_M2_4650
timestamp 1745462530
transform 1 0 3772 0 1 3245
box -3 -3 3 3
use M3_M2  M3_M2_4651
timestamp 1745462530
transform 1 0 3772 0 1 3215
box -3 -3 3 3
use M3_M2  M3_M2_4652
timestamp 1745462530
transform 1 0 3724 0 1 3215
box -3 -3 3 3
use M3_M2  M3_M2_4653
timestamp 1745462530
transform 1 0 3684 0 1 3215
box -3 -3 3 3
use M3_M2  M3_M2_4654
timestamp 1745462530
transform 1 0 3684 0 1 3165
box -3 -3 3 3
use M3_M2  M3_M2_4655
timestamp 1745462530
transform 1 0 2092 0 1 3165
box -3 -3 3 3
use M3_M2  M3_M2_4656
timestamp 1745462530
transform 1 0 2084 0 1 3265
box -3 -3 3 3
use M3_M2  M3_M2_4657
timestamp 1745462530
transform 1 0 2004 0 1 3265
box -3 -3 3 3
use M3_M2  M3_M2_4658
timestamp 1745462530
transform 1 0 1940 0 1 3255
box -3 -3 3 3
use M3_M2  M3_M2_4659
timestamp 1745462530
transform 1 0 1884 0 1 3255
box -3 -3 3 3
use M3_M2  M3_M2_4660
timestamp 1745462530
transform 1 0 1844 0 1 3255
box -3 -3 3 3
use M3_M2  M3_M2_4661
timestamp 1745462530
transform 1 0 3868 0 1 3455
box -3 -3 3 3
use M3_M2  M3_M2_4662
timestamp 1745462530
transform 1 0 3836 0 1 3455
box -3 -3 3 3
use M3_M2  M3_M2_4663
timestamp 1745462530
transform 1 0 3812 0 1 3455
box -3 -3 3 3
use M3_M2  M3_M2_4664
timestamp 1745462530
transform 1 0 3796 0 1 3395
box -3 -3 3 3
use M3_M2  M3_M2_4665
timestamp 1745462530
transform 1 0 3764 0 1 3455
box -3 -3 3 3
use M3_M2  M3_M2_4666
timestamp 1745462530
transform 1 0 3764 0 1 3395
box -3 -3 3 3
use M3_M2  M3_M2_4667
timestamp 1745462530
transform 1 0 3020 0 1 3455
box -3 -3 3 3
use M3_M2  M3_M2_4668
timestamp 1745462530
transform 1 0 2652 0 1 3385
box -3 -3 3 3
use M3_M2  M3_M2_4669
timestamp 1745462530
transform 1 0 2628 0 1 3455
box -3 -3 3 3
use M3_M2  M3_M2_4670
timestamp 1745462530
transform 1 0 2628 0 1 3385
box -3 -3 3 3
use M3_M2  M3_M2_4671
timestamp 1745462530
transform 1 0 2068 0 1 3245
box -3 -3 3 3
use M3_M2  M3_M2_4672
timestamp 1745462530
transform 1 0 1996 0 1 3385
box -3 -3 3 3
use M3_M2  M3_M2_4673
timestamp 1745462530
transform 1 0 1996 0 1 3245
box -3 -3 3 3
use M3_M2  M3_M2_4674
timestamp 1745462530
transform 1 0 1924 0 1 3385
box -3 -3 3 3
use M3_M2  M3_M2_4675
timestamp 1745462530
transform 1 0 3884 0 1 3525
box -3 -3 3 3
use M3_M2  M3_M2_4676
timestamp 1745462530
transform 1 0 3828 0 1 3635
box -3 -3 3 3
use M3_M2  M3_M2_4677
timestamp 1745462530
transform 1 0 3828 0 1 3535
box -3 -3 3 3
use M3_M2  M3_M2_4678
timestamp 1745462530
transform 1 0 3796 0 1 3635
box -3 -3 3 3
use M3_M2  M3_M2_4679
timestamp 1745462530
transform 1 0 3772 0 1 3525
box -3 -3 3 3
use M3_M2  M3_M2_4680
timestamp 1745462530
transform 1 0 3756 0 1 3725
box -3 -3 3 3
use M3_M2  M3_M2_4681
timestamp 1745462530
transform 1 0 3756 0 1 3635
box -3 -3 3 3
use M3_M2  M3_M2_4682
timestamp 1745462530
transform 1 0 3740 0 1 3765
box -3 -3 3 3
use M3_M2  M3_M2_4683
timestamp 1745462530
transform 1 0 3740 0 1 3725
box -3 -3 3 3
use M3_M2  M3_M2_4684
timestamp 1745462530
transform 1 0 3684 0 1 3725
box -3 -3 3 3
use M3_M2  M3_M2_4685
timestamp 1745462530
transform 1 0 2948 0 1 3765
box -3 -3 3 3
use M3_M2  M3_M2_4686
timestamp 1745462530
transform 1 0 2948 0 1 3635
box -3 -3 3 3
use M3_M2  M3_M2_4687
timestamp 1745462530
transform 1 0 2940 0 1 3715
box -3 -3 3 3
use M3_M2  M3_M2_4688
timestamp 1745462530
transform 1 0 2932 0 1 3635
box -3 -3 3 3
use M3_M2  M3_M2_4689
timestamp 1745462530
transform 1 0 2740 0 1 3705
box -3 -3 3 3
use M3_M2  M3_M2_4690
timestamp 1745462530
transform 1 0 2492 0 1 3715
box -3 -3 3 3
use M3_M2  M3_M2_4691
timestamp 1745462530
transform 1 0 2476 0 1 3655
box -3 -3 3 3
use M3_M2  M3_M2_4692
timestamp 1745462530
transform 1 0 2276 0 1 3655
box -3 -3 3 3
use M3_M2  M3_M2_4693
timestamp 1745462530
transform 1 0 2276 0 1 3575
box -3 -3 3 3
use M3_M2  M3_M2_4694
timestamp 1745462530
transform 1 0 2228 0 1 3575
box -3 -3 3 3
use M3_M2  M3_M2_4695
timestamp 1745462530
transform 1 0 3252 0 1 3705
box -3 -3 3 3
use M3_M2  M3_M2_4696
timestamp 1745462530
transform 1 0 3220 0 1 3705
box -3 -3 3 3
use M3_M2  M3_M2_4697
timestamp 1745462530
transform 1 0 3204 0 1 3705
box -3 -3 3 3
use M3_M2  M3_M2_4698
timestamp 1745462530
transform 1 0 3180 0 1 3705
box -3 -3 3 3
use M3_M2  M3_M2_4699
timestamp 1745462530
transform 1 0 3148 0 1 3705
box -3 -3 3 3
use M3_M2  M3_M2_4700
timestamp 1745462530
transform 1 0 3012 0 1 3705
box -3 -3 3 3
use M3_M2  M3_M2_4701
timestamp 1745462530
transform 1 0 2900 0 1 3705
box -3 -3 3 3
use M3_M2  M3_M2_4702
timestamp 1745462530
transform 1 0 2900 0 1 3665
box -3 -3 3 3
use M3_M2  M3_M2_4703
timestamp 1745462530
transform 1 0 2796 0 1 3665
box -3 -3 3 3
use M3_M2  M3_M2_4704
timestamp 1745462530
transform 1 0 2764 0 1 3695
box -3 -3 3 3
use M3_M2  M3_M2_4705
timestamp 1745462530
transform 1 0 2452 0 1 3705
box -3 -3 3 3
use M3_M2  M3_M2_4706
timestamp 1745462530
transform 1 0 2380 0 1 3705
box -3 -3 3 3
use M3_M2  M3_M2_4707
timestamp 1745462530
transform 1 0 2300 0 1 3705
box -3 -3 3 3
use M3_M2  M3_M2_4708
timestamp 1745462530
transform 1 0 2244 0 1 3705
box -3 -3 3 3
use M3_M2  M3_M2_4709
timestamp 1745462530
transform 1 0 3620 0 1 3655
box -3 -3 3 3
use M3_M2  M3_M2_4710
timestamp 1745462530
transform 1 0 3548 0 1 3655
box -3 -3 3 3
use M3_M2  M3_M2_4711
timestamp 1745462530
transform 1 0 3444 0 1 3655
box -3 -3 3 3
use M3_M2  M3_M2_4712
timestamp 1745462530
transform 1 0 3372 0 1 3655
box -3 -3 3 3
use M3_M2  M3_M2_4713
timestamp 1745462530
transform 1 0 3148 0 1 3655
box -3 -3 3 3
use M3_M2  M3_M2_4714
timestamp 1745462530
transform 1 0 3092 0 1 3655
box -3 -3 3 3
use M3_M2  M3_M2_4715
timestamp 1745462530
transform 1 0 2996 0 1 3655
box -3 -3 3 3
use M3_M2  M3_M2_4716
timestamp 1745462530
transform 1 0 2852 0 1 3655
box -3 -3 3 3
use M3_M2  M3_M2_4717
timestamp 1745462530
transform 1 0 2692 0 1 3655
box -3 -3 3 3
use M3_M2  M3_M2_4718
timestamp 1745462530
transform 1 0 2692 0 1 3625
box -3 -3 3 3
use M3_M2  M3_M2_4719
timestamp 1745462530
transform 1 0 2364 0 1 3615
box -3 -3 3 3
use M3_M2  M3_M2_4720
timestamp 1745462530
transform 1 0 2204 0 1 3615
box -3 -3 3 3
use M3_M2  M3_M2_4721
timestamp 1745462530
transform 1 0 2180 0 1 3615
box -3 -3 3 3
use M3_M2  M3_M2_4722
timestamp 1745462530
transform 1 0 2092 0 1 3135
box -3 -3 3 3
use M3_M2  M3_M2_4723
timestamp 1745462530
transform 1 0 2068 0 1 3135
box -3 -3 3 3
use M3_M2  M3_M2_4724
timestamp 1745462530
transform 1 0 2212 0 1 3625
box -3 -3 3 3
use M3_M2  M3_M2_4725
timestamp 1745462530
transform 1 0 2188 0 1 3625
box -3 -3 3 3
use M3_M2  M3_M2_4726
timestamp 1745462530
transform 1 0 2668 0 1 2355
box -3 -3 3 3
use M3_M2  M3_M2_4727
timestamp 1745462530
transform 1 0 2316 0 1 2355
box -3 -3 3 3
use M3_M2  M3_M2_4728
timestamp 1745462530
transform 1 0 2308 0 1 2175
box -3 -3 3 3
use M3_M2  M3_M2_4729
timestamp 1745462530
transform 1 0 2284 0 1 2175
box -3 -3 3 3
use M3_M2  M3_M2_4730
timestamp 1745462530
transform 1 0 2284 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_4731
timestamp 1745462530
transform 1 0 2260 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_4732
timestamp 1745462530
transform 1 0 2252 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_4733
timestamp 1745462530
transform 1 0 2164 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_4734
timestamp 1745462530
transform 1 0 1580 0 1 1835
box -3 -3 3 3
use M3_M2  M3_M2_4735
timestamp 1745462530
transform 1 0 1580 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_4736
timestamp 1745462530
transform 1 0 1508 0 1 1835
box -3 -3 3 3
use M3_M2  M3_M2_4737
timestamp 1745462530
transform 1 0 2988 0 1 2695
box -3 -3 3 3
use M3_M2  M3_M2_4738
timestamp 1745462530
transform 1 0 2956 0 1 2695
box -3 -3 3 3
use M3_M2  M3_M2_4739
timestamp 1745462530
transform 1 0 2684 0 1 2695
box -3 -3 3 3
use M3_M2  M3_M2_4740
timestamp 1745462530
transform 1 0 2684 0 1 2645
box -3 -3 3 3
use M3_M2  M3_M2_4741
timestamp 1745462530
transform 1 0 1300 0 1 2645
box -3 -3 3 3
use M3_M2  M3_M2_4742
timestamp 1745462530
transform 1 0 1292 0 1 2685
box -3 -3 3 3
use M3_M2  M3_M2_4743
timestamp 1745462530
transform 1 0 1220 0 1 2675
box -3 -3 3 3
use M3_M2  M3_M2_4744
timestamp 1745462530
transform 1 0 1212 0 1 2935
box -3 -3 3 3
use M3_M2  M3_M2_4745
timestamp 1745462530
transform 1 0 1188 0 1 2935
box -3 -3 3 3
use M3_M2  M3_M2_4746
timestamp 1745462530
transform 1 0 1180 0 1 3115
box -3 -3 3 3
use M3_M2  M3_M2_4747
timestamp 1745462530
transform 1 0 900 0 1 3115
box -3 -3 3 3
use M3_M2  M3_M2_4748
timestamp 1745462530
transform 1 0 1508 0 1 1935
box -3 -3 3 3
use M3_M2  M3_M2_4749
timestamp 1745462530
transform 1 0 1484 0 1 2385
box -3 -3 3 3
use M3_M2  M3_M2_4750
timestamp 1745462530
transform 1 0 1460 0 1 2385
box -3 -3 3 3
use M3_M2  M3_M2_4751
timestamp 1745462530
transform 1 0 724 0 1 1935
box -3 -3 3 3
use M3_M2  M3_M2_4752
timestamp 1745462530
transform 1 0 644 0 1 1935
box -3 -3 3 3
use M3_M2  M3_M2_4753
timestamp 1745462530
transform 1 0 532 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_4754
timestamp 1745462530
transform 1 0 492 0 1 1935
box -3 -3 3 3
use M3_M2  M3_M2_4755
timestamp 1745462530
transform 1 0 1612 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_4756
timestamp 1745462530
transform 1 0 1500 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_4757
timestamp 1745462530
transform 1 0 1476 0 1 1135
box -3 -3 3 3
use M3_M2  M3_M2_4758
timestamp 1745462530
transform 1 0 1460 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_4759
timestamp 1745462530
transform 1 0 1460 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_4760
timestamp 1745462530
transform 1 0 1092 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_4761
timestamp 1745462530
transform 1 0 1044 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_4762
timestamp 1745462530
transform 1 0 1028 0 1 1135
box -3 -3 3 3
use M3_M2  M3_M2_4763
timestamp 1745462530
transform 1 0 1028 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_4764
timestamp 1745462530
transform 1 0 988 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_4765
timestamp 1745462530
transform 1 0 980 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_4766
timestamp 1745462530
transform 1 0 980 0 1 1085
box -3 -3 3 3
use M3_M2  M3_M2_4767
timestamp 1745462530
transform 1 0 940 0 1 1085
box -3 -3 3 3
use M3_M2  M3_M2_4768
timestamp 1745462530
transform 1 0 932 0 1 975
box -3 -3 3 3
use M3_M2  M3_M2_4769
timestamp 1745462530
transform 1 0 3252 0 1 1015
box -3 -3 3 3
use M3_M2  M3_M2_4770
timestamp 1745462530
transform 1 0 3164 0 1 1015
box -3 -3 3 3
use M3_M2  M3_M2_4771
timestamp 1745462530
transform 1 0 2836 0 1 1015
box -3 -3 3 3
use M3_M2  M3_M2_4772
timestamp 1745462530
transform 1 0 2796 0 1 1015
box -3 -3 3 3
use M3_M2  M3_M2_4773
timestamp 1745462530
transform 1 0 2732 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_4774
timestamp 1745462530
transform 1 0 2708 0 1 1015
box -3 -3 3 3
use M3_M2  M3_M2_4775
timestamp 1745462530
transform 1 0 2404 0 1 2255
box -3 -3 3 3
use M3_M2  M3_M2_4776
timestamp 1745462530
transform 1 0 2356 0 1 2175
box -3 -3 3 3
use M3_M2  M3_M2_4777
timestamp 1745462530
transform 1 0 2340 0 1 2255
box -3 -3 3 3
use M3_M2  M3_M2_4778
timestamp 1745462530
transform 1 0 2340 0 1 2175
box -3 -3 3 3
use M3_M2  M3_M2_4779
timestamp 1745462530
transform 1 0 2340 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_4780
timestamp 1745462530
transform 1 0 2308 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_4781
timestamp 1745462530
transform 1 0 3452 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_4782
timestamp 1745462530
transform 1 0 3452 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_4783
timestamp 1745462530
transform 1 0 3420 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_4784
timestamp 1745462530
transform 1 0 3412 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_4785
timestamp 1745462530
transform 1 0 3412 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_4786
timestamp 1745462530
transform 1 0 3396 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_4787
timestamp 1745462530
transform 1 0 3388 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_4788
timestamp 1745462530
transform 1 0 2180 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_4789
timestamp 1745462530
transform 1 0 2180 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_4790
timestamp 1745462530
transform 1 0 2036 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_4791
timestamp 1745462530
transform 1 0 3148 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_4792
timestamp 1745462530
transform 1 0 3036 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_4793
timestamp 1745462530
transform 1 0 2996 0 1 2415
box -3 -3 3 3
use M3_M2  M3_M2_4794
timestamp 1745462530
transform 1 0 2996 0 1 2325
box -3 -3 3 3
use M3_M2  M3_M2_4795
timestamp 1745462530
transform 1 0 2980 0 1 2415
box -3 -3 3 3
use M3_M2  M3_M2_4796
timestamp 1745462530
transform 1 0 2956 0 1 2325
box -3 -3 3 3
use M3_M2  M3_M2_4797
timestamp 1745462530
transform 1 0 2932 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_4798
timestamp 1745462530
transform 1 0 3092 0 1 2705
box -3 -3 3 3
use M3_M2  M3_M2_4799
timestamp 1745462530
transform 1 0 3060 0 1 2725
box -3 -3 3 3
use M3_M2  M3_M2_4800
timestamp 1745462530
transform 1 0 3060 0 1 2705
box -3 -3 3 3
use M3_M2  M3_M2_4801
timestamp 1745462530
transform 1 0 3044 0 1 2725
box -3 -3 3 3
use M3_M2  M3_M2_4802
timestamp 1745462530
transform 1 0 2844 0 1 2725
box -3 -3 3 3
use M3_M2  M3_M2_4803
timestamp 1745462530
transform 1 0 2724 0 1 2725
box -3 -3 3 3
use M3_M2  M3_M2_4804
timestamp 1745462530
transform 1 0 3004 0 1 2755
box -3 -3 3 3
use M3_M2  M3_M2_4805
timestamp 1745462530
transform 1 0 2956 0 1 2755
box -3 -3 3 3
use M3_M2  M3_M2_4806
timestamp 1745462530
transform 1 0 4124 0 1 1265
box -3 -3 3 3
use M3_M2  M3_M2_4807
timestamp 1745462530
transform 1 0 4108 0 1 655
box -3 -3 3 3
use M3_M2  M3_M2_4808
timestamp 1745462530
transform 1 0 4028 0 1 1615
box -3 -3 3 3
use M3_M2  M3_M2_4809
timestamp 1745462530
transform 1 0 4012 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_4810
timestamp 1745462530
transform 1 0 3988 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_4811
timestamp 1745462530
transform 1 0 3988 0 1 1265
box -3 -3 3 3
use M3_M2  M3_M2_4812
timestamp 1745462530
transform 1 0 3972 0 1 2175
box -3 -3 3 3
use M3_M2  M3_M2_4813
timestamp 1745462530
transform 1 0 3972 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_4814
timestamp 1745462530
transform 1 0 3972 0 1 1935
box -3 -3 3 3
use M3_M2  M3_M2_4815
timestamp 1745462530
transform 1 0 3956 0 1 2445
box -3 -3 3 3
use M3_M2  M3_M2_4816
timestamp 1745462530
transform 1 0 3948 0 1 2665
box -3 -3 3 3
use M3_M2  M3_M2_4817
timestamp 1745462530
transform 1 0 3868 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_4818
timestamp 1745462530
transform 1 0 3868 0 1 85
box -3 -3 3 3
use M3_M2  M3_M2_4819
timestamp 1745462530
transform 1 0 3836 0 1 2445
box -3 -3 3 3
use M3_M2  M3_M2_4820
timestamp 1745462530
transform 1 0 3836 0 1 2175
box -3 -3 3 3
use M3_M2  M3_M2_4821
timestamp 1745462530
transform 1 0 3836 0 1 1935
box -3 -3 3 3
use M3_M2  M3_M2_4822
timestamp 1745462530
transform 1 0 3812 0 1 655
box -3 -3 3 3
use M3_M2  M3_M2_4823
timestamp 1745462530
transform 1 0 3804 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_4824
timestamp 1745462530
transform 1 0 3772 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_4825
timestamp 1745462530
transform 1 0 3764 0 1 2835
box -3 -3 3 3
use M3_M2  M3_M2_4826
timestamp 1745462530
transform 1 0 3764 0 1 2665
box -3 -3 3 3
use M3_M2  M3_M2_4827
timestamp 1745462530
transform 1 0 2868 0 1 2985
box -3 -3 3 3
use M3_M2  M3_M2_4828
timestamp 1745462530
transform 1 0 2868 0 1 2835
box -3 -3 3 3
use M3_M2  M3_M2_4829
timestamp 1745462530
transform 1 0 2660 0 1 2985
box -3 -3 3 3
use M3_M2  M3_M2_4830
timestamp 1745462530
transform 1 0 2532 0 1 3005
box -3 -3 3 3
use M3_M2  M3_M2_4831
timestamp 1745462530
transform 1 0 2532 0 1 2985
box -3 -3 3 3
use M3_M2  M3_M2_4832
timestamp 1745462530
transform 1 0 2468 0 1 3005
box -3 -3 3 3
use M3_M2  M3_M2_4833
timestamp 1745462530
transform 1 0 1284 0 1 85
box -3 -3 3 3
use M3_M2  M3_M2_4834
timestamp 1745462530
transform 1 0 1268 0 1 3005
box -3 -3 3 3
use M3_M2  M3_M2_4835
timestamp 1745462530
transform 1 0 2060 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_4836
timestamp 1745462530
transform 1 0 2060 0 1 1005
box -3 -3 3 3
use M3_M2  M3_M2_4837
timestamp 1745462530
transform 1 0 2044 0 1 1005
box -3 -3 3 3
use M3_M2  M3_M2_4838
timestamp 1745462530
transform 1 0 2044 0 1 665
box -3 -3 3 3
use M3_M2  M3_M2_4839
timestamp 1745462530
transform 1 0 2020 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_4840
timestamp 1745462530
transform 1 0 2020 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_4841
timestamp 1745462530
transform 1 0 1884 0 1 665
box -3 -3 3 3
use M3_M2  M3_M2_4842
timestamp 1745462530
transform 1 0 1452 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_4843
timestamp 1745462530
transform 1 0 1396 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_4844
timestamp 1745462530
transform 1 0 1364 0 1 2575
box -3 -3 3 3
use M3_M2  M3_M2_4845
timestamp 1745462530
transform 1 0 1284 0 1 665
box -3 -3 3 3
use M3_M2  M3_M2_4846
timestamp 1745462530
transform 1 0 1212 0 1 455
box -3 -3 3 3
use M3_M2  M3_M2_4847
timestamp 1745462530
transform 1 0 980 0 1 2565
box -3 -3 3 3
use M3_M2  M3_M2_4848
timestamp 1745462530
transform 1 0 980 0 1 2535
box -3 -3 3 3
use M3_M2  M3_M2_4849
timestamp 1745462530
transform 1 0 956 0 1 2535
box -3 -3 3 3
use M3_M2  M3_M2_4850
timestamp 1745462530
transform 1 0 956 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_4851
timestamp 1745462530
transform 1 0 724 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_4852
timestamp 1745462530
transform 1 0 724 0 1 2385
box -3 -3 3 3
use M3_M2  M3_M2_4853
timestamp 1745462530
transform 1 0 516 0 1 2455
box -3 -3 3 3
use M3_M2  M3_M2_4854
timestamp 1745462530
transform 1 0 500 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_4855
timestamp 1745462530
transform 1 0 500 0 1 455
box -3 -3 3 3
use M3_M2  M3_M2_4856
timestamp 1745462530
transform 1 0 460 0 1 2455
box -3 -3 3 3
use M3_M2  M3_M2_4857
timestamp 1745462530
transform 1 0 460 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_4858
timestamp 1745462530
transform 1 0 420 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_4859
timestamp 1745462530
transform 1 0 2612 0 1 1475
box -3 -3 3 3
use M3_M2  M3_M2_4860
timestamp 1745462530
transform 1 0 2572 0 1 2075
box -3 -3 3 3
use M3_M2  M3_M2_4861
timestamp 1745462530
transform 1 0 2436 0 1 2075
box -3 -3 3 3
use M3_M2  M3_M2_4862
timestamp 1745462530
transform 1 0 2436 0 1 1475
box -3 -3 3 3
use M3_M2  M3_M2_4863
timestamp 1745462530
transform 1 0 1740 0 1 2075
box -3 -3 3 3
use M3_M2  M3_M2_4864
timestamp 1745462530
transform 1 0 1372 0 1 2075
box -3 -3 3 3
use M3_M2  M3_M2_4865
timestamp 1745462530
transform 1 0 1348 0 1 2075
box -3 -3 3 3
use M3_M2  M3_M2_4866
timestamp 1745462530
transform 1 0 1348 0 1 2005
box -3 -3 3 3
use M3_M2  M3_M2_4867
timestamp 1745462530
transform 1 0 1300 0 1 1695
box -3 -3 3 3
use M3_M2  M3_M2_4868
timestamp 1745462530
transform 1 0 1292 0 1 2005
box -3 -3 3 3
use M3_M2  M3_M2_4869
timestamp 1745462530
transform 1 0 1284 0 1 1695
box -3 -3 3 3
use M3_M2  M3_M2_4870
timestamp 1745462530
transform 1 0 1468 0 1 2265
box -3 -3 3 3
use M3_M2  M3_M2_4871
timestamp 1745462530
transform 1 0 1412 0 1 2265
box -3 -3 3 3
use M3_M2  M3_M2_4872
timestamp 1745462530
transform 1 0 1380 0 1 2315
box -3 -3 3 3
use M3_M2  M3_M2_4873
timestamp 1745462530
transform 1 0 1124 0 1 3245
box -3 -3 3 3
use M3_M2  M3_M2_4874
timestamp 1745462530
transform 1 0 1116 0 1 3045
box -3 -3 3 3
use M3_M2  M3_M2_4875
timestamp 1745462530
transform 1 0 1100 0 1 3245
box -3 -3 3 3
use M3_M2  M3_M2_4876
timestamp 1745462530
transform 1 0 1100 0 1 2405
box -3 -3 3 3
use M3_M2  M3_M2_4877
timestamp 1745462530
transform 1 0 1100 0 1 2315
box -3 -3 3 3
use M3_M2  M3_M2_4878
timestamp 1745462530
transform 1 0 1076 0 1 3045
box -3 -3 3 3
use M3_M2  M3_M2_4879
timestamp 1745462530
transform 1 0 1068 0 1 2675
box -3 -3 3 3
use M3_M2  M3_M2_4880
timestamp 1745462530
transform 1 0 956 0 1 2405
box -3 -3 3 3
use M3_M2  M3_M2_4881
timestamp 1745462530
transform 1 0 948 0 1 2675
box -3 -3 3 3
use M3_M2  M3_M2_4882
timestamp 1745462530
transform 1 0 1324 0 1 1525
box -3 -3 3 3
use M3_M2  M3_M2_4883
timestamp 1745462530
transform 1 0 1308 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_4884
timestamp 1745462530
transform 1 0 1308 0 1 495
box -3 -3 3 3
use M3_M2  M3_M2_4885
timestamp 1745462530
transform 1 0 1260 0 1 495
box -3 -3 3 3
use M3_M2  M3_M2_4886
timestamp 1745462530
transform 1 0 996 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_4887
timestamp 1745462530
transform 1 0 980 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_4888
timestamp 1745462530
transform 1 0 740 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_4889
timestamp 1745462530
transform 1 0 540 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_4890
timestamp 1745462530
transform 1 0 540 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_4891
timestamp 1745462530
transform 1 0 540 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_4892
timestamp 1745462530
transform 1 0 468 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_4893
timestamp 1745462530
transform 1 0 460 0 1 865
box -3 -3 3 3
use M3_M2  M3_M2_4894
timestamp 1745462530
transform 1 0 460 0 1 675
box -3 -3 3 3
use M3_M2  M3_M2_4895
timestamp 1745462530
transform 1 0 460 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_4896
timestamp 1745462530
transform 1 0 436 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_4897
timestamp 1745462530
transform 1 0 348 0 1 865
box -3 -3 3 3
use M3_M2  M3_M2_4898
timestamp 1745462530
transform 1 0 348 0 1 675
box -3 -3 3 3
use M3_M2  M3_M2_4899
timestamp 1745462530
transform 1 0 300 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_4900
timestamp 1745462530
transform 1 0 300 0 1 865
box -3 -3 3 3
use M3_M2  M3_M2_4901
timestamp 1745462530
transform 1 0 252 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_4902
timestamp 1745462530
transform 1 0 244 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_4903
timestamp 1745462530
transform 1 0 124 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_4904
timestamp 1745462530
transform 1 0 124 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_4905
timestamp 1745462530
transform 1 0 3820 0 1 485
box -3 -3 3 3
use M3_M2  M3_M2_4906
timestamp 1745462530
transform 1 0 3796 0 1 1485
box -3 -3 3 3
use M3_M2  M3_M2_4907
timestamp 1745462530
transform 1 0 3604 0 1 495
box -3 -3 3 3
use M3_M2  M3_M2_4908
timestamp 1745462530
transform 1 0 3572 0 1 495
box -3 -3 3 3
use M3_M2  M3_M2_4909
timestamp 1745462530
transform 1 0 3532 0 1 495
box -3 -3 3 3
use M3_M2  M3_M2_4910
timestamp 1745462530
transform 1 0 2804 0 1 1475
box -3 -3 3 3
use M3_M2  M3_M2_4911
timestamp 1745462530
transform 1 0 2804 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_4912
timestamp 1745462530
transform 1 0 2676 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_4913
timestamp 1745462530
transform 1 0 2668 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_4914
timestamp 1745462530
transform 1 0 2652 0 1 1475
box -3 -3 3 3
use M3_M2  M3_M2_4915
timestamp 1745462530
transform 1 0 2636 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_4916
timestamp 1745462530
transform 1 0 2596 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_4917
timestamp 1745462530
transform 1 0 2004 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_4918
timestamp 1745462530
transform 1 0 1932 0 1 535
box -3 -3 3 3
use M3_M2  M3_M2_4919
timestamp 1745462530
transform 1 0 4140 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_4920
timestamp 1745462530
transform 1 0 4140 0 1 2045
box -3 -3 3 3
use M3_M2  M3_M2_4921
timestamp 1745462530
transform 1 0 4076 0 1 2045
box -3 -3 3 3
use M3_M2  M3_M2_4922
timestamp 1745462530
transform 1 0 4076 0 1 1895
box -3 -3 3 3
use M3_M2  M3_M2_4923
timestamp 1745462530
transform 1 0 4028 0 1 1895
box -3 -3 3 3
use M3_M2  M3_M2_4924
timestamp 1745462530
transform 1 0 3980 0 1 1895
box -3 -3 3 3
use M3_M2  M3_M2_4925
timestamp 1745462530
transform 1 0 3884 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_4926
timestamp 1745462530
transform 1 0 3868 0 1 1895
box -3 -3 3 3
use M3_M2  M3_M2_4927
timestamp 1745462530
transform 1 0 2604 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_4928
timestamp 1745462530
transform 1 0 1468 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_4929
timestamp 1745462530
transform 1 0 1396 0 1 2125
box -3 -3 3 3
use M3_M2  M3_M2_4930
timestamp 1745462530
transform 1 0 1396 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_4931
timestamp 1745462530
transform 1 0 1268 0 1 2185
box -3 -3 3 3
use M3_M2  M3_M2_4932
timestamp 1745462530
transform 1 0 1268 0 1 2125
box -3 -3 3 3
use M3_M2  M3_M2_4933
timestamp 1745462530
transform 1 0 1260 0 1 2365
box -3 -3 3 3
use M3_M2  M3_M2_4934
timestamp 1745462530
transform 1 0 1252 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_4935
timestamp 1745462530
transform 1 0 1252 0 1 2185
box -3 -3 3 3
use M3_M2  M3_M2_4936
timestamp 1745462530
transform 1 0 1244 0 1 2885
box -3 -3 3 3
use M3_M2  M3_M2_4937
timestamp 1745462530
transform 1 0 1244 0 1 2365
box -3 -3 3 3
use M3_M2  M3_M2_4938
timestamp 1745462530
transform 1 0 1236 0 1 3075
box -3 -3 3 3
use M3_M2  M3_M2_4939
timestamp 1745462530
transform 1 0 1228 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_4940
timestamp 1745462530
transform 1 0 1164 0 1 3075
box -3 -3 3 3
use M3_M2  M3_M2_4941
timestamp 1745462530
transform 1 0 1164 0 1 2885
box -3 -3 3 3
use M3_M2  M3_M2_4942
timestamp 1745462530
transform 1 0 1068 0 1 3075
box -3 -3 3 3
use M3_M2  M3_M2_4943
timestamp 1745462530
transform 1 0 1068 0 1 3025
box -3 -3 3 3
use M3_M2  M3_M2_4944
timestamp 1745462530
transform 1 0 1020 0 1 3025
box -3 -3 3 3
use M3_M2  M3_M2_4945
timestamp 1745462530
transform 1 0 1852 0 1 1655
box -3 -3 3 3
use M3_M2  M3_M2_4946
timestamp 1745462530
transform 1 0 1844 0 1 2245
box -3 -3 3 3
use M3_M2  M3_M2_4947
timestamp 1745462530
transform 1 0 1828 0 1 2245
box -3 -3 3 3
use M3_M2  M3_M2_4948
timestamp 1745462530
transform 1 0 1828 0 1 2125
box -3 -3 3 3
use M3_M2  M3_M2_4949
timestamp 1745462530
transform 1 0 1820 0 1 1655
box -3 -3 3 3
use M3_M2  M3_M2_4950
timestamp 1745462530
transform 1 0 1772 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_4951
timestamp 1745462530
transform 1 0 1772 0 1 1655
box -3 -3 3 3
use M3_M2  M3_M2_4952
timestamp 1745462530
transform 1 0 1764 0 1 2125
box -3 -3 3 3
use M3_M2  M3_M2_4953
timestamp 1745462530
transform 1 0 1676 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_4954
timestamp 1745462530
transform 1 0 1588 0 1 2245
box -3 -3 3 3
use M3_M2  M3_M2_4955
timestamp 1745462530
transform 1 0 3468 0 1 1085
box -3 -3 3 3
use M3_M2  M3_M2_4956
timestamp 1745462530
transform 1 0 3444 0 1 1085
box -3 -3 3 3
use M3_M2  M3_M2_4957
timestamp 1745462530
transform 1 0 3444 0 1 975
box -3 -3 3 3
use M3_M2  M3_M2_4958
timestamp 1745462530
transform 1 0 3396 0 1 1085
box -3 -3 3 3
use M3_M2  M3_M2_4959
timestamp 1745462530
transform 1 0 3276 0 1 975
box -3 -3 3 3
use M3_M2  M3_M2_4960
timestamp 1745462530
transform 1 0 3196 0 1 975
box -3 -3 3 3
use M3_M2  M3_M2_4961
timestamp 1745462530
transform 1 0 3132 0 1 2735
box -3 -3 3 3
use M3_M2  M3_M2_4962
timestamp 1745462530
transform 1 0 3084 0 1 2735
box -3 -3 3 3
use M3_M2  M3_M2_4963
timestamp 1745462530
transform 1 0 3084 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_4964
timestamp 1745462530
transform 1 0 3044 0 1 2735
box -3 -3 3 3
use M3_M2  M3_M2_4965
timestamp 1745462530
transform 1 0 3004 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_4966
timestamp 1745462530
transform 1 0 2988 0 1 1615
box -3 -3 3 3
use M3_M2  M3_M2_4967
timestamp 1745462530
transform 1 0 2932 0 1 1615
box -3 -3 3 3
use M3_M2  M3_M2_4968
timestamp 1745462530
transform 1 0 2932 0 1 1465
box -3 -3 3 3
use M3_M2  M3_M2_4969
timestamp 1745462530
transform 1 0 2868 0 1 1465
box -3 -3 3 3
use M3_M2  M3_M2_4970
timestamp 1745462530
transform 1 0 2868 0 1 975
box -3 -3 3 3
use M3_M2  M3_M2_4971
timestamp 1745462530
transform 1 0 2852 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_4972
timestamp 1745462530
transform 1 0 2820 0 1 975
box -3 -3 3 3
use M3_M2  M3_M2_4973
timestamp 1745462530
transform 1 0 2780 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_4974
timestamp 1745462530
transform 1 0 2780 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_4975
timestamp 1745462530
transform 1 0 2756 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_4976
timestamp 1745462530
transform 1 0 2756 0 1 975
box -3 -3 3 3
use M3_M2  M3_M2_4977
timestamp 1745462530
transform 1 0 2708 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_4978
timestamp 1745462530
transform 1 0 2708 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_4979
timestamp 1745462530
transform 1 0 2436 0 1 3035
box -3 -3 3 3
use M3_M2  M3_M2_4980
timestamp 1745462530
transform 1 0 2436 0 1 2735
box -3 -3 3 3
use M3_M2  M3_M2_4981
timestamp 1745462530
transform 1 0 2340 0 1 975
box -3 -3 3 3
use M3_M2  M3_M2_4982
timestamp 1745462530
transform 1 0 2172 0 1 3025
box -3 -3 3 3
use M3_M2  M3_M2_4983
timestamp 1745462530
transform 1 0 1572 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_4984
timestamp 1745462530
transform 1 0 1540 0 1 3025
box -3 -3 3 3
use M3_M2  M3_M2_4985
timestamp 1745462530
transform 1 0 1492 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_4986
timestamp 1745462530
transform 1 0 1492 0 1 975
box -3 -3 3 3
use M3_M2  M3_M2_4987
timestamp 1745462530
transform 1 0 1156 0 1 3025
box -3 -3 3 3
use M3_M2  M3_M2_4988
timestamp 1745462530
transform 1 0 1124 0 1 975
box -3 -3 3 3
use M3_M2  M3_M2_4989
timestamp 1745462530
transform 1 0 1076 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_4990
timestamp 1745462530
transform 1 0 1044 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_4991
timestamp 1745462530
transform 1 0 1020 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_4992
timestamp 1745462530
transform 1 0 3820 0 1 3885
box -3 -3 3 3
use M3_M2  M3_M2_4993
timestamp 1745462530
transform 1 0 3180 0 1 3885
box -3 -3 3 3
use M3_M2  M3_M2_4994
timestamp 1745462530
transform 1 0 3180 0 1 3815
box -3 -3 3 3
use M3_M2  M3_M2_4995
timestamp 1745462530
transform 1 0 2820 0 1 3985
box -3 -3 3 3
use M3_M2  M3_M2_4996
timestamp 1745462530
transform 1 0 2820 0 1 3815
box -3 -3 3 3
use M3_M2  M3_M2_4997
timestamp 1745462530
transform 1 0 2820 0 1 3765
box -3 -3 3 3
use M3_M2  M3_M2_4998
timestamp 1745462530
transform 1 0 2788 0 1 4325
box -3 -3 3 3
use M3_M2  M3_M2_4999
timestamp 1745462530
transform 1 0 2788 0 1 3985
box -3 -3 3 3
use M3_M2  M3_M2_5000
timestamp 1745462530
transform 1 0 2780 0 1 3765
box -3 -3 3 3
use M3_M2  M3_M2_5001
timestamp 1745462530
transform 1 0 2164 0 1 4115
box -3 -3 3 3
use M3_M2  M3_M2_5002
timestamp 1745462530
transform 1 0 2164 0 1 3945
box -3 -3 3 3
use M3_M2  M3_M2_5003
timestamp 1745462530
transform 1 0 2100 0 1 4115
box -3 -3 3 3
use M3_M2  M3_M2_5004
timestamp 1745462530
transform 1 0 2092 0 1 4325
box -3 -3 3 3
use M3_M2  M3_M2_5005
timestamp 1745462530
transform 1 0 1580 0 1 3945
box -3 -3 3 3
use M3_M2  M3_M2_5006
timestamp 1745462530
transform 1 0 4212 0 1 3195
box -3 -3 3 3
use M3_M2  M3_M2_5007
timestamp 1745462530
transform 1 0 4196 0 1 3195
box -3 -3 3 3
use M3_M2  M3_M2_5008
timestamp 1745462530
transform 1 0 4036 0 1 3205
box -3 -3 3 3
use M3_M2  M3_M2_5009
timestamp 1745462530
transform 1 0 4020 0 1 3475
box -3 -3 3 3
use M3_M2  M3_M2_5010
timestamp 1745462530
transform 1 0 4004 0 1 3475
box -3 -3 3 3
use M3_M2  M3_M2_5011
timestamp 1745462530
transform 1 0 3996 0 1 3635
box -3 -3 3 3
use M3_M2  M3_M2_5012
timestamp 1745462530
transform 1 0 3940 0 1 3205
box -3 -3 3 3
use M3_M2  M3_M2_5013
timestamp 1745462530
transform 1 0 3884 0 1 3905
box -3 -3 3 3
use M3_M2  M3_M2_5014
timestamp 1745462530
transform 1 0 3884 0 1 3635
box -3 -3 3 3
use M3_M2  M3_M2_5015
timestamp 1745462530
transform 1 0 2172 0 1 3975
box -3 -3 3 3
use M3_M2  M3_M2_5016
timestamp 1745462530
transform 1 0 2172 0 1 3905
box -3 -3 3 3
use M3_M2  M3_M2_5017
timestamp 1745462530
transform 1 0 1764 0 1 3975
box -3 -3 3 3
use M3_M2  M3_M2_5018
timestamp 1745462530
transform 1 0 1764 0 1 3915
box -3 -3 3 3
use M3_M2  M3_M2_5019
timestamp 1745462530
transform 1 0 1700 0 1 3915
box -3 -3 3 3
use M3_M2  M3_M2_5020
timestamp 1745462530
transform 1 0 1644 0 1 3915
box -3 -3 3 3
use M3_M2  M3_M2_5021
timestamp 1745462530
transform 1 0 4132 0 1 3415
box -3 -3 3 3
use M3_M2  M3_M2_5022
timestamp 1745462530
transform 1 0 4044 0 1 3595
box -3 -3 3 3
use M3_M2  M3_M2_5023
timestamp 1745462530
transform 1 0 4044 0 1 3525
box -3 -3 3 3
use M3_M2  M3_M2_5024
timestamp 1745462530
transform 1 0 3972 0 1 3415
box -3 -3 3 3
use M3_M2  M3_M2_5025
timestamp 1745462530
transform 1 0 3956 0 1 3915
box -3 -3 3 3
use M3_M2  M3_M2_5026
timestamp 1745462530
transform 1 0 3956 0 1 3595
box -3 -3 3 3
use M3_M2  M3_M2_5027
timestamp 1745462530
transform 1 0 3948 0 1 3525
box -3 -3 3 3
use M3_M2  M3_M2_5028
timestamp 1745462530
transform 1 0 2852 0 1 3925
box -3 -3 3 3
use M3_M2  M3_M2_5029
timestamp 1745462530
transform 1 0 2676 0 1 3925
box -3 -3 3 3
use M3_M2  M3_M2_5030
timestamp 1745462530
transform 1 0 2148 0 1 3925
box -3 -3 3 3
use M3_M2  M3_M2_5031
timestamp 1745462530
transform 1 0 2060 0 1 3955
box -3 -3 3 3
use M3_M2  M3_M2_5032
timestamp 1745462530
transform 1 0 2060 0 1 3925
box -3 -3 3 3
use M3_M2  M3_M2_5033
timestamp 1745462530
transform 1 0 2028 0 1 3925
box -3 -3 3 3
use M3_M2  M3_M2_5034
timestamp 1745462530
transform 1 0 2028 0 1 3705
box -3 -3 3 3
use M3_M2  M3_M2_5035
timestamp 1745462530
transform 1 0 2012 0 1 3955
box -3 -3 3 3
use M3_M2  M3_M2_5036
timestamp 1745462530
transform 1 0 1972 0 1 3705
box -3 -3 3 3
use M3_M2  M3_M2_5037
timestamp 1745462530
transform 1 0 1932 0 1 3955
box -3 -3 3 3
use M3_M2  M3_M2_5038
timestamp 1745462530
transform 1 0 1924 0 1 3925
box -3 -3 3 3
use M3_M2  M3_M2_5039
timestamp 1745462530
transform 1 0 1860 0 1 3925
box -3 -3 3 3
use M3_M2  M3_M2_5040
timestamp 1745462530
transform 1 0 4308 0 1 3665
box -3 -3 3 3
use M3_M2  M3_M2_5041
timestamp 1745462530
transform 1 0 4300 0 1 3775
box -3 -3 3 3
use M3_M2  M3_M2_5042
timestamp 1745462530
transform 1 0 4236 0 1 3655
box -3 -3 3 3
use M3_M2  M3_M2_5043
timestamp 1745462530
transform 1 0 4212 0 1 3775
box -3 -3 3 3
use M3_M2  M3_M2_5044
timestamp 1745462530
transform 1 0 3868 0 1 3655
box -3 -3 3 3
use M3_M2  M3_M2_5045
timestamp 1745462530
transform 1 0 3860 0 1 3985
box -3 -3 3 3
use M3_M2  M3_M2_5046
timestamp 1745462530
transform 1 0 3852 0 1 4095
box -3 -3 3 3
use M3_M2  M3_M2_5047
timestamp 1745462530
transform 1 0 3756 0 1 3985
box -3 -3 3 3
use M3_M2  M3_M2_5048
timestamp 1745462530
transform 1 0 3716 0 1 3985
box -3 -3 3 3
use M3_M2  M3_M2_5049
timestamp 1745462530
transform 1 0 3708 0 1 4095
box -3 -3 3 3
use M3_M2  M3_M2_5050
timestamp 1745462530
transform 1 0 3708 0 1 3935
box -3 -3 3 3
use M3_M2  M3_M2_5051
timestamp 1745462530
transform 1 0 3676 0 1 3935
box -3 -3 3 3
use M3_M2  M3_M2_5052
timestamp 1745462530
transform 1 0 2980 0 1 4095
box -3 -3 3 3
use M3_M2  M3_M2_5053
timestamp 1745462530
transform 1 0 2908 0 1 4095
box -3 -3 3 3
use M3_M2  M3_M2_5054
timestamp 1745462530
transform 1 0 2588 0 1 4105
box -3 -3 3 3
use M3_M2  M3_M2_5055
timestamp 1745462530
transform 1 0 2484 0 1 4105
box -3 -3 3 3
use M3_M2  M3_M2_5056
timestamp 1745462530
transform 1 0 2284 0 1 4105
box -3 -3 3 3
use M3_M2  M3_M2_5057
timestamp 1745462530
transform 1 0 3500 0 1 3985
box -3 -3 3 3
use M3_M2  M3_M2_5058
timestamp 1745462530
transform 1 0 3484 0 1 4185
box -3 -3 3 3
use M3_M2  M3_M2_5059
timestamp 1745462530
transform 1 0 3484 0 1 3985
box -3 -3 3 3
use M3_M2  M3_M2_5060
timestamp 1745462530
transform 1 0 3380 0 1 4185
box -3 -3 3 3
use M3_M2  M3_M2_5061
timestamp 1745462530
transform 1 0 3372 0 1 4125
box -3 -3 3 3
use M3_M2  M3_M2_5062
timestamp 1745462530
transform 1 0 3228 0 1 4145
box -3 -3 3 3
use M3_M2  M3_M2_5063
timestamp 1745462530
transform 1 0 3172 0 1 4145
box -3 -3 3 3
use M3_M2  M3_M2_5064
timestamp 1745462530
transform 1 0 3012 0 1 4145
box -3 -3 3 3
use M3_M2  M3_M2_5065
timestamp 1745462530
transform 1 0 2732 0 1 4125
box -3 -3 3 3
use M3_M2  M3_M2_5066
timestamp 1745462530
transform 1 0 2644 0 1 4125
box -3 -3 3 3
use M3_M2  M3_M2_5067
timestamp 1745462530
transform 1 0 2404 0 1 4125
box -3 -3 3 3
use M3_M2  M3_M2_5068
timestamp 1745462530
transform 1 0 2380 0 1 4125
box -3 -3 3 3
use M3_M2  M3_M2_5069
timestamp 1745462530
transform 1 0 2372 0 1 3945
box -3 -3 3 3
use M3_M2  M3_M2_5070
timestamp 1745462530
transform 1 0 2220 0 1 4125
box -3 -3 3 3
use M3_M2  M3_M2_5071
timestamp 1745462530
transform 1 0 2212 0 1 3945
box -3 -3 3 3
use M3_M2  M3_M2_5072
timestamp 1745462530
transform 1 0 2164 0 1 4125
box -3 -3 3 3
use M3_M2  M3_M2_5073
timestamp 1745462530
transform 1 0 3596 0 1 3965
box -3 -3 3 3
use M3_M2  M3_M2_5074
timestamp 1745462530
transform 1 0 3588 0 1 3725
box -3 -3 3 3
use M3_M2  M3_M2_5075
timestamp 1745462530
transform 1 0 3556 0 1 3965
box -3 -3 3 3
use M3_M2  M3_M2_5076
timestamp 1745462530
transform 1 0 3548 0 1 3725
box -3 -3 3 3
use M3_M2  M3_M2_5077
timestamp 1745462530
transform 1 0 3356 0 1 3965
box -3 -3 3 3
use M3_M2  M3_M2_5078
timestamp 1745462530
transform 1 0 3276 0 1 3965
box -3 -3 3 3
use M3_M2  M3_M2_5079
timestamp 1745462530
transform 1 0 3140 0 1 3945
box -3 -3 3 3
use M3_M2  M3_M2_5080
timestamp 1745462530
transform 1 0 3084 0 1 3945
box -3 -3 3 3
use M3_M2  M3_M2_5081
timestamp 1745462530
transform 1 0 2836 0 1 3965
box -3 -3 3 3
use M3_M2  M3_M2_5082
timestamp 1745462530
transform 1 0 2836 0 1 3945
box -3 -3 3 3
use M3_M2  M3_M2_5083
timestamp 1745462530
transform 1 0 2380 0 1 3965
box -3 -3 3 3
use M3_M2  M3_M2_5084
timestamp 1745462530
transform 1 0 2380 0 1 3845
box -3 -3 3 3
use M3_M2  M3_M2_5085
timestamp 1745462530
transform 1 0 2260 0 1 3835
box -3 -3 3 3
use M3_M2  M3_M2_5086
timestamp 1745462530
transform 1 0 2068 0 1 3965
box -3 -3 3 3
use M3_M2  M3_M2_5087
timestamp 1745462530
transform 1 0 804 0 1 4095
box -3 -3 3 3
use M3_M2  M3_M2_5088
timestamp 1745462530
transform 1 0 628 0 1 4095
box -3 -3 3 3
use M3_M2  M3_M2_5089
timestamp 1745462530
transform 1 0 4156 0 1 4315
box -3 -3 3 3
use M3_M2  M3_M2_5090
timestamp 1745462530
transform 1 0 4156 0 1 4085
box -3 -3 3 3
use M3_M2  M3_M2_5091
timestamp 1745462530
transform 1 0 4100 0 1 4315
box -3 -3 3 3
use M3_M2  M3_M2_5092
timestamp 1745462530
transform 1 0 4068 0 1 4095
box -3 -3 3 3
use M3_M2  M3_M2_5093
timestamp 1745462530
transform 1 0 3988 0 1 4095
box -3 -3 3 3
use M3_M2  M3_M2_5094
timestamp 1745462530
transform 1 0 2908 0 1 4315
box -3 -3 3 3
use M3_M2  M3_M2_5095
timestamp 1745462530
transform 1 0 2908 0 1 4265
box -3 -3 3 3
use M3_M2  M3_M2_5096
timestamp 1745462530
transform 1 0 2668 0 1 4265
box -3 -3 3 3
use M3_M2  M3_M2_5097
timestamp 1745462530
transform 1 0 1940 0 1 4265
box -3 -3 3 3
use M3_M2  M3_M2_5098
timestamp 1745462530
transform 1 0 1940 0 1 4245
box -3 -3 3 3
use M3_M2  M3_M2_5099
timestamp 1745462530
transform 1 0 1892 0 1 4005
box -3 -3 3 3
use M3_M2  M3_M2_5100
timestamp 1745462530
transform 1 0 1812 0 1 4005
box -3 -3 3 3
use M3_M2  M3_M2_5101
timestamp 1745462530
transform 1 0 1804 0 1 4245
box -3 -3 3 3
use M3_M2  M3_M2_5102
timestamp 1745462530
transform 1 0 1348 0 1 4155
box -3 -3 3 3
use M3_M2  M3_M2_5103
timestamp 1745462530
transform 1 0 1348 0 1 4005
box -3 -3 3 3
use M3_M2  M3_M2_5104
timestamp 1745462530
transform 1 0 1324 0 1 4025
box -3 -3 3 3
use M3_M2  M3_M2_5105
timestamp 1745462530
transform 1 0 1260 0 1 4025
box -3 -3 3 3
use M3_M2  M3_M2_5106
timestamp 1745462530
transform 1 0 1084 0 1 4155
box -3 -3 3 3
use M3_M2  M3_M2_5107
timestamp 1745462530
transform 1 0 884 0 1 4155
box -3 -3 3 3
use M3_M2  M3_M2_5108
timestamp 1745462530
transform 1 0 1156 0 1 3345
box -3 -3 3 3
use M3_M2  M3_M2_5109
timestamp 1745462530
transform 1 0 1132 0 1 3345
box -3 -3 3 3
use M3_M2  M3_M2_5110
timestamp 1745462530
transform 1 0 1012 0 1 3345
box -3 -3 3 3
use M3_M2  M3_M2_5111
timestamp 1745462530
transform 1 0 916 0 1 3345
box -3 -3 3 3
use M3_M2  M3_M2_5112
timestamp 1745462530
transform 1 0 3548 0 1 4035
box -3 -3 3 3
use M3_M2  M3_M2_5113
timestamp 1745462530
transform 1 0 3524 0 1 4035
box -3 -3 3 3
use M3_M2  M3_M2_5114
timestamp 1745462530
transform 1 0 3420 0 1 4035
box -3 -3 3 3
use M3_M2  M3_M2_5115
timestamp 1745462530
transform 1 0 3044 0 1 4035
box -3 -3 3 3
use M3_M2  M3_M2_5116
timestamp 1745462530
transform 1 0 2668 0 1 4035
box -3 -3 3 3
use M3_M2  M3_M2_5117
timestamp 1745462530
transform 1 0 2556 0 1 4115
box -3 -3 3 3
use M3_M2  M3_M2_5118
timestamp 1745462530
transform 1 0 2556 0 1 4035
box -3 -3 3 3
use M3_M2  M3_M2_5119
timestamp 1745462530
transform 1 0 2540 0 1 4035
box -3 -3 3 3
use M3_M2  M3_M2_5120
timestamp 1745462530
transform 1 0 2340 0 1 4115
box -3 -3 3 3
use M3_M2  M3_M2_5121
timestamp 1745462530
transform 1 0 2228 0 1 4115
box -3 -3 3 3
use M3_M2  M3_M2_5122
timestamp 1745462530
transform 1 0 2212 0 1 3725
box -3 -3 3 3
use M3_M2  M3_M2_5123
timestamp 1745462530
transform 1 0 2180 0 1 3725
box -3 -3 3 3
use M3_M2  M3_M2_5124
timestamp 1745462530
transform 1 0 3556 0 1 3835
box -3 -3 3 3
use M3_M2  M3_M2_5125
timestamp 1745462530
transform 1 0 3508 0 1 3835
box -3 -3 3 3
use M3_M2  M3_M2_5126
timestamp 1745462530
transform 1 0 3492 0 1 3875
box -3 -3 3 3
use M3_M2  M3_M2_5127
timestamp 1745462530
transform 1 0 3492 0 1 3835
box -3 -3 3 3
use M3_M2  M3_M2_5128
timestamp 1745462530
transform 1 0 3268 0 1 3915
box -3 -3 3 3
use M3_M2  M3_M2_5129
timestamp 1745462530
transform 1 0 3268 0 1 3875
box -3 -3 3 3
use M3_M2  M3_M2_5130
timestamp 1745462530
transform 1 0 3236 0 1 3915
box -3 -3 3 3
use M3_M2  M3_M2_5131
timestamp 1745462530
transform 1 0 3236 0 1 3895
box -3 -3 3 3
use M3_M2  M3_M2_5132
timestamp 1745462530
transform 1 0 3068 0 1 3895
box -3 -3 3 3
use M3_M2  M3_M2_5133
timestamp 1745462530
transform 1 0 2796 0 1 3895
box -3 -3 3 3
use M3_M2  M3_M2_5134
timestamp 1745462530
transform 1 0 2548 0 1 3895
box -3 -3 3 3
use M3_M2  M3_M2_5135
timestamp 1745462530
transform 1 0 2428 0 1 3895
box -3 -3 3 3
use M3_M2  M3_M2_5136
timestamp 1745462530
transform 1 0 2428 0 1 3865
box -3 -3 3 3
use M3_M2  M3_M2_5137
timestamp 1745462530
transform 1 0 2364 0 1 3865
box -3 -3 3 3
use M3_M2  M3_M2_5138
timestamp 1745462530
transform 1 0 2364 0 1 3745
box -3 -3 3 3
use M3_M2  M3_M2_5139
timestamp 1745462530
transform 1 0 2356 0 1 3955
box -3 -3 3 3
use M3_M2  M3_M2_5140
timestamp 1745462530
transform 1 0 2188 0 1 3955
box -3 -3 3 3
use M3_M2  M3_M2_5141
timestamp 1745462530
transform 1 0 2140 0 1 3745
box -3 -3 3 3
use M3_M2  M3_M2_5142
timestamp 1745462530
transform 1 0 3076 0 1 3575
box -3 -3 3 3
use M3_M2  M3_M2_5143
timestamp 1745462530
transform 1 0 3044 0 1 3335
box -3 -3 3 3
use M3_M2  M3_M2_5144
timestamp 1745462530
transform 1 0 3028 0 1 3575
box -3 -3 3 3
use M3_M2  M3_M2_5145
timestamp 1745462530
transform 1 0 3004 0 1 3845
box -3 -3 3 3
use M3_M2  M3_M2_5146
timestamp 1745462530
transform 1 0 2996 0 1 3575
box -3 -3 3 3
use M3_M2  M3_M2_5147
timestamp 1745462530
transform 1 0 2948 0 1 3335
box -3 -3 3 3
use M3_M2  M3_M2_5148
timestamp 1745462530
transform 1 0 2900 0 1 3145
box -3 -3 3 3
use M3_M2  M3_M2_5149
timestamp 1745462530
transform 1 0 2764 0 1 3845
box -3 -3 3 3
use M3_M2  M3_M2_5150
timestamp 1745462530
transform 1 0 2036 0 1 3145
box -3 -3 3 3
use M3_M2  M3_M2_5151
timestamp 1745462530
transform 1 0 3588 0 1 3495
box -3 -3 3 3
use M3_M2  M3_M2_5152
timestamp 1745462530
transform 1 0 3572 0 1 3565
box -3 -3 3 3
use M3_M2  M3_M2_5153
timestamp 1745462530
transform 1 0 3540 0 1 3495
box -3 -3 3 3
use M3_M2  M3_M2_5154
timestamp 1745462530
transform 1 0 3540 0 1 3385
box -3 -3 3 3
use M3_M2  M3_M2_5155
timestamp 1745462530
transform 1 0 3540 0 1 3305
box -3 -3 3 3
use M3_M2  M3_M2_5156
timestamp 1745462530
transform 1 0 3532 0 1 3635
box -3 -3 3 3
use M3_M2  M3_M2_5157
timestamp 1745462530
transform 1 0 3532 0 1 3565
box -3 -3 3 3
use M3_M2  M3_M2_5158
timestamp 1745462530
transform 1 0 3516 0 1 3305
box -3 -3 3 3
use M3_M2  M3_M2_5159
timestamp 1745462530
transform 1 0 3508 0 1 3635
box -3 -3 3 3
use M3_M2  M3_M2_5160
timestamp 1745462530
transform 1 0 3508 0 1 3125
box -3 -3 3 3
use M3_M2  M3_M2_5161
timestamp 1745462530
transform 1 0 3476 0 1 3375
box -3 -3 3 3
use M3_M2  M3_M2_5162
timestamp 1745462530
transform 1 0 3356 0 1 3575
box -3 -3 3 3
use M3_M2  M3_M2_5163
timestamp 1745462530
transform 1 0 3348 0 1 3535
box -3 -3 3 3
use M3_M2  M3_M2_5164
timestamp 1745462530
transform 1 0 3292 0 1 3125
box -3 -3 3 3
use M3_M2  M3_M2_5165
timestamp 1745462530
transform 1 0 3276 0 1 3535
box -3 -3 3 3
use M3_M2  M3_M2_5166
timestamp 1745462530
transform 1 0 3188 0 1 3125
box -3 -3 3 3
use M3_M2  M3_M2_5167
timestamp 1745462530
transform 1 0 2428 0 1 3125
box -3 -3 3 3
use M3_M2  M3_M2_5168
timestamp 1745462530
transform 1 0 2668 0 1 3465
box -3 -3 3 3
use M3_M2  M3_M2_5169
timestamp 1745462530
transform 1 0 2628 0 1 3555
box -3 -3 3 3
use M3_M2  M3_M2_5170
timestamp 1745462530
transform 1 0 2628 0 1 3465
box -3 -3 3 3
use M3_M2  M3_M2_5171
timestamp 1745462530
transform 1 0 2564 0 1 3255
box -3 -3 3 3
use M3_M2  M3_M2_5172
timestamp 1745462530
transform 1 0 2524 0 1 3255
box -3 -3 3 3
use M3_M2  M3_M2_5173
timestamp 1745462530
transform 1 0 2516 0 1 3565
box -3 -3 3 3
use M3_M2  M3_M2_5174
timestamp 1745462530
transform 1 0 2484 0 1 3565
box -3 -3 3 3
use M3_M2  M3_M2_5175
timestamp 1745462530
transform 1 0 2444 0 1 3255
box -3 -3 3 3
use M3_M2  M3_M2_5176
timestamp 1745462530
transform 1 0 2292 0 1 3255
box -3 -3 3 3
use M3_M2  M3_M2_5177
timestamp 1745462530
transform 1 0 3492 0 1 3595
box -3 -3 3 3
use M3_M2  M3_M2_5178
timestamp 1745462530
transform 1 0 3444 0 1 3405
box -3 -3 3 3
use M3_M2  M3_M2_5179
timestamp 1745462530
transform 1 0 3396 0 1 3095
box -3 -3 3 3
use M3_M2  M3_M2_5180
timestamp 1745462530
transform 1 0 3372 0 1 3405
box -3 -3 3 3
use M3_M2  M3_M2_5181
timestamp 1745462530
transform 1 0 3372 0 1 3295
box -3 -3 3 3
use M3_M2  M3_M2_5182
timestamp 1745462530
transform 1 0 3356 0 1 3095
box -3 -3 3 3
use M3_M2  M3_M2_5183
timestamp 1745462530
transform 1 0 3348 0 1 3295
box -3 -3 3 3
use M3_M2  M3_M2_5184
timestamp 1745462530
transform 1 0 3236 0 1 3095
box -3 -3 3 3
use M3_M2  M3_M2_5185
timestamp 1745462530
transform 1 0 3204 0 1 3595
box -3 -3 3 3
use M3_M2  M3_M2_5186
timestamp 1745462530
transform 1 0 3148 0 1 3485
box -3 -3 3 3
use M3_M2  M3_M2_5187
timestamp 1745462530
transform 1 0 3148 0 1 3095
box -3 -3 3 3
use M3_M2  M3_M2_5188
timestamp 1745462530
transform 1 0 3148 0 1 3075
box -3 -3 3 3
use M3_M2  M3_M2_5189
timestamp 1745462530
transform 1 0 3132 0 1 3595
box -3 -3 3 3
use M3_M2  M3_M2_5190
timestamp 1745462530
transform 1 0 3116 0 1 3485
box -3 -3 3 3
use M3_M2  M3_M2_5191
timestamp 1745462530
transform 1 0 2060 0 1 3075
box -3 -3 3 3
use M3_M2  M3_M2_5192
timestamp 1745462530
transform 1 0 3948 0 1 1285
box -3 -3 3 3
use M3_M2  M3_M2_5193
timestamp 1745462530
transform 1 0 3900 0 1 1285
box -3 -3 3 3
use M3_M2  M3_M2_5194
timestamp 1745462530
transform 1 0 3692 0 1 1285
box -3 -3 3 3
use M3_M2  M3_M2_5195
timestamp 1745462530
transform 1 0 3564 0 1 1285
box -3 -3 3 3
use M3_M2  M3_M2_5196
timestamp 1745462530
transform 1 0 3364 0 1 1285
box -3 -3 3 3
use M3_M2  M3_M2_5197
timestamp 1745462530
transform 1 0 3140 0 1 1285
box -3 -3 3 3
use M3_M2  M3_M2_5198
timestamp 1745462530
transform 1 0 3028 0 1 1285
box -3 -3 3 3
use M3_M2  M3_M2_5199
timestamp 1745462530
transform 1 0 2756 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_5200
timestamp 1745462530
transform 1 0 2756 0 1 1285
box -3 -3 3 3
use M3_M2  M3_M2_5201
timestamp 1745462530
transform 1 0 2556 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_5202
timestamp 1745462530
transform 1 0 2476 0 1 1435
box -3 -3 3 3
use M3_M2  M3_M2_5203
timestamp 1745462530
transform 1 0 2476 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_5204
timestamp 1745462530
transform 1 0 2348 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_5205
timestamp 1745462530
transform 1 0 2244 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_5206
timestamp 1745462530
transform 1 0 3100 0 1 2275
box -3 -3 3 3
use M3_M2  M3_M2_5207
timestamp 1745462530
transform 1 0 3076 0 1 2275
box -3 -3 3 3
use M3_M2  M3_M2_5208
timestamp 1745462530
transform 1 0 3052 0 1 2295
box -3 -3 3 3
use M3_M2  M3_M2_5209
timestamp 1745462530
transform 1 0 3052 0 1 2275
box -3 -3 3 3
use M3_M2  M3_M2_5210
timestamp 1745462530
transform 1 0 2996 0 1 2295
box -3 -3 3 3
use M3_M2  M3_M2_5211
timestamp 1745462530
transform 1 0 2956 0 1 2295
box -3 -3 3 3
use M3_M2  M3_M2_5212
timestamp 1745462530
transform 1 0 2924 0 1 1685
box -3 -3 3 3
use M3_M2  M3_M2_5213
timestamp 1745462530
transform 1 0 2916 0 1 2295
box -3 -3 3 3
use M3_M2  M3_M2_5214
timestamp 1745462530
transform 1 0 2916 0 1 2275
box -3 -3 3 3
use M3_M2  M3_M2_5215
timestamp 1745462530
transform 1 0 2748 0 1 2275
box -3 -3 3 3
use M3_M2  M3_M2_5216
timestamp 1745462530
transform 1 0 2748 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_5217
timestamp 1745462530
transform 1 0 2692 0 1 2075
box -3 -3 3 3
use M3_M2  M3_M2_5218
timestamp 1745462530
transform 1 0 2692 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_5219
timestamp 1745462530
transform 1 0 2684 0 1 1685
box -3 -3 3 3
use M3_M2  M3_M2_5220
timestamp 1745462530
transform 1 0 2652 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_5221
timestamp 1745462530
transform 1 0 2652 0 1 1685
box -3 -3 3 3
use M3_M2  M3_M2_5222
timestamp 1745462530
transform 1 0 2564 0 1 2065
box -3 -3 3 3
use M3_M2  M3_M2_5223
timestamp 1745462530
transform 1 0 2244 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_5224
timestamp 1745462530
transform 1 0 2084 0 1 1835
box -3 -3 3 3
use M3_M2  M3_M2_5225
timestamp 1745462530
transform 1 0 2036 0 1 1835
box -3 -3 3 3
use M3_M2  M3_M2_5226
timestamp 1745462530
transform 1 0 1940 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_5227
timestamp 1745462530
transform 1 0 1588 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_5228
timestamp 1745462530
transform 1 0 1588 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_5229
timestamp 1745462530
transform 1 0 1540 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_5230
timestamp 1745462530
transform 1 0 1380 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_5231
timestamp 1745462530
transform 1 0 1284 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_5232
timestamp 1745462530
transform 1 0 1180 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_5233
timestamp 1745462530
transform 1 0 1044 0 1 1815
box -3 -3 3 3
use M3_M2  M3_M2_5234
timestamp 1745462530
transform 1 0 1020 0 1 1815
box -3 -3 3 3
use M3_M2  M3_M2_5235
timestamp 1745462530
transform 1 0 1012 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_5236
timestamp 1745462530
transform 1 0 932 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_5237
timestamp 1745462530
transform 1 0 2140 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_5238
timestamp 1745462530
transform 1 0 2116 0 1 1485
box -3 -3 3 3
use M3_M2  M3_M2_5239
timestamp 1745462530
transform 1 0 2116 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_5240
timestamp 1745462530
transform 1 0 1916 0 1 1485
box -3 -3 3 3
use M3_M2  M3_M2_5241
timestamp 1745462530
transform 1 0 1740 0 1 1495
box -3 -3 3 3
use M3_M2  M3_M2_5242
timestamp 1745462530
transform 1 0 1740 0 1 1485
box -3 -3 3 3
use M3_M2  M3_M2_5243
timestamp 1745462530
transform 1 0 1532 0 1 1495
box -3 -3 3 3
use M3_M2  M3_M2_5244
timestamp 1745462530
transform 1 0 1284 0 1 1495
box -3 -3 3 3
use M3_M2  M3_M2_5245
timestamp 1745462530
transform 1 0 1284 0 1 1475
box -3 -3 3 3
use M3_M2  M3_M2_5246
timestamp 1745462530
transform 1 0 1244 0 1 1475
box -3 -3 3 3
use M3_M2  M3_M2_5247
timestamp 1745462530
transform 1 0 1212 0 1 1475
box -3 -3 3 3
use M3_M2  M3_M2_5248
timestamp 1745462530
transform 1 0 1212 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_5249
timestamp 1745462530
transform 1 0 1180 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_5250
timestamp 1745462530
transform 1 0 1132 0 1 1475
box -3 -3 3 3
use M3_M2  M3_M2_5251
timestamp 1745462530
transform 1 0 1076 0 1 1475
box -3 -3 3 3
use M3_M2  M3_M2_5252
timestamp 1745462530
transform 1 0 1044 0 1 1475
box -3 -3 3 3
use M3_M2  M3_M2_5253
timestamp 1745462530
transform 1 0 1044 0 1 1415
box -3 -3 3 3
use M3_M2  M3_M2_5254
timestamp 1745462530
transform 1 0 964 0 1 1415
box -3 -3 3 3
use M3_M2  M3_M2_5255
timestamp 1745462530
transform 1 0 500 0 1 3555
box -3 -3 3 3
use M3_M2  M3_M2_5256
timestamp 1745462530
transform 1 0 340 0 1 3555
box -3 -3 3 3
use M3_M2  M3_M2_5257
timestamp 1745462530
transform 1 0 284 0 1 3555
box -3 -3 3 3
use M3_M2  M3_M2_5258
timestamp 1745462530
transform 1 0 252 0 1 3555
box -3 -3 3 3
use M3_M2  M3_M2_5259
timestamp 1745462530
transform 1 0 220 0 1 3555
box -3 -3 3 3
use M3_M2  M3_M2_5260
timestamp 1745462530
transform 1 0 284 0 1 3525
box -3 -3 3 3
use M3_M2  M3_M2_5261
timestamp 1745462530
transform 1 0 164 0 1 3525
box -3 -3 3 3
use M3_M2  M3_M2_5262
timestamp 1745462530
transform 1 0 412 0 1 3505
box -3 -3 3 3
use M3_M2  M3_M2_5263
timestamp 1745462530
transform 1 0 356 0 1 3505
box -3 -3 3 3
use M3_M2  M3_M2_5264
timestamp 1745462530
transform 1 0 276 0 1 3435
box -3 -3 3 3
use M3_M2  M3_M2_5265
timestamp 1745462530
transform 1 0 268 0 1 3605
box -3 -3 3 3
use M3_M2  M3_M2_5266
timestamp 1745462530
transform 1 0 236 0 1 3425
box -3 -3 3 3
use M3_M2  M3_M2_5267
timestamp 1745462530
transform 1 0 196 0 1 3605
box -3 -3 3 3
use M3_M2  M3_M2_5268
timestamp 1745462530
transform 1 0 180 0 1 3425
box -3 -3 3 3
use M3_M2  M3_M2_5269
timestamp 1745462530
transform 1 0 116 0 1 3425
box -3 -3 3 3
use M3_M2  M3_M2_5270
timestamp 1745462530
transform 1 0 276 0 1 3635
box -3 -3 3 3
use M3_M2  M3_M2_5271
timestamp 1745462530
transform 1 0 212 0 1 3645
box -3 -3 3 3
use M3_M2  M3_M2_5272
timestamp 1745462530
transform 1 0 428 0 1 3585
box -3 -3 3 3
use M3_M2  M3_M2_5273
timestamp 1745462530
transform 1 0 348 0 1 3585
box -3 -3 3 3
use M3_M2  M3_M2_5274
timestamp 1745462530
transform 1 0 204 0 1 3405
box -3 -3 3 3
use M3_M2  M3_M2_5275
timestamp 1745462530
transform 1 0 140 0 1 3405
box -3 -3 3 3
use M3_M2  M3_M2_5276
timestamp 1745462530
transform 1 0 268 0 1 3345
box -3 -3 3 3
use M3_M2  M3_M2_5277
timestamp 1745462530
transform 1 0 196 0 1 3345
box -3 -3 3 3
use M3_M2  M3_M2_5278
timestamp 1745462530
transform 1 0 2972 0 1 2685
box -3 -3 3 3
use M3_M2  M3_M2_5279
timestamp 1745462530
transform 1 0 2924 0 1 2685
box -3 -3 3 3
use M3_M2  M3_M2_5280
timestamp 1745462530
transform 1 0 2756 0 1 2325
box -3 -3 3 3
use M3_M2  M3_M2_5281
timestamp 1745462530
transform 1 0 2716 0 1 2325
box -3 -3 3 3
use M3_M2  M3_M2_5282
timestamp 1745462530
transform 1 0 3140 0 1 2455
box -3 -3 3 3
use M3_M2  M3_M2_5283
timestamp 1745462530
transform 1 0 3076 0 1 2385
box -3 -3 3 3
use M3_M2  M3_M2_5284
timestamp 1745462530
transform 1 0 3028 0 1 2455
box -3 -3 3 3
use M3_M2  M3_M2_5285
timestamp 1745462530
transform 1 0 3028 0 1 2385
box -3 -3 3 3
use M3_M2  M3_M2_5286
timestamp 1745462530
transform 1 0 2876 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_5287
timestamp 1745462530
transform 1 0 2820 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_5288
timestamp 1745462530
transform 1 0 3044 0 1 2545
box -3 -3 3 3
use M3_M2  M3_M2_5289
timestamp 1745462530
transform 1 0 2916 0 1 2545
box -3 -3 3 3
use M3_M2  M3_M2_5290
timestamp 1745462530
transform 1 0 4148 0 1 2835
box -3 -3 3 3
use M3_M2  M3_M2_5291
timestamp 1745462530
transform 1 0 4076 0 1 2545
box -3 -3 3 3
use M3_M2  M3_M2_5292
timestamp 1745462530
transform 1 0 4068 0 1 2835
box -3 -3 3 3
use M3_M2  M3_M2_5293
timestamp 1745462530
transform 1 0 4044 0 1 2545
box -3 -3 3 3
use M3_M2  M3_M2_5294
timestamp 1745462530
transform 1 0 4220 0 1 2635
box -3 -3 3 3
use M3_M2  M3_M2_5295
timestamp 1745462530
transform 1 0 4204 0 1 2895
box -3 -3 3 3
use M3_M2  M3_M2_5296
timestamp 1745462530
transform 1 0 4100 0 1 2895
box -3 -3 3 3
use M3_M2  M3_M2_5297
timestamp 1745462530
transform 1 0 4052 0 1 2625
box -3 -3 3 3
use M3_M2  M3_M2_5298
timestamp 1745462530
transform 1 0 3900 0 1 3075
box -3 -3 3 3
use M3_M2  M3_M2_5299
timestamp 1745462530
transform 1 0 3820 0 1 3075
box -3 -3 3 3
use M3_M2  M3_M2_5300
timestamp 1745462530
transform 1 0 3820 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_5301
timestamp 1745462530
transform 1 0 3700 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_5302
timestamp 1745462530
transform 1 0 3316 0 1 2805
box -3 -3 3 3
use M3_M2  M3_M2_5303
timestamp 1745462530
transform 1 0 3292 0 1 2845
box -3 -3 3 3
use M3_M2  M3_M2_5304
timestamp 1745462530
transform 1 0 3292 0 1 2805
box -3 -3 3 3
use M3_M2  M3_M2_5305
timestamp 1745462530
transform 1 0 2948 0 1 2845
box -3 -3 3 3
use M3_M2  M3_M2_5306
timestamp 1745462530
transform 1 0 3532 0 1 2555
box -3 -3 3 3
use M3_M2  M3_M2_5307
timestamp 1745462530
transform 1 0 3508 0 1 2555
box -3 -3 3 3
use M3_M2  M3_M2_5308
timestamp 1745462530
transform 1 0 3468 0 1 2555
box -3 -3 3 3
use M3_M2  M3_M2_5309
timestamp 1745462530
transform 1 0 4372 0 1 2365
box -3 -3 3 3
use M3_M2  M3_M2_5310
timestamp 1745462530
transform 1 0 4260 0 1 2365
box -3 -3 3 3
use M3_M2  M3_M2_5311
timestamp 1745462530
transform 1 0 4100 0 1 2365
box -3 -3 3 3
use M3_M2  M3_M2_5312
timestamp 1745462530
transform 1 0 4236 0 1 2175
box -3 -3 3 3
use M3_M2  M3_M2_5313
timestamp 1745462530
transform 1 0 4132 0 1 2175
box -3 -3 3 3
use M3_M2  M3_M2_5314
timestamp 1745462530
transform 1 0 4092 0 1 2175
box -3 -3 3 3
use M3_M2  M3_M2_5315
timestamp 1745462530
transform 1 0 4060 0 1 2315
box -3 -3 3 3
use M3_M2  M3_M2_5316
timestamp 1745462530
transform 1 0 3892 0 1 2315
box -3 -3 3 3
use M3_M2  M3_M2_5317
timestamp 1745462530
transform 1 0 3804 0 1 2315
box -3 -3 3 3
use M3_M2  M3_M2_5318
timestamp 1745462530
transform 1 0 3500 0 1 2385
box -3 -3 3 3
use M3_M2  M3_M2_5319
timestamp 1745462530
transform 1 0 3316 0 1 2385
box -3 -3 3 3
use M3_M2  M3_M2_5320
timestamp 1745462530
transform 1 0 3748 0 1 2245
box -3 -3 3 3
use M3_M2  M3_M2_5321
timestamp 1745462530
transform 1 0 3540 0 1 2245
box -3 -3 3 3
use M3_M2  M3_M2_5322
timestamp 1745462530
transform 1 0 4372 0 1 2565
box -3 -3 3 3
use M3_M2  M3_M2_5323
timestamp 1745462530
transform 1 0 4244 0 1 2565
box -3 -3 3 3
use M3_M2  M3_M2_5324
timestamp 1745462530
transform 1 0 4116 0 1 2565
box -3 -3 3 3
use M3_M2  M3_M2_5325
timestamp 1745462530
transform 1 0 3356 0 1 2545
box -3 -3 3 3
use M3_M2  M3_M2_5326
timestamp 1745462530
transform 1 0 3252 0 1 2545
box -3 -3 3 3
use M3_M2  M3_M2_5327
timestamp 1745462530
transform 1 0 3212 0 1 2545
box -3 -3 3 3
use M3_M2  M3_M2_5328
timestamp 1745462530
transform 1 0 4356 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_5329
timestamp 1745462530
transform 1 0 4188 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_5330
timestamp 1745462530
transform 1 0 4076 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_5331
timestamp 1745462530
transform 1 0 3972 0 1 2555
box -3 -3 3 3
use M3_M2  M3_M2_5332
timestamp 1745462530
transform 1 0 3796 0 1 2555
box -3 -3 3 3
use M3_M2  M3_M2_5333
timestamp 1745462530
transform 1 0 3764 0 1 2555
box -3 -3 3 3
use M3_M2  M3_M2_5334
timestamp 1745462530
transform 1 0 3460 0 1 2535
box -3 -3 3 3
use M3_M2  M3_M2_5335
timestamp 1745462530
transform 1 0 3436 0 1 2435
box -3 -3 3 3
use M3_M2  M3_M2_5336
timestamp 1745462530
transform 1 0 3412 0 1 2535
box -3 -3 3 3
use M3_M2  M3_M2_5337
timestamp 1745462530
transform 1 0 3412 0 1 2435
box -3 -3 3 3
use M3_M2  M3_M2_5338
timestamp 1745462530
transform 1 0 3796 0 1 2385
box -3 -3 3 3
use M3_M2  M3_M2_5339
timestamp 1745462530
transform 1 0 3612 0 1 2385
box -3 -3 3 3
use M3_M2  M3_M2_5340
timestamp 1745462530
transform 1 0 4332 0 1 2985
box -3 -3 3 3
use M3_M2  M3_M2_5341
timestamp 1745462530
transform 1 0 4324 0 1 2765
box -3 -3 3 3
use M3_M2  M3_M2_5342
timestamp 1745462530
transform 1 0 4308 0 1 2355
box -3 -3 3 3
use M3_M2  M3_M2_5343
timestamp 1745462530
transform 1 0 4204 0 1 2985
box -3 -3 3 3
use M3_M2  M3_M2_5344
timestamp 1745462530
transform 1 0 4148 0 1 2355
box -3 -3 3 3
use M3_M2  M3_M2_5345
timestamp 1745462530
transform 1 0 4076 0 1 2765
box -3 -3 3 3
use M3_M2  M3_M2_5346
timestamp 1745462530
transform 1 0 3220 0 1 2605
box -3 -3 3 3
use M3_M2  M3_M2_5347
timestamp 1745462530
transform 1 0 3188 0 1 2695
box -3 -3 3 3
use M3_M2  M3_M2_5348
timestamp 1745462530
transform 1 0 3188 0 1 2605
box -3 -3 3 3
use M3_M2  M3_M2_5349
timestamp 1745462530
transform 1 0 3164 0 1 2985
box -3 -3 3 3
use M3_M2  M3_M2_5350
timestamp 1745462530
transform 1 0 3036 0 1 2985
box -3 -3 3 3
use M3_M2  M3_M2_5351
timestamp 1745462530
transform 1 0 3036 0 1 2695
box -3 -3 3 3
use M3_M2  M3_M2_5352
timestamp 1745462530
transform 1 0 4372 0 1 2885
box -3 -3 3 3
use M3_M2  M3_M2_5353
timestamp 1745462530
transform 1 0 4268 0 1 2885
box -3 -3 3 3
use M3_M2  M3_M2_5354
timestamp 1745462530
transform 1 0 4228 0 1 2885
box -3 -3 3 3
use M3_M2  M3_M2_5355
timestamp 1745462530
transform 1 0 4228 0 1 2705
box -3 -3 3 3
use M3_M2  M3_M2_5356
timestamp 1745462530
transform 1 0 4124 0 1 2705
box -3 -3 3 3
use M3_M2  M3_M2_5357
timestamp 1745462530
transform 1 0 4076 0 1 2885
box -3 -3 3 3
use M3_M2  M3_M2_5358
timestamp 1745462530
transform 1 0 3876 0 1 2865
box -3 -3 3 3
use M3_M2  M3_M2_5359
timestamp 1745462530
transform 1 0 3844 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_5360
timestamp 1745462530
transform 1 0 3820 0 1 2865
box -3 -3 3 3
use M3_M2  M3_M2_5361
timestamp 1745462530
transform 1 0 3780 0 1 2535
box -3 -3 3 3
use M3_M2  M3_M2_5362
timestamp 1745462530
transform 1 0 3780 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_5363
timestamp 1745462530
transform 1 0 3764 0 1 2865
box -3 -3 3 3
use M3_M2  M3_M2_5364
timestamp 1745462530
transform 1 0 3732 0 1 2865
box -3 -3 3 3
use M3_M2  M3_M2_5365
timestamp 1745462530
transform 1 0 3732 0 1 2535
box -3 -3 3 3
use M3_M2  M3_M2_5366
timestamp 1745462530
transform 1 0 3444 0 1 2945
box -3 -3 3 3
use M3_M2  M3_M2_5367
timestamp 1745462530
transform 1 0 3348 0 1 2945
box -3 -3 3 3
use M3_M2  M3_M2_5368
timestamp 1745462530
transform 1 0 3324 0 1 2945
box -3 -3 3 3
use M3_M2  M3_M2_5369
timestamp 1745462530
transform 1 0 3684 0 1 2905
box -3 -3 3 3
use M3_M2  M3_M2_5370
timestamp 1745462530
transform 1 0 3596 0 1 2905
box -3 -3 3 3
use M3_M2  M3_M2_5371
timestamp 1745462530
transform 1 0 4268 0 1 2775
box -3 -3 3 3
use M3_M2  M3_M2_5372
timestamp 1745462530
transform 1 0 4084 0 1 2775
box -3 -3 3 3
use M3_M2  M3_M2_5373
timestamp 1745462530
transform 1 0 3148 0 1 2805
box -3 -3 3 3
use M3_M2  M3_M2_5374
timestamp 1745462530
transform 1 0 3004 0 1 2805
box -3 -3 3 3
use M3_M2  M3_M2_5375
timestamp 1745462530
transform 1 0 4372 0 1 2785
box -3 -3 3 3
use M3_M2  M3_M2_5376
timestamp 1745462530
transform 1 0 4116 0 1 2785
box -3 -3 3 3
use M3_M2  M3_M2_5377
timestamp 1745462530
transform 1 0 4028 0 1 2785
box -3 -3 3 3
use M3_M2  M3_M2_5378
timestamp 1745462530
transform 1 0 3988 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_5379
timestamp 1745462530
transform 1 0 3820 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_5380
timestamp 1745462530
transform 1 0 3788 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_5381
timestamp 1745462530
transform 1 0 3436 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_5382
timestamp 1745462530
transform 1 0 3356 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_5383
timestamp 1745462530
transform 1 0 3316 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_5384
timestamp 1745462530
transform 1 0 3772 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_5385
timestamp 1745462530
transform 1 0 3580 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_5386
timestamp 1745462530
transform 1 0 4076 0 1 3005
box -3 -3 3 3
use M3_M2  M3_M2_5387
timestamp 1745462530
transform 1 0 3964 0 1 3005
box -3 -3 3 3
use M3_M2  M3_M2_5388
timestamp 1745462530
transform 1 0 3124 0 1 2605
box -3 -3 3 3
use M3_M2  M3_M2_5389
timestamp 1745462530
transform 1 0 3068 0 1 2605
box -3 -3 3 3
use M3_M2  M3_M2_5390
timestamp 1745462530
transform 1 0 2988 0 1 2605
box -3 -3 3 3
use M3_M2  M3_M2_5391
timestamp 1745462530
transform 1 0 4044 0 1 2935
box -3 -3 3 3
use M3_M2  M3_M2_5392
timestamp 1745462530
transform 1 0 4012 0 1 2575
box -3 -3 3 3
use M3_M2  M3_M2_5393
timestamp 1745462530
transform 1 0 4004 0 1 2935
box -3 -3 3 3
use M3_M2  M3_M2_5394
timestamp 1745462530
transform 1 0 3988 0 1 2575
box -3 -3 3 3
use M3_M2  M3_M2_5395
timestamp 1745462530
transform 1 0 3940 0 1 2935
box -3 -3 3 3
use M3_M2  M3_M2_5396
timestamp 1745462530
transform 1 0 3772 0 1 2695
box -3 -3 3 3
use M3_M2  M3_M2_5397
timestamp 1745462530
transform 1 0 3772 0 1 2565
box -3 -3 3 3
use M3_M2  M3_M2_5398
timestamp 1745462530
transform 1 0 3732 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_5399
timestamp 1745462530
transform 1 0 3724 0 1 2925
box -3 -3 3 3
use M3_M2  M3_M2_5400
timestamp 1745462530
transform 1 0 3724 0 1 2695
box -3 -3 3 3
use M3_M2  M3_M2_5401
timestamp 1745462530
transform 1 0 3692 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_5402
timestamp 1745462530
transform 1 0 3684 0 1 2935
box -3 -3 3 3
use M3_M2  M3_M2_5403
timestamp 1745462530
transform 1 0 3652 0 1 2565
box -3 -3 3 3
use M3_M2  M3_M2_5404
timestamp 1745462530
transform 1 0 3404 0 1 2685
box -3 -3 3 3
use M3_M2  M3_M2_5405
timestamp 1745462530
transform 1 0 3332 0 1 2925
box -3 -3 3 3
use M3_M2  M3_M2_5406
timestamp 1745462530
transform 1 0 3308 0 1 2685
box -3 -3 3 3
use M3_M2  M3_M2_5407
timestamp 1745462530
transform 1 0 3268 0 1 2925
box -3 -3 3 3
use M3_M2  M3_M2_5408
timestamp 1745462530
transform 1 0 3268 0 1 2685
box -3 -3 3 3
use M3_M2  M3_M2_5409
timestamp 1745462530
transform 1 0 3604 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_5410
timestamp 1745462530
transform 1 0 3500 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_5411
timestamp 1745462530
transform 1 0 4340 0 1 2715
box -3 -3 3 3
use M3_M2  M3_M2_5412
timestamp 1745462530
transform 1 0 4156 0 1 2725
box -3 -3 3 3
use M3_M2  M3_M2_5413
timestamp 1745462530
transform 1 0 3932 0 1 2735
box -3 -3 3 3
use M3_M2  M3_M2_5414
timestamp 1745462530
transform 1 0 3252 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_5415
timestamp 1745462530
transform 1 0 3172 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_5416
timestamp 1745462530
transform 1 0 3092 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_5417
timestamp 1745462530
transform 1 0 4340 0 1 2625
box -3 -3 3 3
use M3_M2  M3_M2_5418
timestamp 1745462530
transform 1 0 4172 0 1 2625
box -3 -3 3 3
use M3_M2  M3_M2_5419
timestamp 1745462530
transform 1 0 4172 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_5420
timestamp 1745462530
transform 1 0 3980 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_5421
timestamp 1745462530
transform 1 0 3956 0 1 2695
box -3 -3 3 3
use M3_M2  M3_M2_5422
timestamp 1745462530
transform 1 0 3820 0 1 2695
box -3 -3 3 3
use M3_M2  M3_M2_5423
timestamp 1745462530
transform 1 0 3812 0 1 2725
box -3 -3 3 3
use M3_M2  M3_M2_5424
timestamp 1745462530
transform 1 0 3740 0 1 2725
box -3 -3 3 3
use M3_M2  M3_M2_5425
timestamp 1745462530
transform 1 0 3540 0 1 2805
box -3 -3 3 3
use M3_M2  M3_M2_5426
timestamp 1745462530
transform 1 0 3492 0 1 2805
box -3 -3 3 3
use M3_M2  M3_M2_5427
timestamp 1745462530
transform 1 0 3484 0 1 2695
box -3 -3 3 3
use M3_M2  M3_M2_5428
timestamp 1745462530
transform 1 0 3372 0 1 2695
box -3 -3 3 3
use M3_M2  M3_M2_5429
timestamp 1745462530
transform 1 0 3716 0 1 2725
box -3 -3 3 3
use M3_M2  M3_M2_5430
timestamp 1745462530
transform 1 0 3628 0 1 2725
box -3 -3 3 3
use M3_M2  M3_M2_5431
timestamp 1745462530
transform 1 0 3572 0 1 2725
box -3 -3 3 3
use M3_M2  M3_M2_5432
timestamp 1745462530
transform 1 0 3092 0 1 2135
box -3 -3 3 3
use M3_M2  M3_M2_5433
timestamp 1745462530
transform 1 0 3020 0 1 2135
box -3 -3 3 3
use M3_M2  M3_M2_5434
timestamp 1745462530
transform 1 0 2980 0 1 2135
box -3 -3 3 3
use M3_M2  M3_M2_5435
timestamp 1745462530
transform 1 0 2948 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_5436
timestamp 1745462530
transform 1 0 2900 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_5437
timestamp 1745462530
transform 1 0 2900 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_5438
timestamp 1745462530
transform 1 0 2820 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_5439
timestamp 1745462530
transform 1 0 2884 0 1 1695
box -3 -3 3 3
use M3_M2  M3_M2_5440
timestamp 1745462530
transform 1 0 2716 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_5441
timestamp 1745462530
transform 1 0 2676 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_5442
timestamp 1745462530
transform 1 0 2676 0 1 1695
box -3 -3 3 3
use M3_M2  M3_M2_5443
timestamp 1745462530
transform 1 0 2636 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_5444
timestamp 1745462530
transform 1 0 2604 0 1 1695
box -3 -3 3 3
use M3_M2  M3_M2_5445
timestamp 1745462530
transform 1 0 3012 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_5446
timestamp 1745462530
transform 1 0 2636 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_5447
timestamp 1745462530
transform 1 0 2988 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_5448
timestamp 1745462530
transform 1 0 2572 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_5449
timestamp 1745462530
transform 1 0 3028 0 1 2055
box -3 -3 3 3
use M3_M2  M3_M2_5450
timestamp 1745462530
transform 1 0 2716 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_5451
timestamp 1745462530
transform 1 0 2716 0 1 2055
box -3 -3 3 3
use M3_M2  M3_M2_5452
timestamp 1745462530
transform 1 0 2684 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_5453
timestamp 1745462530
transform 1 0 3932 0 1 2135
box -3 -3 3 3
use M3_M2  M3_M2_5454
timestamp 1745462530
transform 1 0 3276 0 1 2175
box -3 -3 3 3
use M3_M2  M3_M2_5455
timestamp 1745462530
transform 1 0 3276 0 1 2135
box -3 -3 3 3
use M3_M2  M3_M2_5456
timestamp 1745462530
transform 1 0 3172 0 1 2165
box -3 -3 3 3
use M3_M2  M3_M2_5457
timestamp 1745462530
transform 1 0 2988 0 1 2165
box -3 -3 3 3
use M3_M2  M3_M2_5458
timestamp 1745462530
transform 1 0 3148 0 1 1665
box -3 -3 3 3
use M3_M2  M3_M2_5459
timestamp 1745462530
transform 1 0 2908 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_5460
timestamp 1745462530
transform 1 0 2908 0 1 1665
box -3 -3 3 3
use M3_M2  M3_M2_5461
timestamp 1745462530
transform 1 0 2868 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_5462
timestamp 1745462530
transform 1 0 3044 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_5463
timestamp 1745462530
transform 1 0 2932 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_5464
timestamp 1745462530
transform 1 0 2852 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_5465
timestamp 1745462530
transform 1 0 3284 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_5466
timestamp 1745462530
transform 1 0 3284 0 1 1465
box -3 -3 3 3
use M3_M2  M3_M2_5467
timestamp 1745462530
transform 1 0 3236 0 1 1465
box -3 -3 3 3
use M3_M2  M3_M2_5468
timestamp 1745462530
transform 1 0 3148 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_5469
timestamp 1745462530
transform 1 0 3028 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_5470
timestamp 1745462530
transform 1 0 3028 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_5471
timestamp 1745462530
transform 1 0 2980 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_5472
timestamp 1745462530
transform 1 0 3060 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_5473
timestamp 1745462530
transform 1 0 2908 0 1 2205
box -3 -3 3 3
use M3_M2  M3_M2_5474
timestamp 1745462530
transform 1 0 2908 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_5475
timestamp 1745462530
transform 1 0 2756 0 1 2205
box -3 -3 3 3
use M3_M2  M3_M2_5476
timestamp 1745462530
transform 1 0 3244 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_5477
timestamp 1745462530
transform 1 0 2988 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_5478
timestamp 1745462530
transform 1 0 2988 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_5479
timestamp 1745462530
transform 1 0 2900 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_5480
timestamp 1745462530
transform 1 0 4036 0 1 2235
box -3 -3 3 3
use M3_M2  M3_M2_5481
timestamp 1745462530
transform 1 0 4028 0 1 2125
box -3 -3 3 3
use M3_M2  M3_M2_5482
timestamp 1745462530
transform 1 0 3924 0 1 2045
box -3 -3 3 3
use M3_M2  M3_M2_5483
timestamp 1745462530
transform 1 0 3892 0 1 2235
box -3 -3 3 3
use M3_M2  M3_M2_5484
timestamp 1745462530
transform 1 0 3852 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_5485
timestamp 1745462530
transform 1 0 3852 0 1 2045
box -3 -3 3 3
use M3_M2  M3_M2_5486
timestamp 1745462530
transform 1 0 3340 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_5487
timestamp 1745462530
transform 1 0 3220 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_5488
timestamp 1745462530
transform 1 0 3116 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_5489
timestamp 1745462530
transform 1 0 3388 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_5490
timestamp 1745462530
transform 1 0 3388 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_5491
timestamp 1745462530
transform 1 0 3332 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_5492
timestamp 1745462530
transform 1 0 3220 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_5493
timestamp 1745462530
transform 1 0 4044 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_5494
timestamp 1745462530
transform 1 0 3916 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_5495
timestamp 1745462530
transform 1 0 3828 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_5496
timestamp 1745462530
transform 1 0 3708 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_5497
timestamp 1745462530
transform 1 0 3532 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_5498
timestamp 1745462530
transform 1 0 3468 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_5499
timestamp 1745462530
transform 1 0 3332 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_5500
timestamp 1745462530
transform 1 0 3324 0 1 2175
box -3 -3 3 3
use M3_M2  M3_M2_5501
timestamp 1745462530
transform 1 0 3300 0 1 2175
box -3 -3 3 3
use M3_M2  M3_M2_5502
timestamp 1745462530
transform 1 0 3724 0 1 2175
box -3 -3 3 3
use M3_M2  M3_M2_5503
timestamp 1745462530
transform 1 0 3588 0 1 2175
box -3 -3 3 3
use M3_M2  M3_M2_5504
timestamp 1745462530
transform 1 0 3588 0 1 2075
box -3 -3 3 3
use M3_M2  M3_M2_5505
timestamp 1745462530
transform 1 0 3532 0 1 2075
box -3 -3 3 3
use M3_M2  M3_M2_5506
timestamp 1745462530
transform 1 0 3356 0 1 2075
box -3 -3 3 3
use M3_M2  M3_M2_5507
timestamp 1745462530
transform 1 0 4276 0 1 2095
box -3 -3 3 3
use M3_M2  M3_M2_5508
timestamp 1745462530
transform 1 0 4180 0 1 2095
box -3 -3 3 3
use M3_M2  M3_M2_5509
timestamp 1745462530
transform 1 0 3996 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_5510
timestamp 1745462530
transform 1 0 3820 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_5511
timestamp 1745462530
transform 1 0 4292 0 1 1695
box -3 -3 3 3
use M3_M2  M3_M2_5512
timestamp 1745462530
transform 1 0 4132 0 1 1695
box -3 -3 3 3
use M3_M2  M3_M2_5513
timestamp 1745462530
transform 1 0 3300 0 1 1695
box -3 -3 3 3
use M3_M2  M3_M2_5514
timestamp 1745462530
transform 1 0 3292 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_5515
timestamp 1745462530
transform 1 0 3188 0 1 1695
box -3 -3 3 3
use M3_M2  M3_M2_5516
timestamp 1745462530
transform 1 0 3156 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_5517
timestamp 1745462530
transform 1 0 4356 0 1 1665
box -3 -3 3 3
use M3_M2  M3_M2_5518
timestamp 1745462530
transform 1 0 3316 0 1 1665
box -3 -3 3 3
use M3_M2  M3_M2_5519
timestamp 1745462530
transform 1 0 3308 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_5520
timestamp 1745462530
transform 1 0 3220 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_5521
timestamp 1745462530
transform 1 0 4068 0 1 1685
box -3 -3 3 3
use M3_M2  M3_M2_5522
timestamp 1745462530
transform 1 0 3916 0 1 1685
box -3 -3 3 3
use M3_M2  M3_M2_5523
timestamp 1745462530
transform 1 0 3916 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_5524
timestamp 1745462530
transform 1 0 3796 0 1 1685
box -3 -3 3 3
use M3_M2  M3_M2_5525
timestamp 1745462530
transform 1 0 3708 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_5526
timestamp 1745462530
transform 1 0 4180 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_5527
timestamp 1745462530
transform 1 0 4100 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_5528
timestamp 1745462530
transform 1 0 4100 0 1 2065
box -3 -3 3 3
use M3_M2  M3_M2_5529
timestamp 1745462530
transform 1 0 3444 0 1 2065
box -3 -3 3 3
use M3_M2  M3_M2_5530
timestamp 1745462530
transform 1 0 4372 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_5531
timestamp 1745462530
transform 1 0 4324 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_5532
timestamp 1745462530
transform 1 0 3540 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_5533
timestamp 1745462530
transform 1 0 3396 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_5534
timestamp 1745462530
transform 1 0 4084 0 1 2015
box -3 -3 3 3
use M3_M2  M3_M2_5535
timestamp 1745462530
transform 1 0 3996 0 1 2015
box -3 -3 3 3
use M3_M2  M3_M2_5536
timestamp 1745462530
transform 1 0 3900 0 1 2015
box -3 -3 3 3
use M3_M2  M3_M2_5537
timestamp 1745462530
transform 1 0 3540 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_5538
timestamp 1745462530
transform 1 0 3412 0 1 1575
box -3 -3 3 3
use M3_M2  M3_M2_5539
timestamp 1745462530
transform 1 0 3156 0 1 1575
box -3 -3 3 3
use M3_M2  M3_M2_5540
timestamp 1745462530
transform 1 0 3684 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_5541
timestamp 1745462530
transform 1 0 3604 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_5542
timestamp 1745462530
transform 1 0 3604 0 1 1485
box -3 -3 3 3
use M3_M2  M3_M2_5543
timestamp 1745462530
transform 1 0 3244 0 1 1495
box -3 -3 3 3
use M3_M2  M3_M2_5544
timestamp 1745462530
transform 1 0 3956 0 1 1575
box -3 -3 3 3
use M3_M2  M3_M2_5545
timestamp 1745462530
transform 1 0 3844 0 1 1575
box -3 -3 3 3
use M3_M2  M3_M2_5546
timestamp 1745462530
transform 1 0 3748 0 1 1575
box -3 -3 3 3
use M3_M2  M3_M2_5547
timestamp 1745462530
transform 1 0 3700 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_5548
timestamp 1745462530
transform 1 0 3636 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_5549
timestamp 1745462530
transform 1 0 3348 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_5550
timestamp 1745462530
transform 1 0 3796 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_5551
timestamp 1745462530
transform 1 0 3732 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_5552
timestamp 1745462530
transform 1 0 3708 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_5553
timestamp 1745462530
transform 1 0 3700 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_5554
timestamp 1745462530
transform 1 0 3428 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_5555
timestamp 1745462530
transform 1 0 4372 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_5556
timestamp 1745462530
transform 1 0 4260 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_5557
timestamp 1745462530
transform 1 0 4196 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_5558
timestamp 1745462530
transform 1 0 4028 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_5559
timestamp 1745462530
transform 1 0 4364 0 1 1525
box -3 -3 3 3
use M3_M2  M3_M2_5560
timestamp 1745462530
transform 1 0 4268 0 1 1525
box -3 -3 3 3
use M3_M2  M3_M2_5561
timestamp 1745462530
transform 1 0 4364 0 1 1405
box -3 -3 3 3
use M3_M2  M3_M2_5562
timestamp 1745462530
transform 1 0 4260 0 1 1405
box -3 -3 3 3
use M3_M2  M3_M2_5563
timestamp 1745462530
transform 1 0 4156 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_5564
timestamp 1745462530
transform 1 0 4092 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_5565
timestamp 1745462530
transform 1 0 4380 0 1 1895
box -3 -3 3 3
use M3_M2  M3_M2_5566
timestamp 1745462530
transform 1 0 4268 0 1 1895
box -3 -3 3 3
use M3_M2  M3_M2_5567
timestamp 1745462530
transform 1 0 4052 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_5568
timestamp 1745462530
transform 1 0 4052 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_5569
timestamp 1745462530
transform 1 0 3940 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_5570
timestamp 1745462530
transform 1 0 3916 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_5571
timestamp 1745462530
transform 1 0 3588 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_5572
timestamp 1745462530
transform 1 0 3468 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_5573
timestamp 1745462530
transform 1 0 3460 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_5574
timestamp 1745462530
transform 1 0 3084 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_5575
timestamp 1745462530
transform 1 0 3716 0 1 1375
box -3 -3 3 3
use M3_M2  M3_M2_5576
timestamp 1745462530
transform 1 0 3636 0 1 1375
box -3 -3 3 3
use M3_M2  M3_M2_5577
timestamp 1745462530
transform 1 0 3596 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_5578
timestamp 1745462530
transform 1 0 2988 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_5579
timestamp 1745462530
transform 1 0 3836 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_5580
timestamp 1745462530
transform 1 0 3172 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_5581
timestamp 1745462530
transform 1 0 3428 0 1 1815
box -3 -3 3 3
use M3_M2  M3_M2_5582
timestamp 1745462530
transform 1 0 3028 0 1 1815
box -3 -3 3 3
use M3_M2  M3_M2_5583
timestamp 1745462530
transform 1 0 3636 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_5584
timestamp 1745462530
transform 1 0 3196 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_5585
timestamp 1745462530
transform 1 0 4156 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_5586
timestamp 1745462530
transform 1 0 4044 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_5587
timestamp 1745462530
transform 1 0 4364 0 1 1335
box -3 -3 3 3
use M3_M2  M3_M2_5588
timestamp 1745462530
transform 1 0 4260 0 1 1335
box -3 -3 3 3
use M3_M2  M3_M2_5589
timestamp 1745462530
transform 1 0 4268 0 1 1285
box -3 -3 3 3
use M3_M2  M3_M2_5590
timestamp 1745462530
transform 1 0 4172 0 1 1285
box -3 -3 3 3
use M3_M2  M3_M2_5591
timestamp 1745462530
transform 1 0 4028 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_5592
timestamp 1745462530
transform 1 0 3932 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_5593
timestamp 1745462530
transform 1 0 4356 0 1 1815
box -3 -3 3 3
use M3_M2  M3_M2_5594
timestamp 1745462530
transform 1 0 4260 0 1 1815
box -3 -3 3 3
use M3_M2  M3_M2_5595
timestamp 1745462530
transform 1 0 4164 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_5596
timestamp 1745462530
transform 1 0 3844 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_5597
timestamp 1745462530
transform 1 0 3308 0 1 1215
box -3 -3 3 3
use M3_M2  M3_M2_5598
timestamp 1745462530
transform 1 0 3100 0 1 1215
box -3 -3 3 3
use M3_M2  M3_M2_5599
timestamp 1745462530
transform 1 0 4076 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_5600
timestamp 1745462530
transform 1 0 3964 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_5601
timestamp 1745462530
transform 1 0 3924 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_5602
timestamp 1745462530
transform 1 0 3788 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_5603
timestamp 1745462530
transform 1 0 3740 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_5604
timestamp 1745462530
transform 1 0 3700 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_5605
timestamp 1745462530
transform 1 0 3692 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_5606
timestamp 1745462530
transform 1 0 3668 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_5607
timestamp 1745462530
transform 1 0 3564 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_5608
timestamp 1745462530
transform 1 0 3420 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_5609
timestamp 1745462530
transform 1 0 3412 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_5610
timestamp 1745462530
transform 1 0 3340 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_5611
timestamp 1745462530
transform 1 0 3676 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_5612
timestamp 1745462530
transform 1 0 3572 0 1 1215
box -3 -3 3 3
use M3_M2  M3_M2_5613
timestamp 1745462530
transform 1 0 3540 0 1 1215
box -3 -3 3 3
use M3_M2  M3_M2_5614
timestamp 1745462530
transform 1 0 3540 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_5615
timestamp 1745462530
transform 1 0 4268 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_5616
timestamp 1745462530
transform 1 0 4092 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_5617
timestamp 1745462530
transform 1 0 3964 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_5618
timestamp 1745462530
transform 1 0 3812 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_5619
timestamp 1745462530
transform 1 0 3340 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_5620
timestamp 1745462530
transform 1 0 3340 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_5621
timestamp 1745462530
transform 1 0 3316 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_5622
timestamp 1745462530
transform 1 0 3308 0 1 1015
box -3 -3 3 3
use M3_M2  M3_M2_5623
timestamp 1745462530
transform 1 0 3276 0 1 1015
box -3 -3 3 3
use M3_M2  M3_M2_5624
timestamp 1745462530
transform 1 0 3172 0 1 865
box -3 -3 3 3
use M3_M2  M3_M2_5625
timestamp 1745462530
transform 1 0 4364 0 1 1135
box -3 -3 3 3
use M3_M2  M3_M2_5626
timestamp 1745462530
transform 1 0 4260 0 1 1135
box -3 -3 3 3
use M3_M2  M3_M2_5627
timestamp 1745462530
transform 1 0 4004 0 1 1135
box -3 -3 3 3
use M3_M2  M3_M2_5628
timestamp 1745462530
transform 1 0 3868 0 1 1135
box -3 -3 3 3
use M3_M2  M3_M2_5629
timestamp 1745462530
transform 1 0 3836 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_5630
timestamp 1745462530
transform 1 0 3748 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_5631
timestamp 1745462530
transform 1 0 3676 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_5632
timestamp 1745462530
transform 1 0 3516 0 1 1055
box -3 -3 3 3
use M3_M2  M3_M2_5633
timestamp 1745462530
transform 1 0 3500 0 1 1055
box -3 -3 3 3
use M3_M2  M3_M2_5634
timestamp 1745462530
transform 1 0 3340 0 1 1055
box -3 -3 3 3
use M3_M2  M3_M2_5635
timestamp 1745462530
transform 1 0 4188 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_5636
timestamp 1745462530
transform 1 0 4124 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_5637
timestamp 1745462530
transform 1 0 3612 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_5638
timestamp 1745462530
transform 1 0 4372 0 1 1035
box -3 -3 3 3
use M3_M2  M3_M2_5639
timestamp 1745462530
transform 1 0 4364 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_5640
timestamp 1745462530
transform 1 0 3980 0 1 1075
box -3 -3 3 3
use M3_M2  M3_M2_5641
timestamp 1745462530
transform 1 0 4068 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_5642
timestamp 1745462530
transform 1 0 3988 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_5643
timestamp 1745462530
transform 1 0 3356 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_5644
timestamp 1745462530
transform 1 0 3356 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_5645
timestamp 1745462530
transform 1 0 3188 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_5646
timestamp 1745462530
transform 1 0 4372 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_5647
timestamp 1745462530
transform 1 0 4180 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_5648
timestamp 1745462530
transform 1 0 4036 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_5649
timestamp 1745462530
transform 1 0 3980 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_5650
timestamp 1745462530
transform 1 0 4212 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_5651
timestamp 1745462530
transform 1 0 4092 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_5652
timestamp 1745462530
transform 1 0 3900 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_5653
timestamp 1745462530
transform 1 0 3900 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_5654
timestamp 1745462530
transform 1 0 3804 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_5655
timestamp 1745462530
transform 1 0 3916 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_5656
timestamp 1745462530
transform 1 0 3516 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_5657
timestamp 1745462530
transform 1 0 3364 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_5658
timestamp 1745462530
transform 1 0 4372 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_5659
timestamp 1745462530
transform 1 0 4188 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_5660
timestamp 1745462530
transform 1 0 3692 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_5661
timestamp 1745462530
transform 1 0 4244 0 1 335
box -3 -3 3 3
use M3_M2  M3_M2_5662
timestamp 1745462530
transform 1 0 4116 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_5663
timestamp 1745462530
transform 1 0 4116 0 1 335
box -3 -3 3 3
use M3_M2  M3_M2_5664
timestamp 1745462530
transform 1 0 3948 0 1 975
box -3 -3 3 3
use M3_M2  M3_M2_5665
timestamp 1745462530
transform 1 0 3940 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_5666
timestamp 1745462530
transform 1 0 3916 0 1 975
box -3 -3 3 3
use M3_M2  M3_M2_5667
timestamp 1745462530
transform 1 0 4284 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_5668
timestamp 1745462530
transform 1 0 4076 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_5669
timestamp 1745462530
transform 1 0 3324 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_5670
timestamp 1745462530
transform 1 0 3324 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_5671
timestamp 1745462530
transform 1 0 3276 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_5672
timestamp 1745462530
transform 1 0 4380 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_5673
timestamp 1745462530
transform 1 0 4036 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_5674
timestamp 1745462530
transform 1 0 3916 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_5675
timestamp 1745462530
transform 1 0 4372 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_5676
timestamp 1745462530
transform 1 0 4260 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_5677
timestamp 1745462530
transform 1 0 4260 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_5678
timestamp 1745462530
transform 1 0 3844 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_5679
timestamp 1745462530
transform 1 0 3748 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_5680
timestamp 1745462530
transform 1 0 4036 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_5681
timestamp 1745462530
transform 1 0 3492 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_5682
timestamp 1745462530
transform 1 0 3476 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_5683
timestamp 1745462530
transform 1 0 3380 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_5684
timestamp 1745462530
transform 1 0 4372 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_5685
timestamp 1745462530
transform 1 0 4228 0 1 725
box -3 -3 3 3
use M3_M2  M3_M2_5686
timestamp 1745462530
transform 1 0 3612 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_5687
timestamp 1745462530
transform 1 0 4116 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_5688
timestamp 1745462530
transform 1 0 4036 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_5689
timestamp 1745462530
transform 1 0 3428 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_5690
timestamp 1745462530
transform 1 0 3324 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_5691
timestamp 1745462530
transform 1 0 3244 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_5692
timestamp 1745462530
transform 1 0 3244 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_5693
timestamp 1745462530
transform 1 0 3228 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_5694
timestamp 1745462530
transform 1 0 4132 0 1 375
box -3 -3 3 3
use M3_M2  M3_M2_5695
timestamp 1745462530
transform 1 0 4068 0 1 375
box -3 -3 3 3
use M3_M2  M3_M2_5696
timestamp 1745462530
transform 1 0 3972 0 1 375
box -3 -3 3 3
use M3_M2  M3_M2_5697
timestamp 1745462530
transform 1 0 3924 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_5698
timestamp 1745462530
transform 1 0 3836 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_5699
timestamp 1745462530
transform 1 0 3548 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_5700
timestamp 1745462530
transform 1 0 3396 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_5701
timestamp 1745462530
transform 1 0 3708 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_5702
timestamp 1745462530
transform 1 0 3684 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_5703
timestamp 1745462530
transform 1 0 4220 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_5704
timestamp 1745462530
transform 1 0 4108 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_5705
timestamp 1745462530
transform 1 0 4196 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_5706
timestamp 1745462530
transform 1 0 4092 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_5707
timestamp 1745462530
transform 1 0 4356 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_5708
timestamp 1745462530
transform 1 0 4244 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_5709
timestamp 1745462530
transform 1 0 4372 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_5710
timestamp 1745462530
transform 1 0 4260 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_5711
timestamp 1745462530
transform 1 0 4084 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_5712
timestamp 1745462530
transform 1 0 3964 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_5713
timestamp 1745462530
transform 1 0 3764 0 1 155
box -3 -3 3 3
use M3_M2  M3_M2_5714
timestamp 1745462530
transform 1 0 3708 0 1 155
box -3 -3 3 3
use M3_M2  M3_M2_5715
timestamp 1745462530
transform 1 0 4020 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_5716
timestamp 1745462530
transform 1 0 4020 0 1 575
box -3 -3 3 3
use M3_M2  M3_M2_5717
timestamp 1745462530
transform 1 0 3972 0 1 575
box -3 -3 3 3
use M3_M2  M3_M2_5718
timestamp 1745462530
transform 1 0 3924 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_5719
timestamp 1745462530
transform 1 0 3196 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_5720
timestamp 1745462530
transform 1 0 3084 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_5721
timestamp 1745462530
transform 1 0 3996 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_5722
timestamp 1745462530
transform 1 0 3956 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_5723
timestamp 1745462530
transform 1 0 3956 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_5724
timestamp 1745462530
transform 1 0 3876 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_5725
timestamp 1745462530
transform 1 0 3828 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_5726
timestamp 1745462530
transform 1 0 3772 0 1 535
box -3 -3 3 3
use M3_M2  M3_M2_5727
timestamp 1745462530
transform 1 0 3660 0 1 535
box -3 -3 3 3
use M3_M2  M3_M2_5728
timestamp 1745462530
transform 1 0 3492 0 1 495
box -3 -3 3 3
use M3_M2  M3_M2_5729
timestamp 1745462530
transform 1 0 3412 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_5730
timestamp 1745462530
transform 1 0 3412 0 1 495
box -3 -3 3 3
use M3_M2  M3_M2_5731
timestamp 1745462530
transform 1 0 3324 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_5732
timestamp 1745462530
transform 1 0 3300 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_5733
timestamp 1745462530
transform 1 0 3276 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_5734
timestamp 1745462530
transform 1 0 3644 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_5735
timestamp 1745462530
transform 1 0 3604 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_5736
timestamp 1745462530
transform 1 0 3564 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_5737
timestamp 1745462530
transform 1 0 3084 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_5738
timestamp 1745462530
transform 1 0 2972 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_5739
timestamp 1745462530
transform 1 0 2860 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_5740
timestamp 1745462530
transform 1 0 3044 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_5741
timestamp 1745462530
transform 1 0 3044 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_5742
timestamp 1745462530
transform 1 0 3028 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_5743
timestamp 1745462530
transform 1 0 3004 0 1 1435
box -3 -3 3 3
use M3_M2  M3_M2_5744
timestamp 1745462530
transform 1 0 3004 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_5745
timestamp 1745462530
transform 1 0 2892 0 1 1435
box -3 -3 3 3
use M3_M2  M3_M2_5746
timestamp 1745462530
transform 1 0 2468 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_5747
timestamp 1745462530
transform 1 0 2324 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_5748
timestamp 1745462530
transform 1 0 2652 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_5749
timestamp 1745462530
transform 1 0 2548 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_5750
timestamp 1745462530
transform 1 0 2540 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_5751
timestamp 1745462530
transform 1 0 2516 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_5752
timestamp 1745462530
transform 1 0 2532 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_5753
timestamp 1745462530
transform 1 0 2452 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_5754
timestamp 1745462530
transform 1 0 2812 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_5755
timestamp 1745462530
transform 1 0 2756 0 1 1435
box -3 -3 3 3
use M3_M2  M3_M2_5756
timestamp 1745462530
transform 1 0 2708 0 1 1435
box -3 -3 3 3
use M3_M2  M3_M2_5757
timestamp 1745462530
transform 1 0 2708 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_5758
timestamp 1745462530
transform 1 0 3172 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_5759
timestamp 1745462530
transform 1 0 3084 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_5760
timestamp 1745462530
transform 1 0 2908 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_5761
timestamp 1745462530
transform 1 0 3100 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_5762
timestamp 1745462530
transform 1 0 2972 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_5763
timestamp 1745462530
transform 1 0 2868 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_5764
timestamp 1745462530
transform 1 0 2428 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_5765
timestamp 1745462530
transform 1 0 2268 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_5766
timestamp 1745462530
transform 1 0 2268 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_5767
timestamp 1745462530
transform 1 0 2244 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_5768
timestamp 1745462530
transform 1 0 2668 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_5769
timestamp 1745462530
transform 1 0 2564 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_5770
timestamp 1745462530
transform 1 0 2524 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_5771
timestamp 1745462530
transform 1 0 2484 0 1 1205
box -3 -3 3 3
use M3_M2  M3_M2_5772
timestamp 1745462530
transform 1 0 2412 0 1 1205
box -3 -3 3 3
use M3_M2  M3_M2_5773
timestamp 1745462530
transform 1 0 2788 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_5774
timestamp 1745462530
transform 1 0 2716 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_5775
timestamp 1745462530
transform 1 0 3100 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_5776
timestamp 1745462530
transform 1 0 3036 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_5777
timestamp 1745462530
transform 1 0 3012 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_5778
timestamp 1745462530
transform 1 0 2956 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_5779
timestamp 1745462530
transform 1 0 3076 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_5780
timestamp 1745462530
transform 1 0 2988 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_5781
timestamp 1745462530
transform 1 0 2988 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_5782
timestamp 1745462530
transform 1 0 2892 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_5783
timestamp 1745462530
transform 1 0 2500 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_5784
timestamp 1745462530
transform 1 0 2404 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_5785
timestamp 1745462530
transform 1 0 2316 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_5786
timestamp 1745462530
transform 1 0 2276 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_5787
timestamp 1745462530
transform 1 0 2532 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_5788
timestamp 1745462530
transform 1 0 2396 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_5789
timestamp 1745462530
transform 1 0 2308 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_5790
timestamp 1745462530
transform 1 0 2244 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_5791
timestamp 1745462530
transform 1 0 2692 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_5792
timestamp 1745462530
transform 1 0 2692 0 1 865
box -3 -3 3 3
use M3_M2  M3_M2_5793
timestamp 1745462530
transform 1 0 2668 0 1 865
box -3 -3 3 3
use M3_M2  M3_M2_5794
timestamp 1745462530
transform 1 0 2516 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_5795
timestamp 1745462530
transform 1 0 2428 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_5796
timestamp 1745462530
transform 1 0 2868 0 1 865
box -3 -3 3 3
use M3_M2  M3_M2_5797
timestamp 1745462530
transform 1 0 2764 0 1 865
box -3 -3 3 3
use M3_M2  M3_M2_5798
timestamp 1745462530
transform 1 0 3204 0 1 165
box -3 -3 3 3
use M3_M2  M3_M2_5799
timestamp 1745462530
transform 1 0 3156 0 1 165
box -3 -3 3 3
use M3_M2  M3_M2_5800
timestamp 1745462530
transform 1 0 3148 0 1 675
box -3 -3 3 3
use M3_M2  M3_M2_5801
timestamp 1745462530
transform 1 0 3116 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_5802
timestamp 1745462530
transform 1 0 3100 0 1 845
box -3 -3 3 3
use M3_M2  M3_M2_5803
timestamp 1745462530
transform 1 0 3100 0 1 675
box -3 -3 3 3
use M3_M2  M3_M2_5804
timestamp 1745462530
transform 1 0 3076 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_5805
timestamp 1745462530
transform 1 0 3060 0 1 845
box -3 -3 3 3
use M3_M2  M3_M2_5806
timestamp 1745462530
transform 1 0 3116 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_5807
timestamp 1745462530
transform 1 0 2996 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_5808
timestamp 1745462530
transform 1 0 2468 0 1 875
box -3 -3 3 3
use M3_M2  M3_M2_5809
timestamp 1745462530
transform 1 0 2444 0 1 875
box -3 -3 3 3
use M3_M2  M3_M2_5810
timestamp 1745462530
transform 1 0 2236 0 1 865
box -3 -3 3 3
use M3_M2  M3_M2_5811
timestamp 1745462530
transform 1 0 2676 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_5812
timestamp 1745462530
transform 1 0 2628 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_5813
timestamp 1745462530
transform 1 0 2604 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_5814
timestamp 1745462530
transform 1 0 2580 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_5815
timestamp 1745462530
transform 1 0 2452 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_5816
timestamp 1745462530
transform 1 0 3092 0 1 285
box -3 -3 3 3
use M3_M2  M3_M2_5817
timestamp 1745462530
transform 1 0 2980 0 1 285
box -3 -3 3 3
use M3_M2  M3_M2_5818
timestamp 1745462530
transform 1 0 2828 0 1 845
box -3 -3 3 3
use M3_M2  M3_M2_5819
timestamp 1745462530
transform 1 0 2820 0 1 285
box -3 -3 3 3
use M3_M2  M3_M2_5820
timestamp 1745462530
transform 1 0 2780 0 1 845
box -3 -3 3 3
use M3_M2  M3_M2_5821
timestamp 1745462530
transform 1 0 3084 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_5822
timestamp 1745462530
transform 1 0 3052 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_5823
timestamp 1745462530
transform 1 0 2972 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_5824
timestamp 1745462530
transform 1 0 3156 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_5825
timestamp 1745462530
transform 1 0 3044 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_5826
timestamp 1745462530
transform 1 0 2380 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_5827
timestamp 1745462530
transform 1 0 2196 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_5828
timestamp 1745462530
transform 1 0 2436 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_5829
timestamp 1745462530
transform 1 0 2412 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_5830
timestamp 1745462530
transform 1 0 2356 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_5831
timestamp 1745462530
transform 1 0 2460 0 1 475
box -3 -3 3 3
use M3_M2  M3_M2_5832
timestamp 1745462530
transform 1 0 2340 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_5833
timestamp 1745462530
transform 1 0 2212 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_5834
timestamp 1745462530
transform 1 0 2844 0 1 655
box -3 -3 3 3
use M3_M2  M3_M2_5835
timestamp 1745462530
transform 1 0 2804 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_5836
timestamp 1745462530
transform 1 0 2748 0 1 655
box -3 -3 3 3
use M3_M2  M3_M2_5837
timestamp 1745462530
transform 1 0 2748 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_5838
timestamp 1745462530
transform 1 0 3196 0 1 645
box -3 -3 3 3
use M3_M2  M3_M2_5839
timestamp 1745462530
transform 1 0 3132 0 1 645
box -3 -3 3 3
use M3_M2  M3_M2_5840
timestamp 1745462530
transform 1 0 3068 0 1 645
box -3 -3 3 3
use M3_M2  M3_M2_5841
timestamp 1745462530
transform 1 0 3228 0 1 685
box -3 -3 3 3
use M3_M2  M3_M2_5842
timestamp 1745462530
transform 1 0 3116 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_5843
timestamp 1745462530
transform 1 0 3116 0 1 685
box -3 -3 3 3
use M3_M2  M3_M2_5844
timestamp 1745462530
transform 1 0 3108 0 1 1005
box -3 -3 3 3
use M3_M2  M3_M2_5845
timestamp 1745462530
transform 1 0 3092 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_5846
timestamp 1745462530
transform 1 0 3076 0 1 1005
box -3 -3 3 3
use M3_M2  M3_M2_5847
timestamp 1745462530
transform 1 0 2196 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_5848
timestamp 1745462530
transform 1 0 2172 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_5849
timestamp 1745462530
transform 1 0 2484 0 1 775
box -3 -3 3 3
use M3_M2  M3_M2_5850
timestamp 1745462530
transform 1 0 2428 0 1 775
box -3 -3 3 3
use M3_M2  M3_M2_5851
timestamp 1745462530
transform 1 0 2372 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_5852
timestamp 1745462530
transform 1 0 2244 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_5853
timestamp 1745462530
transform 1 0 2244 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_5854
timestamp 1745462530
transform 1 0 2180 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_5855
timestamp 1745462530
transform 1 0 2868 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_5856
timestamp 1745462530
transform 1 0 2860 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_5857
timestamp 1745462530
transform 1 0 2788 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_5858
timestamp 1745462530
transform 1 0 2740 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_5859
timestamp 1745462530
transform 1 0 2932 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_5860
timestamp 1745462530
transform 1 0 2884 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_5861
timestamp 1745462530
transform 1 0 2772 0 1 165
box -3 -3 3 3
use M3_M2  M3_M2_5862
timestamp 1745462530
transform 1 0 2700 0 1 165
box -3 -3 3 3
use M3_M2  M3_M2_5863
timestamp 1745462530
transform 1 0 1788 0 1 1295
box -3 -3 3 3
use M3_M2  M3_M2_5864
timestamp 1745462530
transform 1 0 1748 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_5865
timestamp 1745462530
transform 1 0 1724 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_5866
timestamp 1745462530
transform 1 0 1708 0 1 1295
box -3 -3 3 3
use M3_M2  M3_M2_5867
timestamp 1745462530
transform 1 0 1660 0 1 1535
box -3 -3 3 3
use M3_M2  M3_M2_5868
timestamp 1745462530
transform 1 0 1644 0 1 1535
box -3 -3 3 3
use M3_M2  M3_M2_5869
timestamp 1745462530
transform 1 0 1556 0 1 1535
box -3 -3 3 3
use M3_M2  M3_M2_5870
timestamp 1745462530
transform 1 0 1508 0 1 1525
box -3 -3 3 3
use M3_M2  M3_M2_5871
timestamp 1745462530
transform 1 0 1948 0 1 1375
box -3 -3 3 3
use M3_M2  M3_M2_5872
timestamp 1745462530
transform 1 0 1892 0 1 1375
box -3 -3 3 3
use M3_M2  M3_M2_5873
timestamp 1745462530
transform 1 0 2164 0 1 1275
box -3 -3 3 3
use M3_M2  M3_M2_5874
timestamp 1745462530
transform 1 0 2108 0 1 1275
box -3 -3 3 3
use M3_M2  M3_M2_5875
timestamp 1745462530
transform 1 0 2068 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_5876
timestamp 1745462530
transform 1 0 2068 0 1 1275
box -3 -3 3 3
use M3_M2  M3_M2_5877
timestamp 1745462530
transform 1 0 2052 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_5878
timestamp 1745462530
transform 1 0 1460 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_5879
timestamp 1745462530
transform 1 0 1284 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_5880
timestamp 1745462530
transform 1 0 1252 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_5881
timestamp 1745462530
transform 1 0 2100 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_5882
timestamp 1745462530
transform 1 0 1972 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_5883
timestamp 1745462530
transform 1 0 1340 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_5884
timestamp 1745462530
transform 1 0 1340 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_5885
timestamp 1745462530
transform 1 0 1220 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_5886
timestamp 1745462530
transform 1 0 1796 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_5887
timestamp 1745462530
transform 1 0 1748 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_5888
timestamp 1745462530
transform 1 0 1636 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_5889
timestamp 1745462530
transform 1 0 1636 0 1 1135
box -3 -3 3 3
use M3_M2  M3_M2_5890
timestamp 1745462530
transform 1 0 1588 0 1 1135
box -3 -3 3 3
use M3_M2  M3_M2_5891
timestamp 1745462530
transform 1 0 1580 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_5892
timestamp 1745462530
transform 1 0 1532 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_5893
timestamp 1745462530
transform 1 0 1484 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_5894
timestamp 1745462530
transform 1 0 1972 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_5895
timestamp 1745462530
transform 1 0 1924 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_5896
timestamp 1745462530
transform 1 0 1924 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_5897
timestamp 1745462530
transform 1 0 1884 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_5898
timestamp 1745462530
transform 1 0 2228 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_5899
timestamp 1745462530
transform 1 0 2188 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_5900
timestamp 1745462530
transform 1 0 2116 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_5901
timestamp 1745462530
transform 1 0 2028 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_5902
timestamp 1745462530
transform 1 0 1396 0 1 1335
box -3 -3 3 3
use M3_M2  M3_M2_5903
timestamp 1745462530
transform 1 0 1244 0 1 1335
box -3 -3 3 3
use M3_M2  M3_M2_5904
timestamp 1745462530
transform 1 0 1244 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_5905
timestamp 1745462530
transform 1 0 1148 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_5906
timestamp 1745462530
transform 1 0 1372 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_5907
timestamp 1745462530
transform 1 0 1324 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_5908
timestamp 1745462530
transform 1 0 1252 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_5909
timestamp 1745462530
transform 1 0 1036 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_5910
timestamp 1745462530
transform 1 0 1828 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_5911
timestamp 1745462530
transform 1 0 1764 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_5912
timestamp 1745462530
transform 1 0 1700 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_5913
timestamp 1745462530
transform 1 0 1700 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_5914
timestamp 1745462530
transform 1 0 1604 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_5915
timestamp 1745462530
transform 1 0 1556 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_5916
timestamp 1745462530
transform 1 0 1500 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_5917
timestamp 1745462530
transform 1 0 1396 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_5918
timestamp 1745462530
transform 1 0 1972 0 1 1015
box -3 -3 3 3
use M3_M2  M3_M2_5919
timestamp 1745462530
transform 1 0 1924 0 1 1075
box -3 -3 3 3
use M3_M2  M3_M2_5920
timestamp 1745462530
transform 1 0 1924 0 1 1015
box -3 -3 3 3
use M3_M2  M3_M2_5921
timestamp 1745462530
transform 1 0 1836 0 1 1075
box -3 -3 3 3
use M3_M2  M3_M2_5922
timestamp 1745462530
transform 1 0 2140 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_5923
timestamp 1745462530
transform 1 0 2092 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_5924
timestamp 1745462530
transform 1 0 1988 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_5925
timestamp 1745462530
transform 1 0 1980 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_5926
timestamp 1745462530
transform 1 0 1964 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_5927
timestamp 1745462530
transform 1 0 1372 0 1 975
box -3 -3 3 3
use M3_M2  M3_M2_5928
timestamp 1745462530
transform 1 0 1252 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_5929
timestamp 1745462530
transform 1 0 1252 0 1 975
box -3 -3 3 3
use M3_M2  M3_M2_5930
timestamp 1745462530
transform 1 0 1116 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_5931
timestamp 1745462530
transform 1 0 1372 0 1 885
box -3 -3 3 3
use M3_M2  M3_M2_5932
timestamp 1745462530
transform 1 0 1252 0 1 885
box -3 -3 3 3
use M3_M2  M3_M2_5933
timestamp 1745462530
transform 1 0 1116 0 1 885
box -3 -3 3 3
use M3_M2  M3_M2_5934
timestamp 1745462530
transform 1 0 1796 0 1 535
box -3 -3 3 3
use M3_M2  M3_M2_5935
timestamp 1745462530
transform 1 0 1796 0 1 375
box -3 -3 3 3
use M3_M2  M3_M2_5936
timestamp 1745462530
transform 1 0 1684 0 1 375
box -3 -3 3 3
use M3_M2  M3_M2_5937
timestamp 1745462530
transform 1 0 1612 0 1 535
box -3 -3 3 3
use M3_M2  M3_M2_5938
timestamp 1745462530
transform 1 0 1652 0 1 155
box -3 -3 3 3
use M3_M2  M3_M2_5939
timestamp 1745462530
transform 1 0 1548 0 1 495
box -3 -3 3 3
use M3_M2  M3_M2_5940
timestamp 1745462530
transform 1 0 1540 0 1 155
box -3 -3 3 3
use M3_M2  M3_M2_5941
timestamp 1745462530
transform 1 0 1484 0 1 495
box -3 -3 3 3
use M3_M2  M3_M2_5942
timestamp 1745462530
transform 1 0 2060 0 1 155
box -3 -3 3 3
use M3_M2  M3_M2_5943
timestamp 1745462530
transform 1 0 1948 0 1 155
box -3 -3 3 3
use M3_M2  M3_M2_5944
timestamp 1745462530
transform 1 0 1940 0 1 405
box -3 -3 3 3
use M3_M2  M3_M2_5945
timestamp 1745462530
transform 1 0 1884 0 1 775
box -3 -3 3 3
use M3_M2  M3_M2_5946
timestamp 1745462530
transform 1 0 1788 0 1 405
box -3 -3 3 3
use M3_M2  M3_M2_5947
timestamp 1745462530
transform 1 0 1772 0 1 775
box -3 -3 3 3
use M3_M2  M3_M2_5948
timestamp 1745462530
transform 1 0 2068 0 1 335
box -3 -3 3 3
use M3_M2  M3_M2_5949
timestamp 1745462530
transform 1 0 2028 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_5950
timestamp 1745462530
transform 1 0 2020 0 1 335
box -3 -3 3 3
use M3_M2  M3_M2_5951
timestamp 1745462530
transform 1 0 1996 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_5952
timestamp 1745462530
transform 1 0 1956 0 1 335
box -3 -3 3 3
use M3_M2  M3_M2_5953
timestamp 1745462530
transform 1 0 1948 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_5954
timestamp 1745462530
transform 1 0 1356 0 1 375
box -3 -3 3 3
use M3_M2  M3_M2_5955
timestamp 1745462530
transform 1 0 1348 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_5956
timestamp 1745462530
transform 1 0 1340 0 1 405
box -3 -3 3 3
use M3_M2  M3_M2_5957
timestamp 1745462530
transform 1 0 1308 0 1 405
box -3 -3 3 3
use M3_M2  M3_M2_5958
timestamp 1745462530
transform 1 0 1308 0 1 375
box -3 -3 3 3
use M3_M2  M3_M2_5959
timestamp 1745462530
transform 1 0 1196 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_5960
timestamp 1745462530
transform 1 0 1108 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_5961
timestamp 1745462530
transform 1 0 1108 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_5962
timestamp 1745462530
transform 1 0 1076 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_5963
timestamp 1745462530
transform 1 0 1228 0 1 865
box -3 -3 3 3
use M3_M2  M3_M2_5964
timestamp 1745462530
transform 1 0 1196 0 1 865
box -3 -3 3 3
use M3_M2  M3_M2_5965
timestamp 1745462530
transform 1 0 1044 0 1 865
box -3 -3 3 3
use M3_M2  M3_M2_5966
timestamp 1745462530
transform 1 0 1756 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_5967
timestamp 1745462530
transform 1 0 1676 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_5968
timestamp 1745462530
transform 1 0 1468 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_5969
timestamp 1745462530
transform 1 0 1404 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_5970
timestamp 1745462530
transform 1 0 1900 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_5971
timestamp 1745462530
transform 1 0 1788 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_5972
timestamp 1745462530
transform 1 0 2124 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_5973
timestamp 1745462530
transform 1 0 2060 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_5974
timestamp 1745462530
transform 1 0 1940 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_5975
timestamp 1745462530
transform 1 0 1268 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_5976
timestamp 1745462530
transform 1 0 1220 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_5977
timestamp 1745462530
transform 1 0 1204 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_5978
timestamp 1745462530
transform 1 0 1172 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_5979
timestamp 1745462530
transform 1 0 1460 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_5980
timestamp 1745462530
transform 1 0 1412 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_5981
timestamp 1745462530
transform 1 0 2060 0 1 205
box -3 -3 3 3
use M3_M2  M3_M2_5982
timestamp 1745462530
transform 1 0 1956 0 1 205
box -3 -3 3 3
use M3_M2  M3_M2_5983
timestamp 1745462530
transform 1 0 1276 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_5984
timestamp 1745462530
transform 1 0 1212 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_5985
timestamp 1745462530
transform 1 0 1332 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_5986
timestamp 1745462530
transform 1 0 1220 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_5987
timestamp 1745462530
transform 1 0 1828 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_5988
timestamp 1745462530
transform 1 0 1724 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_5989
timestamp 1745462530
transform 1 0 1580 0 1 535
box -3 -3 3 3
use M3_M2  M3_M2_5990
timestamp 1745462530
transform 1 0 1540 0 1 535
box -3 -3 3 3
use M3_M2  M3_M2_5991
timestamp 1745462530
transform 1 0 1476 0 1 535
box -3 -3 3 3
use M3_M2  M3_M2_5992
timestamp 1745462530
transform 1 0 1892 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_5993
timestamp 1745462530
transform 1 0 1852 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_5994
timestamp 1745462530
transform 1 0 1844 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_5995
timestamp 1745462530
transform 1 0 1820 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_5996
timestamp 1745462530
transform 1 0 2132 0 1 605
box -3 -3 3 3
use M3_M2  M3_M2_5997
timestamp 1745462530
transform 1 0 2052 0 1 605
box -3 -3 3 3
use M3_M2  M3_M2_5998
timestamp 1745462530
transform 1 0 1108 0 1 575
box -3 -3 3 3
use M3_M2  M3_M2_5999
timestamp 1745462530
transform 1 0 1084 0 1 575
box -3 -3 3 3
use M3_M2  M3_M2_6000
timestamp 1745462530
transform 1 0 1044 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_6001
timestamp 1745462530
transform 1 0 1044 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_6002
timestamp 1745462530
transform 1 0 996 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_6003
timestamp 1745462530
transform 1 0 980 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_6004
timestamp 1745462530
transform 1 0 1652 0 1 325
box -3 -3 3 3
use M3_M2  M3_M2_6005
timestamp 1745462530
transform 1 0 1572 0 1 325
box -3 -3 3 3
use M3_M2  M3_M2_6006
timestamp 1745462530
transform 1 0 924 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_6007
timestamp 1745462530
transform 1 0 772 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_6008
timestamp 1745462530
transform 1 0 668 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_6009
timestamp 1745462530
transform 1 0 668 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_6010
timestamp 1745462530
transform 1 0 644 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_6011
timestamp 1745462530
transform 1 0 996 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_6012
timestamp 1745462530
transform 1 0 740 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_6013
timestamp 1745462530
transform 1 0 740 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_6014
timestamp 1745462530
transform 1 0 724 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_6015
timestamp 1745462530
transform 1 0 660 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_6016
timestamp 1745462530
transform 1 0 660 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_6017
timestamp 1745462530
transform 1 0 932 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_6018
timestamp 1745462530
transform 1 0 764 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_6019
timestamp 1745462530
transform 1 0 1020 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_6020
timestamp 1745462530
transform 1 0 900 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_6021
timestamp 1745462530
transform 1 0 900 0 1 1435
box -3 -3 3 3
use M3_M2  M3_M2_6022
timestamp 1745462530
transform 1 0 836 0 1 1435
box -3 -3 3 3
use M3_M2  M3_M2_6023
timestamp 1745462530
transform 1 0 1148 0 1 1285
box -3 -3 3 3
use M3_M2  M3_M2_6024
timestamp 1745462530
transform 1 0 1100 0 1 1285
box -3 -3 3 3
use M3_M2  M3_M2_6025
timestamp 1745462530
transform 1 0 1012 0 1 1285
box -3 -3 3 3
use M3_M2  M3_M2_6026
timestamp 1745462530
transform 1 0 988 0 1 1285
box -3 -3 3 3
use M3_M2  M3_M2_6027
timestamp 1745462530
transform 1 0 1084 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_6028
timestamp 1745462530
transform 1 0 908 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_6029
timestamp 1745462530
transform 1 0 900 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_6030
timestamp 1745462530
transform 1 0 836 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_6031
timestamp 1745462530
transform 1 0 628 0 1 1285
box -3 -3 3 3
use M3_M2  M3_M2_6032
timestamp 1745462530
transform 1 0 540 0 1 1285
box -3 -3 3 3
use M3_M2  M3_M2_6033
timestamp 1745462530
transform 1 0 524 0 1 1285
box -3 -3 3 3
use M3_M2  M3_M2_6034
timestamp 1745462530
transform 1 0 668 0 1 1135
box -3 -3 3 3
use M3_M2  M3_M2_6035
timestamp 1745462530
transform 1 0 612 0 1 1135
box -3 -3 3 3
use M3_M2  M3_M2_6036
timestamp 1745462530
transform 1 0 540 0 1 1135
box -3 -3 3 3
use M3_M2  M3_M2_6037
timestamp 1745462530
transform 1 0 420 0 1 1135
box -3 -3 3 3
use M3_M2  M3_M2_6038
timestamp 1745462530
transform 1 0 708 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_6039
timestamp 1745462530
transform 1 0 596 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_6040
timestamp 1745462530
transform 1 0 364 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_6041
timestamp 1745462530
transform 1 0 788 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_6042
timestamp 1745462530
transform 1 0 748 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_6043
timestamp 1745462530
transform 1 0 196 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_6044
timestamp 1745462530
transform 1 0 148 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_6045
timestamp 1745462530
transform 1 0 148 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_6046
timestamp 1745462530
transform 1 0 956 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_6047
timestamp 1745462530
transform 1 0 908 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_6048
timestamp 1745462530
transform 1 0 908 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_6049
timestamp 1745462530
transform 1 0 180 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_6050
timestamp 1745462530
transform 1 0 908 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_6051
timestamp 1745462530
transform 1 0 780 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_6052
timestamp 1745462530
transform 1 0 460 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_6053
timestamp 1745462530
transform 1 0 844 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_6054
timestamp 1745462530
transform 1 0 828 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_6055
timestamp 1745462530
transform 1 0 724 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_6056
timestamp 1745462530
transform 1 0 724 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_6057
timestamp 1745462530
transform 1 0 1020 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_6058
timestamp 1745462530
transform 1 0 1004 0 1 205
box -3 -3 3 3
use M3_M2  M3_M2_6059
timestamp 1745462530
transform 1 0 980 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_6060
timestamp 1745462530
transform 1 0 940 0 1 205
box -3 -3 3 3
use M3_M2  M3_M2_6061
timestamp 1745462530
transform 1 0 716 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_6062
timestamp 1745462530
transform 1 0 964 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_6063
timestamp 1745462530
transform 1 0 900 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_6064
timestamp 1745462530
transform 1 0 900 0 1 485
box -3 -3 3 3
use M3_M2  M3_M2_6065
timestamp 1745462530
transform 1 0 868 0 1 485
box -3 -3 3 3
use M3_M2  M3_M2_6066
timestamp 1745462530
transform 1 0 804 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_6067
timestamp 1745462530
transform 1 0 980 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_6068
timestamp 1745462530
transform 1 0 972 0 1 375
box -3 -3 3 3
use M3_M2  M3_M2_6069
timestamp 1745462530
transform 1 0 956 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_6070
timestamp 1745462530
transform 1 0 940 0 1 375
box -3 -3 3 3
use M3_M2  M3_M2_6071
timestamp 1745462530
transform 1 0 964 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_6072
timestamp 1745462530
transform 1 0 948 0 1 665
box -3 -3 3 3
use M3_M2  M3_M2_6073
timestamp 1745462530
transform 1 0 948 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_6074
timestamp 1745462530
transform 1 0 924 0 1 665
box -3 -3 3 3
use M3_M2  M3_M2_6075
timestamp 1745462530
transform 1 0 1004 0 1 845
box -3 -3 3 3
use M3_M2  M3_M2_6076
timestamp 1745462530
transform 1 0 820 0 1 845
box -3 -3 3 3
use M3_M2  M3_M2_6077
timestamp 1745462530
transform 1 0 820 0 1 375
box -3 -3 3 3
use M3_M2  M3_M2_6078
timestamp 1745462530
transform 1 0 804 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_6079
timestamp 1745462530
transform 1 0 780 0 1 375
box -3 -3 3 3
use M3_M2  M3_M2_6080
timestamp 1745462530
transform 1 0 780 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_6081
timestamp 1745462530
transform 1 0 772 0 1 105
box -3 -3 3 3
use M3_M2  M3_M2_6082
timestamp 1745462530
transform 1 0 668 0 1 105
box -3 -3 3 3
use M3_M2  M3_M2_6083
timestamp 1745462530
transform 1 0 612 0 1 105
box -3 -3 3 3
use M3_M2  M3_M2_6084
timestamp 1745462530
transform 1 0 716 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_6085
timestamp 1745462530
transform 1 0 572 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_6086
timestamp 1745462530
transform 1 0 916 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_6087
timestamp 1745462530
transform 1 0 892 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_6088
timestamp 1745462530
transform 1 0 844 0 1 405
box -3 -3 3 3
use M3_M2  M3_M2_6089
timestamp 1745462530
transform 1 0 804 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_6090
timestamp 1745462530
transform 1 0 756 0 1 405
box -3 -3 3 3
use M3_M2  M3_M2_6091
timestamp 1745462530
transform 1 0 844 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_6092
timestamp 1745462530
transform 1 0 740 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_6093
timestamp 1745462530
transform 1 0 780 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_6094
timestamp 1745462530
transform 1 0 756 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_6095
timestamp 1745462530
transform 1 0 748 0 1 325
box -3 -3 3 3
use M3_M2  M3_M2_6096
timestamp 1745462530
transform 1 0 700 0 1 325
box -3 -3 3 3
use M3_M2  M3_M2_6097
timestamp 1745462530
transform 1 0 668 0 1 325
box -3 -3 3 3
use M3_M2  M3_M2_6098
timestamp 1745462530
transform 1 0 900 0 1 975
box -3 -3 3 3
use M3_M2  M3_M2_6099
timestamp 1745462530
transform 1 0 764 0 1 975
box -3 -3 3 3
use M3_M2  M3_M2_6100
timestamp 1745462530
transform 1 0 764 0 1 535
box -3 -3 3 3
use M3_M2  M3_M2_6101
timestamp 1745462530
transform 1 0 652 0 1 535
box -3 -3 3 3
use M3_M2  M3_M2_6102
timestamp 1745462530
transform 1 0 620 0 1 535
box -3 -3 3 3
use M3_M2  M3_M2_6103
timestamp 1745462530
transform 1 0 1068 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_6104
timestamp 1745462530
transform 1 0 476 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_6105
timestamp 1745462530
transform 1 0 1012 0 1 415
box -3 -3 3 3
use M3_M2  M3_M2_6106
timestamp 1745462530
transform 1 0 372 0 1 415
box -3 -3 3 3
use M3_M2  M3_M2_6107
timestamp 1745462530
transform 1 0 1036 0 1 775
box -3 -3 3 3
use M3_M2  M3_M2_6108
timestamp 1745462530
transform 1 0 276 0 1 415
box -3 -3 3 3
use M3_M2  M3_M2_6109
timestamp 1745462530
transform 1 0 260 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_6110
timestamp 1745462530
transform 1 0 172 0 1 415
box -3 -3 3 3
use M3_M2  M3_M2_6111
timestamp 1745462530
transform 1 0 980 0 1 885
box -3 -3 3 3
use M3_M2  M3_M2_6112
timestamp 1745462530
transform 1 0 300 0 1 645
box -3 -3 3 3
use M3_M2  M3_M2_6113
timestamp 1745462530
transform 1 0 292 0 1 885
box -3 -3 3 3
use M3_M2  M3_M2_6114
timestamp 1745462530
transform 1 0 180 0 1 645
box -3 -3 3 3
use M3_M2  M3_M2_6115
timestamp 1745462530
transform 1 0 1052 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_6116
timestamp 1745462530
transform 1 0 588 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_6117
timestamp 1745462530
transform 1 0 588 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_6118
timestamp 1745462530
transform 1 0 532 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_6119
timestamp 1745462530
transform 1 0 508 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_6120
timestamp 1745462530
transform 1 0 284 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_6121
timestamp 1745462530
transform 1 0 180 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_6122
timestamp 1745462530
transform 1 0 548 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_6123
timestamp 1745462530
transform 1 0 428 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_6124
timestamp 1745462530
transform 1 0 564 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_6125
timestamp 1745462530
transform 1 0 420 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_6126
timestamp 1745462530
transform 1 0 420 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_6127
timestamp 1745462530
transform 1 0 356 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_6128
timestamp 1745462530
transform 1 0 708 0 1 975
box -3 -3 3 3
use M3_M2  M3_M2_6129
timestamp 1745462530
transform 1 0 316 0 1 975
box -3 -3 3 3
use M3_M2  M3_M2_6130
timestamp 1745462530
transform 1 0 316 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_6131
timestamp 1745462530
transform 1 0 236 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_6132
timestamp 1745462530
transform 1 0 188 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_6133
timestamp 1745462530
transform 1 0 844 0 1 1015
box -3 -3 3 3
use M3_M2  M3_M2_6134
timestamp 1745462530
transform 1 0 244 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_6135
timestamp 1745462530
transform 1 0 180 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_6136
timestamp 1745462530
transform 1 0 844 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_6137
timestamp 1745462530
transform 1 0 412 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_6138
timestamp 1745462530
transform 1 0 348 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_6139
timestamp 1745462530
transform 1 0 332 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_6140
timestamp 1745462530
transform 1 0 940 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_6141
timestamp 1745462530
transform 1 0 756 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_6142
timestamp 1745462530
transform 1 0 668 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_6143
timestamp 1745462530
transform 1 0 668 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_6144
timestamp 1745462530
transform 1 0 620 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_6145
timestamp 1745462530
transform 1 0 988 0 1 1865
box -3 -3 3 3
use M3_M2  M3_M2_6146
timestamp 1745462530
transform 1 0 916 0 1 1865
box -3 -3 3 3
use M3_M2  M3_M2_6147
timestamp 1745462530
transform 1 0 812 0 1 1865
box -3 -3 3 3
use M3_M2  M3_M2_6148
timestamp 1745462530
transform 1 0 900 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_6149
timestamp 1745462530
transform 1 0 756 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_6150
timestamp 1745462530
transform 1 0 748 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_6151
timestamp 1745462530
transform 1 0 676 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_6152
timestamp 1745462530
transform 1 0 628 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_6153
timestamp 1745462530
transform 1 0 900 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_6154
timestamp 1745462530
transform 1 0 836 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_6155
timestamp 1745462530
transform 1 0 724 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_6156
timestamp 1745462530
transform 1 0 980 0 1 1615
box -3 -3 3 3
use M3_M2  M3_M2_6157
timestamp 1745462530
transform 1 0 868 0 1 1615
box -3 -3 3 3
use M3_M2  M3_M2_6158
timestamp 1745462530
transform 1 0 748 0 1 1615
box -3 -3 3 3
use M3_M2  M3_M2_6159
timestamp 1745462530
transform 1 0 852 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_6160
timestamp 1745462530
transform 1 0 836 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_6161
timestamp 1745462530
transform 1 0 580 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_6162
timestamp 1745462530
transform 1 0 692 0 1 2095
box -3 -3 3 3
use M3_M2  M3_M2_6163
timestamp 1745462530
transform 1 0 548 0 1 2095
box -3 -3 3 3
use M3_M2  M3_M2_6164
timestamp 1745462530
transform 1 0 316 0 1 2095
box -3 -3 3 3
use M3_M2  M3_M2_6165
timestamp 1745462530
transform 1 0 820 0 1 2285
box -3 -3 3 3
use M3_M2  M3_M2_6166
timestamp 1745462530
transform 1 0 820 0 1 2065
box -3 -3 3 3
use M3_M2  M3_M2_6167
timestamp 1745462530
transform 1 0 764 0 1 2065
box -3 -3 3 3
use M3_M2  M3_M2_6168
timestamp 1745462530
transform 1 0 764 0 1 1885
box -3 -3 3 3
use M3_M2  M3_M2_6169
timestamp 1745462530
transform 1 0 668 0 1 2285
box -3 -3 3 3
use M3_M2  M3_M2_6170
timestamp 1745462530
transform 1 0 452 0 1 1885
box -3 -3 3 3
use M3_M2  M3_M2_6171
timestamp 1745462530
transform 1 0 644 0 1 1685
box -3 -3 3 3
use M3_M2  M3_M2_6172
timestamp 1745462530
transform 1 0 524 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_6173
timestamp 1745462530
transform 1 0 524 0 1 1685
box -3 -3 3 3
use M3_M2  M3_M2_6174
timestamp 1745462530
transform 1 0 468 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_6175
timestamp 1745462530
transform 1 0 836 0 1 1845
box -3 -3 3 3
use M3_M2  M3_M2_6176
timestamp 1745462530
transform 1 0 748 0 1 2295
box -3 -3 3 3
use M3_M2  M3_M2_6177
timestamp 1745462530
transform 1 0 708 0 1 2295
box -3 -3 3 3
use M3_M2  M3_M2_6178
timestamp 1745462530
transform 1 0 700 0 1 1845
box -3 -3 3 3
use M3_M2  M3_M2_6179
timestamp 1745462530
transform 1 0 380 0 1 1845
box -3 -3 3 3
use M3_M2  M3_M2_6180
timestamp 1745462530
transform 1 0 908 0 1 1885
box -3 -3 3 3
use M3_M2  M3_M2_6181
timestamp 1745462530
transform 1 0 884 0 1 2055
box -3 -3 3 3
use M3_M2  M3_M2_6182
timestamp 1745462530
transform 1 0 852 0 1 1885
box -3 -3 3 3
use M3_M2  M3_M2_6183
timestamp 1745462530
transform 1 0 852 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_6184
timestamp 1745462530
transform 1 0 820 0 1 2055
box -3 -3 3 3
use M3_M2  M3_M2_6185
timestamp 1745462530
transform 1 0 820 0 1 1885
box -3 -3 3 3
use M3_M2  M3_M2_6186
timestamp 1745462530
transform 1 0 268 0 1 1775
box -3 -3 3 3
use M3_M2  M3_M2_6187
timestamp 1745462530
transform 1 0 268 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_6188
timestamp 1745462530
transform 1 0 204 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_6189
timestamp 1745462530
transform 1 0 772 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_6190
timestamp 1745462530
transform 1 0 180 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_6191
timestamp 1745462530
transform 1 0 892 0 1 2205
box -3 -3 3 3
use M3_M2  M3_M2_6192
timestamp 1745462530
transform 1 0 652 0 1 2205
box -3 -3 3 3
use M3_M2  M3_M2_6193
timestamp 1745462530
transform 1 0 308 0 1 2205
box -3 -3 3 3
use M3_M2  M3_M2_6194
timestamp 1745462530
transform 1 0 1036 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_6195
timestamp 1745462530
transform 1 0 668 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_6196
timestamp 1745462530
transform 1 0 556 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_6197
timestamp 1745462530
transform 1 0 460 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_6198
timestamp 1745462530
transform 1 0 860 0 1 2155
box -3 -3 3 3
use M3_M2  M3_M2_6199
timestamp 1745462530
transform 1 0 628 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_6200
timestamp 1745462530
transform 1 0 500 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_6201
timestamp 1745462530
transform 1 0 932 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_6202
timestamp 1745462530
transform 1 0 828 0 1 2005
box -3 -3 3 3
use M3_M2  M3_M2_6203
timestamp 1745462530
transform 1 0 828 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_6204
timestamp 1745462530
transform 1 0 388 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_6205
timestamp 1745462530
transform 1 0 1020 0 1 2135
box -3 -3 3 3
use M3_M2  M3_M2_6206
timestamp 1745462530
transform 1 0 844 0 1 2135
box -3 -3 3 3
use M3_M2  M3_M2_6207
timestamp 1745462530
transform 1 0 172 0 1 2135
box -3 -3 3 3
use M3_M2  M3_M2_6208
timestamp 1745462530
transform 1 0 972 0 1 2095
box -3 -3 3 3
use M3_M2  M3_M2_6209
timestamp 1745462530
transform 1 0 812 0 1 2275
box -3 -3 3 3
use M3_M2  M3_M2_6210
timestamp 1745462530
transform 1 0 812 0 1 2095
box -3 -3 3 3
use M3_M2  M3_M2_6211
timestamp 1745462530
transform 1 0 812 0 1 2045
box -3 -3 3 3
use M3_M2  M3_M2_6212
timestamp 1745462530
transform 1 0 740 0 1 2275
box -3 -3 3 3
use M3_M2  M3_M2_6213
timestamp 1745462530
transform 1 0 180 0 1 2045
box -3 -3 3 3
use M3_M2  M3_M2_6214
timestamp 1745462530
transform 1 0 604 0 1 2275
box -3 -3 3 3
use M3_M2  M3_M2_6215
timestamp 1745462530
transform 1 0 540 0 1 2275
box -3 -3 3 3
use M3_M2  M3_M2_6216
timestamp 1745462530
transform 1 0 516 0 1 2375
box -3 -3 3 3
use M3_M2  M3_M2_6217
timestamp 1745462530
transform 1 0 364 0 1 2375
box -3 -3 3 3
use M3_M2  M3_M2_6218
timestamp 1745462530
transform 1 0 364 0 1 2355
box -3 -3 3 3
use M3_M2  M3_M2_6219
timestamp 1745462530
transform 1 0 308 0 1 2355
box -3 -3 3 3
use M3_M2  M3_M2_6220
timestamp 1745462530
transform 1 0 620 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_6221
timestamp 1745462530
transform 1 0 612 0 1 2465
box -3 -3 3 3
use M3_M2  M3_M2_6222
timestamp 1745462530
transform 1 0 588 0 1 2465
box -3 -3 3 3
use M3_M2  M3_M2_6223
timestamp 1745462530
transform 1 0 588 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_6224
timestamp 1745462530
transform 1 0 500 0 1 2485
box -3 -3 3 3
use M3_M2  M3_M2_6225
timestamp 1745462530
transform 1 0 436 0 1 2485
box -3 -3 3 3
use M3_M2  M3_M2_6226
timestamp 1745462530
transform 1 0 580 0 1 2385
box -3 -3 3 3
use M3_M2  M3_M2_6227
timestamp 1745462530
transform 1 0 508 0 1 2385
box -3 -3 3 3
use M3_M2  M3_M2_6228
timestamp 1745462530
transform 1 0 508 0 1 2355
box -3 -3 3 3
use M3_M2  M3_M2_6229
timestamp 1745462530
transform 1 0 388 0 1 2355
box -3 -3 3 3
use M3_M2  M3_M2_6230
timestamp 1745462530
transform 1 0 796 0 1 2265
box -3 -3 3 3
use M3_M2  M3_M2_6231
timestamp 1745462530
transform 1 0 796 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_6232
timestamp 1745462530
transform 1 0 772 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_6233
timestamp 1745462530
transform 1 0 756 0 1 2265
box -3 -3 3 3
use M3_M2  M3_M2_6234
timestamp 1745462530
transform 1 0 436 0 1 2265
box -3 -3 3 3
use M3_M2  M3_M2_6235
timestamp 1745462530
transform 1 0 436 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_6236
timestamp 1745462530
transform 1 0 364 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_6237
timestamp 1745462530
transform 1 0 852 0 1 2255
box -3 -3 3 3
use M3_M2  M3_M2_6238
timestamp 1745462530
transform 1 0 804 0 1 2255
box -3 -3 3 3
use M3_M2  M3_M2_6239
timestamp 1745462530
transform 1 0 180 0 1 2255
box -3 -3 3 3
use M3_M2  M3_M2_6240
timestamp 1745462530
transform 1 0 780 0 1 2425
box -3 -3 3 3
use M3_M2  M3_M2_6241
timestamp 1745462530
transform 1 0 692 0 1 2425
box -3 -3 3 3
use M3_M2  M3_M2_6242
timestamp 1745462530
transform 1 0 244 0 1 2405
box -3 -3 3 3
use M3_M2  M3_M2_6243
timestamp 1745462530
transform 1 0 172 0 1 2405
box -3 -3 3 3
use M3_M2  M3_M2_6244
timestamp 1745462530
transform 1 0 988 0 1 2365
box -3 -3 3 3
use M3_M2  M3_M2_6245
timestamp 1745462530
transform 1 0 940 0 1 2365
box -3 -3 3 3
use M3_M2  M3_M2_6246
timestamp 1745462530
transform 1 0 900 0 1 2365
box -3 -3 3 3
use M3_M2  M3_M2_6247
timestamp 1745462530
transform 1 0 1204 0 1 2835
box -3 -3 3 3
use M3_M2  M3_M2_6248
timestamp 1745462530
transform 1 0 1076 0 1 2075
box -3 -3 3 3
use M3_M2  M3_M2_6249
timestamp 1745462530
transform 1 0 1052 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_6250
timestamp 1745462530
transform 1 0 1052 0 1 2075
box -3 -3 3 3
use M3_M2  M3_M2_6251
timestamp 1745462530
transform 1 0 1036 0 1 2835
box -3 -3 3 3
use M3_M2  M3_M2_6252
timestamp 1745462530
transform 1 0 1036 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_6253
timestamp 1745462530
transform 1 0 1036 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_6254
timestamp 1745462530
transform 1 0 1004 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_6255
timestamp 1745462530
transform 1 0 1092 0 1 2575
box -3 -3 3 3
use M3_M2  M3_M2_6256
timestamp 1745462530
transform 1 0 924 0 1 2575
box -3 -3 3 3
use M3_M2  M3_M2_6257
timestamp 1745462530
transform 1 0 1092 0 1 2875
box -3 -3 3 3
use M3_M2  M3_M2_6258
timestamp 1745462530
transform 1 0 956 0 1 2075
box -3 -3 3 3
use M3_M2  M3_M2_6259
timestamp 1745462530
transform 1 0 908 0 1 2895
box -3 -3 3 3
use M3_M2  M3_M2_6260
timestamp 1745462530
transform 1 0 908 0 1 2875
box -3 -3 3 3
use M3_M2  M3_M2_6261
timestamp 1745462530
transform 1 0 348 0 1 2895
box -3 -3 3 3
use M3_M2  M3_M2_6262
timestamp 1745462530
transform 1 0 348 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_6263
timestamp 1745462530
transform 1 0 340 0 1 2075
box -3 -3 3 3
use M3_M2  M3_M2_6264
timestamp 1745462530
transform 1 0 332 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_6265
timestamp 1745462530
transform 1 0 1084 0 1 2655
box -3 -3 3 3
use M3_M2  M3_M2_6266
timestamp 1745462530
transform 1 0 1020 0 1 2655
box -3 -3 3 3
use M3_M2  M3_M2_6267
timestamp 1745462530
transform 1 0 1060 0 1 2705
box -3 -3 3 3
use M3_M2  M3_M2_6268
timestamp 1745462530
transform 1 0 1044 0 1 2705
box -3 -3 3 3
use M3_M2  M3_M2_6269
timestamp 1745462530
transform 1 0 1036 0 1 2065
box -3 -3 3 3
use M3_M2  M3_M2_6270
timestamp 1745462530
transform 1 0 1020 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_6271
timestamp 1745462530
transform 1 0 972 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_6272
timestamp 1745462530
transform 1 0 964 0 1 2705
box -3 -3 3 3
use M3_M2  M3_M2_6273
timestamp 1745462530
transform 1 0 964 0 1 2065
box -3 -3 3 3
use M3_M2  M3_M2_6274
timestamp 1745462530
transform 1 0 596 0 1 2375
box -3 -3 3 3
use M3_M2  M3_M2_6275
timestamp 1745462530
transform 1 0 532 0 1 2375
box -3 -3 3 3
use M3_M2  M3_M2_6276
timestamp 1745462530
transform 1 0 596 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_6277
timestamp 1745462530
transform 1 0 596 0 1 2185
box -3 -3 3 3
use M3_M2  M3_M2_6278
timestamp 1745462530
transform 1 0 564 0 1 2185
box -3 -3 3 3
use M3_M2  M3_M2_6279
timestamp 1745462530
transform 1 0 556 0 1 2615
box -3 -3 3 3
use M3_M2  M3_M2_6280
timestamp 1745462530
transform 1 0 556 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_6281
timestamp 1745462530
transform 1 0 492 0 1 2615
box -3 -3 3 3
use M3_M2  M3_M2_6282
timestamp 1745462530
transform 1 0 724 0 1 2875
box -3 -3 3 3
use M3_M2  M3_M2_6283
timestamp 1745462530
transform 1 0 716 0 1 2375
box -3 -3 3 3
use M3_M2  M3_M2_6284
timestamp 1745462530
transform 1 0 620 0 1 2405
box -3 -3 3 3
use M3_M2  M3_M2_6285
timestamp 1745462530
transform 1 0 620 0 1 2375
box -3 -3 3 3
use M3_M2  M3_M2_6286
timestamp 1745462530
transform 1 0 492 0 1 2875
box -3 -3 3 3
use M3_M2  M3_M2_6287
timestamp 1745462530
transform 1 0 484 0 1 2405
box -3 -3 3 3
use M3_M2  M3_M2_6288
timestamp 1745462530
transform 1 0 892 0 1 2535
box -3 -3 3 3
use M3_M2  M3_M2_6289
timestamp 1745462530
transform 1 0 860 0 1 2555
box -3 -3 3 3
use M3_M2  M3_M2_6290
timestamp 1745462530
transform 1 0 860 0 1 2535
box -3 -3 3 3
use M3_M2  M3_M2_6291
timestamp 1745462530
transform 1 0 812 0 1 2555
box -3 -3 3 3
use M3_M2  M3_M2_6292
timestamp 1745462530
transform 1 0 732 0 1 2535
box -3 -3 3 3
use M3_M2  M3_M2_6293
timestamp 1745462530
transform 1 0 572 0 1 2535
box -3 -3 3 3
use M3_M2  M3_M2_6294
timestamp 1745462530
transform 1 0 412 0 1 2855
box -3 -3 3 3
use M3_M2  M3_M2_6295
timestamp 1745462530
transform 1 0 364 0 1 2855
box -3 -3 3 3
use M3_M2  M3_M2_6296
timestamp 1745462530
transform 1 0 2004 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_6297
timestamp 1745462530
transform 1 0 1844 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_6298
timestamp 1745462530
transform 1 0 1316 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_6299
timestamp 1745462530
transform 1 0 1220 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_6300
timestamp 1745462530
transform 1 0 1636 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_6301
timestamp 1745462530
transform 1 0 1524 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_6302
timestamp 1745462530
transform 1 0 1972 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_6303
timestamp 1745462530
transform 1 0 1972 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_6304
timestamp 1745462530
transform 1 0 1908 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_6305
timestamp 1745462530
transform 1 0 1852 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_6306
timestamp 1745462530
transform 1 0 1204 0 1 1975
box -3 -3 3 3
use M3_M2  M3_M2_6307
timestamp 1745462530
transform 1 0 1148 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_6308
timestamp 1745462530
transform 1 0 1124 0 1 1975
box -3 -3 3 3
use M3_M2  M3_M2_6309
timestamp 1745462530
transform 1 0 1116 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_6310
timestamp 1745462530
transform 1 0 1372 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_6311
timestamp 1745462530
transform 1 0 1340 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_6312
timestamp 1745462530
transform 1 0 2036 0 1 2475
box -3 -3 3 3
use M3_M2  M3_M2_6313
timestamp 1745462530
transform 1 0 1820 0 1 2475
box -3 -3 3 3
use M3_M2  M3_M2_6314
timestamp 1745462530
transform 1 0 1372 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_6315
timestamp 1745462530
transform 1 0 1276 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_6316
timestamp 1745462530
transform 1 0 1684 0 1 2565
box -3 -3 3 3
use M3_M2  M3_M2_6317
timestamp 1745462530
transform 1 0 1660 0 1 2565
box -3 -3 3 3
use M3_M2  M3_M2_6318
timestamp 1745462530
transform 1 0 1572 0 1 2565
box -3 -3 3 3
use M3_M2  M3_M2_6319
timestamp 1745462530
transform 1 0 1996 0 1 2545
box -3 -3 3 3
use M3_M2  M3_M2_6320
timestamp 1745462530
transform 1 0 1812 0 1 2545
box -3 -3 3 3
use M3_M2  M3_M2_6321
timestamp 1745462530
transform 1 0 1180 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_6322
timestamp 1745462530
transform 1 0 1156 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_6323
timestamp 1745462530
transform 1 0 1500 0 1 2685
box -3 -3 3 3
use M3_M2  M3_M2_6324
timestamp 1745462530
transform 1 0 1468 0 1 2685
box -3 -3 3 3
use M3_M2  M3_M2_6325
timestamp 1745462530
transform 1 0 1396 0 1 2685
box -3 -3 3 3
use M3_M2  M3_M2_6326
timestamp 1745462530
transform 1 0 2172 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_6327
timestamp 1745462530
transform 1 0 2036 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_6328
timestamp 1745462530
transform 1 0 2004 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_6329
timestamp 1745462530
transform 1 0 1388 0 1 1975
box -3 -3 3 3
use M3_M2  M3_M2_6330
timestamp 1745462530
transform 1 0 1316 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_6331
timestamp 1745462530
transform 1 0 1764 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_6332
timestamp 1745462530
transform 1 0 1644 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_6333
timestamp 1745462530
transform 1 0 2060 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_6334
timestamp 1745462530
transform 1 0 1900 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_6335
timestamp 1745462530
transform 1 0 1132 0 1 2155
box -3 -3 3 3
use M3_M2  M3_M2_6336
timestamp 1745462530
transform 1 0 1084 0 1 2155
box -3 -3 3 3
use M3_M2  M3_M2_6337
timestamp 1745462530
transform 1 0 2092 0 1 2545
box -3 -3 3 3
use M3_M2  M3_M2_6338
timestamp 1745462530
transform 1 0 2020 0 1 2545
box -3 -3 3 3
use M3_M2  M3_M2_6339
timestamp 1745462530
transform 1 0 1324 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_6340
timestamp 1745462530
transform 1 0 1308 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_6341
timestamp 1745462530
transform 1 0 1844 0 1 2725
box -3 -3 3 3
use M3_M2  M3_M2_6342
timestamp 1745462530
transform 1 0 1844 0 1 2705
box -3 -3 3 3
use M3_M2  M3_M2_6343
timestamp 1745462530
transform 1 0 1820 0 1 2705
box -3 -3 3 3
use M3_M2  M3_M2_6344
timestamp 1745462530
transform 1 0 1644 0 1 2725
box -3 -3 3 3
use M3_M2  M3_M2_6345
timestamp 1745462530
transform 1 0 1628 0 1 2725
box -3 -3 3 3
use M3_M2  M3_M2_6346
timestamp 1745462530
transform 1 0 1948 0 1 2705
box -3 -3 3 3
use M3_M2  M3_M2_6347
timestamp 1745462530
transform 1 0 1868 0 1 2705
box -3 -3 3 3
use M3_M2  M3_M2_6348
timestamp 1745462530
transform 1 0 1204 0 1 2705
box -3 -3 3 3
use M3_M2  M3_M2_6349
timestamp 1745462530
transform 1 0 1164 0 1 2705
box -3 -3 3 3
use M3_M2  M3_M2_6350
timestamp 1745462530
transform 1 0 1604 0 1 2765
box -3 -3 3 3
use M3_M2  M3_M2_6351
timestamp 1745462530
transform 1 0 1604 0 1 2705
box -3 -3 3 3
use M3_M2  M3_M2_6352
timestamp 1745462530
transform 1 0 1516 0 1 2705
box -3 -3 3 3
use M3_M2  M3_M2_6353
timestamp 1745462530
transform 1 0 1468 0 1 2765
box -3 -3 3 3
use M3_M2  M3_M2_6354
timestamp 1745462530
transform 1 0 2132 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_6355
timestamp 1745462530
transform 1 0 2068 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_6356
timestamp 1745462530
transform 1 0 2036 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_6357
timestamp 1745462530
transform 1 0 1396 0 1 2265
box -3 -3 3 3
use M3_M2  M3_M2_6358
timestamp 1745462530
transform 1 0 1364 0 1 2185
box -3 -3 3 3
use M3_M2  M3_M2_6359
timestamp 1745462530
transform 1 0 1340 0 1 2265
box -3 -3 3 3
use M3_M2  M3_M2_6360
timestamp 1745462530
transform 1 0 1340 0 1 2185
box -3 -3 3 3
use M3_M2  M3_M2_6361
timestamp 1745462530
transform 1 0 1748 0 1 2165
box -3 -3 3 3
use M3_M2  M3_M2_6362
timestamp 1745462530
transform 1 0 1732 0 1 2165
box -3 -3 3 3
use M3_M2  M3_M2_6363
timestamp 1745462530
transform 1 0 1732 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_6364
timestamp 1745462530
transform 1 0 1724 0 1 2315
box -3 -3 3 3
use M3_M2  M3_M2_6365
timestamp 1745462530
transform 1 0 1700 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_6366
timestamp 1745462530
transform 1 0 1692 0 1 2315
box -3 -3 3 3
use M3_M2  M3_M2_6367
timestamp 1745462530
transform 1 0 1668 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_6368
timestamp 1745462530
transform 1 0 1988 0 1 2125
box -3 -3 3 3
use M3_M2  M3_M2_6369
timestamp 1745462530
transform 1 0 1948 0 1 2125
box -3 -3 3 3
use M3_M2  M3_M2_6370
timestamp 1745462530
transform 1 0 1236 0 1 2385
box -3 -3 3 3
use M3_M2  M3_M2_6371
timestamp 1745462530
transform 1 0 1188 0 1 2385
box -3 -3 3 3
use M3_M2  M3_M2_6372
timestamp 1745462530
transform 1 0 1188 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_6373
timestamp 1745462530
transform 1 0 1124 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_6374
timestamp 1745462530
transform 1 0 1628 0 1 2165
box -3 -3 3 3
use M3_M2  M3_M2_6375
timestamp 1745462530
transform 1 0 1556 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_6376
timestamp 1745462530
transform 1 0 1516 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_6377
timestamp 1745462530
transform 1 0 1516 0 1 2165
box -3 -3 3 3
use M3_M2  M3_M2_6378
timestamp 1745462530
transform 1 0 2020 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_6379
timestamp 1745462530
transform 1 0 1980 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_6380
timestamp 1745462530
transform 1 0 1980 0 1 2635
box -3 -3 3 3
use M3_M2  M3_M2_6381
timestamp 1745462530
transform 1 0 1964 0 1 2635
box -3 -3 3 3
use M3_M2  M3_M2_6382
timestamp 1745462530
transform 1 0 1420 0 1 2905
box -3 -3 3 3
use M3_M2  M3_M2_6383
timestamp 1745462530
transform 1 0 1380 0 1 2905
box -3 -3 3 3
use M3_M2  M3_M2_6384
timestamp 1745462530
transform 1 0 1380 0 1 2565
box -3 -3 3 3
use M3_M2  M3_M2_6385
timestamp 1745462530
transform 1 0 1348 0 1 2565
box -3 -3 3 3
use M3_M2  M3_M2_6386
timestamp 1745462530
transform 1 0 1788 0 1 2815
box -3 -3 3 3
use M3_M2  M3_M2_6387
timestamp 1745462530
transform 1 0 1772 0 1 2525
box -3 -3 3 3
use M3_M2  M3_M2_6388
timestamp 1745462530
transform 1 0 1716 0 1 2815
box -3 -3 3 3
use M3_M2  M3_M2_6389
timestamp 1745462530
transform 1 0 1652 0 1 2525
box -3 -3 3 3
use M3_M2  M3_M2_6390
timestamp 1745462530
transform 1 0 1948 0 1 2755
box -3 -3 3 3
use M3_M2  M3_M2_6391
timestamp 1745462530
transform 1 0 1940 0 1 2635
box -3 -3 3 3
use M3_M2  M3_M2_6392
timestamp 1745462530
transform 1 0 1924 0 1 2635
box -3 -3 3 3
use M3_M2  M3_M2_6393
timestamp 1745462530
transform 1 0 1908 0 1 2755
box -3 -3 3 3
use M3_M2  M3_M2_6394
timestamp 1745462530
transform 1 0 1892 0 1 2925
box -3 -3 3 3
use M3_M2  M3_M2_6395
timestamp 1745462530
transform 1 0 1852 0 1 2925
box -3 -3 3 3
use M3_M2  M3_M2_6396
timestamp 1745462530
transform 1 0 1180 0 1 2475
box -3 -3 3 3
use M3_M2  M3_M2_6397
timestamp 1745462530
transform 1 0 1132 0 1 2475
box -3 -3 3 3
use M3_M2  M3_M2_6398
timestamp 1745462530
transform 1 0 1636 0 1 2835
box -3 -3 3 3
use M3_M2  M3_M2_6399
timestamp 1745462530
transform 1 0 1564 0 1 2835
box -3 -3 3 3
use M3_M2  M3_M2_6400
timestamp 1745462530
transform 1 0 1564 0 1 2525
box -3 -3 3 3
use M3_M2  M3_M2_6401
timestamp 1745462530
transform 1 0 1532 0 1 2525
box -3 -3 3 3
use M3_M2  M3_M2_6402
timestamp 1745462530
transform 1 0 2852 0 1 2905
box -3 -3 3 3
use M3_M2  M3_M2_6403
timestamp 1745462530
transform 1 0 2748 0 1 2905
box -3 -3 3 3
use M3_M2  M3_M2_6404
timestamp 1745462530
transform 1 0 2036 0 1 2925
box -3 -3 3 3
use M3_M2  M3_M2_6405
timestamp 1745462530
transform 1 0 2020 0 1 2915
box -3 -3 3 3
use M3_M2  M3_M2_6406
timestamp 1745462530
transform 1 0 2764 0 1 2715
box -3 -3 3 3
use M3_M2  M3_M2_6407
timestamp 1745462530
transform 1 0 1452 0 1 2765
box -3 -3 3 3
use M3_M2  M3_M2_6408
timestamp 1745462530
transform 1 0 1364 0 1 2765
box -3 -3 3 3
use M3_M2  M3_M2_6409
timestamp 1745462530
transform 1 0 1364 0 1 2715
box -3 -3 3 3
use M3_M2  M3_M2_6410
timestamp 1745462530
transform 1 0 1340 0 1 2715
box -3 -3 3 3
use M3_M2  M3_M2_6411
timestamp 1745462530
transform 1 0 2548 0 1 2695
box -3 -3 3 3
use M3_M2  M3_M2_6412
timestamp 1745462530
transform 1 0 1692 0 1 2695
box -3 -3 3 3
use M3_M2  M3_M2_6413
timestamp 1745462530
transform 1 0 1636 0 1 2695
box -3 -3 3 3
use M3_M2  M3_M2_6414
timestamp 1745462530
transform 1 0 2468 0 1 2835
box -3 -3 3 3
use M3_M2  M3_M2_6415
timestamp 1745462530
transform 1 0 2468 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_6416
timestamp 1745462530
transform 1 0 1964 0 1 2835
box -3 -3 3 3
use M3_M2  M3_M2_6417
timestamp 1745462530
transform 1 0 1948 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_6418
timestamp 1745462530
transform 1 0 2740 0 1 2975
box -3 -3 3 3
use M3_M2  M3_M2_6419
timestamp 1745462530
transform 1 0 2740 0 1 2915
box -3 -3 3 3
use M3_M2  M3_M2_6420
timestamp 1745462530
transform 1 0 2660 0 1 2915
box -3 -3 3 3
use M3_M2  M3_M2_6421
timestamp 1745462530
transform 1 0 1468 0 1 2975
box -3 -3 3 3
use M3_M2  M3_M2_6422
timestamp 1745462530
transform 1 0 1468 0 1 2935
box -3 -3 3 3
use M3_M2  M3_M2_6423
timestamp 1745462530
transform 1 0 1364 0 1 2935
box -3 -3 3 3
use M3_M2  M3_M2_6424
timestamp 1745462530
transform 1 0 1364 0 1 2885
box -3 -3 3 3
use M3_M2  M3_M2_6425
timestamp 1745462530
transform 1 0 1156 0 1 2875
box -3 -3 3 3
use M3_M2  M3_M2_6426
timestamp 1745462530
transform 1 0 2596 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_6427
timestamp 1745462530
transform 1 0 2556 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_6428
timestamp 1745462530
transform 1 0 1516 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_6429
timestamp 1745462530
transform 1 0 1444 0 1 2635
box -3 -3 3 3
use M3_M2  M3_M2_6430
timestamp 1745462530
transform 1 0 1428 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_6431
timestamp 1745462530
transform 1 0 1428 0 1 2635
box -3 -3 3 3
use M3_M2  M3_M2_6432
timestamp 1745462530
transform 1 0 3196 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_6433
timestamp 1745462530
transform 1 0 3092 0 1 2775
box -3 -3 3 3
use M3_M2  M3_M2_6434
timestamp 1745462530
transform 1 0 3028 0 1 2775
box -3 -3 3 3
use M3_M2  M3_M2_6435
timestamp 1745462530
transform 1 0 2996 0 1 2775
box -3 -3 3 3
use M3_M2  M3_M2_6436
timestamp 1745462530
transform 1 0 2956 0 1 2285
box -3 -3 3 3
use M3_M2  M3_M2_6437
timestamp 1745462530
transform 1 0 2956 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_6438
timestamp 1745462530
transform 1 0 2852 0 1 2775
box -3 -3 3 3
use M3_M2  M3_M2_6439
timestamp 1745462530
transform 1 0 2844 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_6440
timestamp 1745462530
transform 1 0 2820 0 1 2285
box -3 -3 3 3
use M3_M2  M3_M2_6441
timestamp 1745462530
transform 1 0 2428 0 1 2275
box -3 -3 3 3
use M3_M2  M3_M2_6442
timestamp 1745462530
transform 1 0 1540 0 1 2385
box -3 -3 3 3
use M3_M2  M3_M2_6443
timestamp 1745462530
transform 1 0 1508 0 1 2385
box -3 -3 3 3
use M3_M2  M3_M2_6444
timestamp 1745462530
transform 1 0 1492 0 1 2785
box -3 -3 3 3
use M3_M2  M3_M2_6445
timestamp 1745462530
transform 1 0 1492 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_6446
timestamp 1745462530
transform 1 0 1476 0 1 3045
box -3 -3 3 3
use M3_M2  M3_M2_6447
timestamp 1745462530
transform 1 0 1476 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_6448
timestamp 1745462530
transform 1 0 1468 0 1 2785
box -3 -3 3 3
use M3_M2  M3_M2_6449
timestamp 1745462530
transform 1 0 1404 0 1 3045
box -3 -3 3 3
use M3_M2  M3_M2_6450
timestamp 1745462530
transform 1 0 1396 0 1 3165
box -3 -3 3 3
use M3_M2  M3_M2_6451
timestamp 1745462530
transform 1 0 1340 0 1 3165
box -3 -3 3 3
use M3_M2  M3_M2_6452
timestamp 1745462530
transform 1 0 1284 0 1 3375
box -3 -3 3 3
use M3_M2  M3_M2_6453
timestamp 1745462530
transform 1 0 956 0 1 1055
box -3 -3 3 3
use M3_M2  M3_M2_6454
timestamp 1745462530
transform 1 0 948 0 1 3375
box -3 -3 3 3
use M3_M2  M3_M2_6455
timestamp 1745462530
transform 1 0 908 0 1 3375
box -3 -3 3 3
use M3_M2  M3_M2_6456
timestamp 1745462530
transform 1 0 748 0 1 1865
box -3 -3 3 3
use M3_M2  M3_M2_6457
timestamp 1745462530
transform 1 0 660 0 1 2065
box -3 -3 3 3
use M3_M2  M3_M2_6458
timestamp 1745462530
transform 1 0 644 0 1 3375
box -3 -3 3 3
use M3_M2  M3_M2_6459
timestamp 1745462530
transform 1 0 644 0 1 3245
box -3 -3 3 3
use M3_M2  M3_M2_6460
timestamp 1745462530
transform 1 0 572 0 1 2065
box -3 -3 3 3
use M3_M2  M3_M2_6461
timestamp 1745462530
transform 1 0 572 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_6462
timestamp 1745462530
transform 1 0 572 0 1 1865
box -3 -3 3 3
use M3_M2  M3_M2_6463
timestamp 1745462530
transform 1 0 556 0 1 2245
box -3 -3 3 3
use M3_M2  M3_M2_6464
timestamp 1745462530
transform 1 0 548 0 1 1865
box -3 -3 3 3
use M3_M2  M3_M2_6465
timestamp 1745462530
transform 1 0 540 0 1 3245
box -3 -3 3 3
use M3_M2  M3_M2_6466
timestamp 1745462530
transform 1 0 516 0 1 1055
box -3 -3 3 3
use M3_M2  M3_M2_6467
timestamp 1745462530
transform 1 0 500 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_6468
timestamp 1745462530
transform 1 0 132 0 1 3245
box -3 -3 3 3
use M3_M2  M3_M2_6469
timestamp 1745462530
transform 1 0 132 0 1 2245
box -3 -3 3 3
use M3_M2  M3_M2_6470
timestamp 1745462530
transform 1 0 1332 0 1 3305
box -3 -3 3 3
use M3_M2  M3_M2_6471
timestamp 1745462530
transform 1 0 1220 0 1 3305
box -3 -3 3 3
use M3_M2  M3_M2_6472
timestamp 1745462530
transform 1 0 1404 0 1 3405
box -3 -3 3 3
use M3_M2  M3_M2_6473
timestamp 1745462530
transform 1 0 1340 0 1 3405
box -3 -3 3 3
use M3_M2  M3_M2_6474
timestamp 1745462530
transform 1 0 1476 0 1 3425
box -3 -3 3 3
use M3_M2  M3_M2_6475
timestamp 1745462530
transform 1 0 1228 0 1 3425
box -3 -3 3 3
use M3_M2  M3_M2_6476
timestamp 1745462530
transform 1 0 1428 0 1 3515
box -3 -3 3 3
use M3_M2  M3_M2_6477
timestamp 1745462530
transform 1 0 1324 0 1 3515
box -3 -3 3 3
use M3_M2  M3_M2_6478
timestamp 1745462530
transform 1 0 1284 0 1 3715
box -3 -3 3 3
use M3_M2  M3_M2_6479
timestamp 1745462530
transform 1 0 1212 0 1 3715
box -3 -3 3 3
use M3_M2  M3_M2_6480
timestamp 1745462530
transform 1 0 1420 0 1 3625
box -3 -3 3 3
use M3_M2  M3_M2_6481
timestamp 1745462530
transform 1 0 1220 0 1 3625
box -3 -3 3 3
use M3_M2  M3_M2_6482
timestamp 1745462530
transform 1 0 2292 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_6483
timestamp 1745462530
transform 1 0 2260 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_6484
timestamp 1745462530
transform 1 0 2252 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_6485
timestamp 1745462530
transform 1 0 1604 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_6486
timestamp 1745462530
transform 1 0 1532 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_6487
timestamp 1745462530
transform 1 0 1124 0 1 3175
box -3 -3 3 3
use M3_M2  M3_M2_6488
timestamp 1745462530
transform 1 0 1068 0 1 3175
box -3 -3 3 3
use M3_M2  M3_M2_6489
timestamp 1745462530
transform 1 0 980 0 1 3385
box -3 -3 3 3
use M3_M2  M3_M2_6490
timestamp 1745462530
transform 1 0 884 0 1 3385
box -3 -3 3 3
use M3_M2  M3_M2_6491
timestamp 1745462530
transform 1 0 228 0 1 3155
box -3 -3 3 3
use M3_M2  M3_M2_6492
timestamp 1745462530
transform 1 0 140 0 1 3155
box -3 -3 3 3
use M3_M2  M3_M2_6493
timestamp 1745462530
transform 1 0 2092 0 1 3065
box -3 -3 3 3
use M3_M2  M3_M2_6494
timestamp 1745462530
transform 1 0 2020 0 1 3065
box -3 -3 3 3
use M3_M2  M3_M2_6495
timestamp 1745462530
transform 1 0 2020 0 1 2945
box -3 -3 3 3
use M3_M2  M3_M2_6496
timestamp 1745462530
transform 1 0 1260 0 1 3035
box -3 -3 3 3
use M3_M2  M3_M2_6497
timestamp 1745462530
transform 1 0 1260 0 1 2945
box -3 -3 3 3
use M3_M2  M3_M2_6498
timestamp 1745462530
transform 1 0 860 0 1 3035
box -3 -3 3 3
use M3_M2  M3_M2_6499
timestamp 1745462530
transform 1 0 2196 0 1 2955
box -3 -3 3 3
use M3_M2  M3_M2_6500
timestamp 1745462530
transform 1 0 708 0 1 2955
box -3 -3 3 3
use M3_M2  M3_M2_6501
timestamp 1745462530
transform 1 0 2188 0 1 3015
box -3 -3 3 3
use M3_M2  M3_M2_6502
timestamp 1745462530
transform 1 0 636 0 1 3025
box -3 -3 3 3
use M3_M2  M3_M2_6503
timestamp 1745462530
transform 1 0 2124 0 1 2985
box -3 -3 3 3
use M3_M2  M3_M2_6504
timestamp 1745462530
transform 1 0 532 0 1 2985
box -3 -3 3 3
use M3_M2  M3_M2_6505
timestamp 1745462530
transform 1 0 2068 0 1 2895
box -3 -3 3 3
use M3_M2  M3_M2_6506
timestamp 1745462530
transform 1 0 1796 0 1 2925
box -3 -3 3 3
use M3_M2  M3_M2_6507
timestamp 1745462530
transform 1 0 1796 0 1 2895
box -3 -3 3 3
use M3_M2  M3_M2_6508
timestamp 1745462530
transform 1 0 788 0 1 3035
box -3 -3 3 3
use M3_M2  M3_M2_6509
timestamp 1745462530
transform 1 0 788 0 1 2925
box -3 -3 3 3
use M3_M2  M3_M2_6510
timestamp 1745462530
transform 1 0 412 0 1 3035
box -3 -3 3 3
use M3_M2  M3_M2_6511
timestamp 1745462530
transform 1 0 2140 0 1 2945
box -3 -3 3 3
use M3_M2  M3_M2_6512
timestamp 1745462530
transform 1 0 2132 0 1 3435
box -3 -3 3 3
use M3_M2  M3_M2_6513
timestamp 1745462530
transform 1 0 2116 0 1 2945
box -3 -3 3 3
use M3_M2  M3_M2_6514
timestamp 1745462530
transform 1 0 292 0 1 3435
box -3 -3 3 3
use M3_M2  M3_M2_6515
timestamp 1745462530
transform 1 0 2404 0 1 2615
box -3 -3 3 3
use M3_M2  M3_M2_6516
timestamp 1745462530
transform 1 0 2356 0 1 2635
box -3 -3 3 3
use M3_M2  M3_M2_6517
timestamp 1745462530
transform 1 0 2356 0 1 2615
box -3 -3 3 3
use M3_M2  M3_M2_6518
timestamp 1745462530
transform 1 0 2268 0 1 2635
box -3 -3 3 3
use M3_M2  M3_M2_6519
timestamp 1745462530
transform 1 0 2140 0 1 2635
box -3 -3 3 3
use M3_M2  M3_M2_6520
timestamp 1745462530
transform 1 0 2532 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_6521
timestamp 1745462530
transform 1 0 2492 0 1 2045
box -3 -3 3 3
use M3_M2  M3_M2_6522
timestamp 1745462530
transform 1 0 2492 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_6523
timestamp 1745462530
transform 1 0 2460 0 1 1575
box -3 -3 3 3
use M3_M2  M3_M2_6524
timestamp 1745462530
transform 1 0 2460 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_6525
timestamp 1745462530
transform 1 0 2420 0 1 2705
box -3 -3 3 3
use M3_M2  M3_M2_6526
timestamp 1745462530
transform 1 0 2420 0 1 2045
box -3 -3 3 3
use M3_M2  M3_M2_6527
timestamp 1745462530
transform 1 0 2420 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_6528
timestamp 1745462530
transform 1 0 2388 0 1 1575
box -3 -3 3 3
use M3_M2  M3_M2_6529
timestamp 1745462530
transform 1 0 2340 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_6530
timestamp 1745462530
transform 1 0 2340 0 1 1575
box -3 -3 3 3
use M3_M2  M3_M2_6531
timestamp 1745462530
transform 1 0 2324 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_6532
timestamp 1745462530
transform 1 0 2324 0 1 1575
box -3 -3 3 3
use M3_M2  M3_M2_6533
timestamp 1745462530
transform 1 0 2316 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_6534
timestamp 1745462530
transform 1 0 2236 0 1 2705
box -3 -3 3 3
use M3_M2  M3_M2_6535
timestamp 1745462530
transform 1 0 2084 0 1 2705
box -3 -3 3 3
use M3_M2  M3_M2_6536
timestamp 1745462530
transform 1 0 2204 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_6537
timestamp 1745462530
transform 1 0 2132 0 1 2665
box -3 -3 3 3
use M3_M2  M3_M2_6538
timestamp 1745462530
transform 1 0 2132 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_6539
timestamp 1745462530
transform 1 0 2060 0 1 2665
box -3 -3 3 3
use M3_M2  M3_M2_6540
timestamp 1745462530
transform 1 0 2180 0 1 1835
box -3 -3 3 3
use M3_M2  M3_M2_6541
timestamp 1745462530
transform 1 0 2164 0 1 2915
box -3 -3 3 3
use M3_M2  M3_M2_6542
timestamp 1745462530
transform 1 0 2164 0 1 1835
box -3 -3 3 3
use M3_M2  M3_M2_6543
timestamp 1745462530
transform 1 0 2108 0 1 2915
box -3 -3 3 3
use M3_M2  M3_M2_6544
timestamp 1745462530
transform 1 0 3548 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_6545
timestamp 1745462530
transform 1 0 3524 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_6546
timestamp 1745462530
transform 1 0 3516 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_6547
timestamp 1745462530
transform 1 0 2780 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_6548
timestamp 1745462530
transform 1 0 2660 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_6549
timestamp 1745462530
transform 1 0 2620 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_6550
timestamp 1745462530
transform 1 0 2620 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_6551
timestamp 1745462530
transform 1 0 2596 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_6552
timestamp 1745462530
transform 1 0 2596 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_6553
timestamp 1745462530
transform 1 0 2580 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_6554
timestamp 1745462530
transform 1 0 2580 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_6555
timestamp 1745462530
transform 1 0 2580 0 1 405
box -3 -3 3 3
use M3_M2  M3_M2_6556
timestamp 1745462530
transform 1 0 2524 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_6557
timestamp 1745462530
transform 1 0 2516 0 1 265
box -3 -3 3 3
use M3_M2  M3_M2_6558
timestamp 1745462530
transform 1 0 2420 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_6559
timestamp 1745462530
transform 1 0 2412 0 1 1655
box -3 -3 3 3
use M3_M2  M3_M2_6560
timestamp 1745462530
transform 1 0 2364 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_6561
timestamp 1745462530
transform 1 0 2364 0 1 1655
box -3 -3 3 3
use M3_M2  M3_M2_6562
timestamp 1745462530
transform 1 0 2300 0 1 3055
box -3 -3 3 3
use M3_M2  M3_M2_6563
timestamp 1745462530
transform 1 0 2300 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_6564
timestamp 1745462530
transform 1 0 2268 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_6565
timestamp 1745462530
transform 1 0 2268 0 1 2565
box -3 -3 3 3
use M3_M2  M3_M2_6566
timestamp 1745462530
transform 1 0 2252 0 1 3055
box -3 -3 3 3
use M3_M2  M3_M2_6567
timestamp 1745462530
transform 1 0 2252 0 1 2565
box -3 -3 3 3
use M3_M2  M3_M2_6568
timestamp 1745462530
transform 1 0 2252 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_6569
timestamp 1745462530
transform 1 0 2228 0 1 3525
box -3 -3 3 3
use M3_M2  M3_M2_6570
timestamp 1745462530
transform 1 0 2228 0 1 3475
box -3 -3 3 3
use M3_M2  M3_M2_6571
timestamp 1745462530
transform 1 0 2212 0 1 3765
box -3 -3 3 3
use M3_M2  M3_M2_6572
timestamp 1745462530
transform 1 0 2196 0 1 3765
box -3 -3 3 3
use M3_M2  M3_M2_6573
timestamp 1745462530
transform 1 0 2196 0 1 3535
box -3 -3 3 3
use M3_M2  M3_M2_6574
timestamp 1745462530
transform 1 0 2196 0 1 3475
box -3 -3 3 3
use M3_M2  M3_M2_6575
timestamp 1745462530
transform 1 0 2196 0 1 3055
box -3 -3 3 3
use M3_M2  M3_M2_6576
timestamp 1745462530
transform 1 0 1972 0 1 265
box -3 -3 3 3
use M3_M2  M3_M2_6577
timestamp 1745462530
transform 1 0 1628 0 1 3055
box -3 -3 3 3
use M3_M2  M3_M2_6578
timestamp 1745462530
transform 1 0 1140 0 1 3765
box -3 -3 3 3
use M3_M2  M3_M2_6579
timestamp 1745462530
transform 1 0 1236 0 1 3245
box -3 -3 3 3
use M3_M2  M3_M2_6580
timestamp 1745462530
transform 1 0 1220 0 1 3485
box -3 -3 3 3
use M3_M2  M3_M2_6581
timestamp 1745462530
transform 1 0 1212 0 1 3245
box -3 -3 3 3
use M3_M2  M3_M2_6582
timestamp 1745462530
transform 1 0 1148 0 1 3585
box -3 -3 3 3
use M3_M2  M3_M2_6583
timestamp 1745462530
transform 1 0 1092 0 1 3585
box -3 -3 3 3
use M3_M2  M3_M2_6584
timestamp 1745462530
transform 1 0 1092 0 1 3485
box -3 -3 3 3
use M3_M2  M3_M2_6585
timestamp 1745462530
transform 1 0 1724 0 1 2965
box -3 -3 3 3
use M3_M2  M3_M2_6586
timestamp 1745462530
transform 1 0 1212 0 1 2965
box -3 -3 3 3
use M3_M2  M3_M2_6587
timestamp 1745462530
transform 1 0 1356 0 1 3045
box -3 -3 3 3
use M3_M2  M3_M2_6588
timestamp 1745462530
transform 1 0 1188 0 1 3045
box -3 -3 3 3
use M3_M2  M3_M2_6589
timestamp 1745462530
transform 1 0 1524 0 1 2125
box -3 -3 3 3
use M3_M2  M3_M2_6590
timestamp 1745462530
transform 1 0 1452 0 1 2125
box -3 -3 3 3
use M3_M2  M3_M2_6591
timestamp 1745462530
transform 1 0 1444 0 1 2735
box -3 -3 3 3
use M3_M2  M3_M2_6592
timestamp 1745462530
transform 1 0 1412 0 1 2735
box -3 -3 3 3
use M3_M2  M3_M2_6593
timestamp 1745462530
transform 1 0 1236 0 1 2185
box -3 -3 3 3
use M3_M2  M3_M2_6594
timestamp 1745462530
transform 1 0 1188 0 1 2185
box -3 -3 3 3
use M3_M2  M3_M2_6595
timestamp 1745462530
transform 1 0 1780 0 1 3085
box -3 -3 3 3
use M3_M2  M3_M2_6596
timestamp 1745462530
transform 1 0 1708 0 1 3085
box -3 -3 3 3
use M3_M2  M3_M2_6597
timestamp 1745462530
transform 1 0 1820 0 1 3035
box -3 -3 3 3
use M3_M2  M3_M2_6598
timestamp 1745462530
transform 1 0 1724 0 1 3035
box -3 -3 3 3
use M3_M2  M3_M2_6599
timestamp 1745462530
transform 1 0 1876 0 1 2965
box -3 -3 3 3
use M3_M2  M3_M2_6600
timestamp 1745462530
transform 1 0 1796 0 1 2965
box -3 -3 3 3
use M3_M2  M3_M2_6601
timestamp 1745462530
transform 1 0 1812 0 1 3075
box -3 -3 3 3
use M3_M2  M3_M2_6602
timestamp 1745462530
transform 1 0 1796 0 1 3075
box -3 -3 3 3
use M3_M2  M3_M2_6603
timestamp 1745462530
transform 1 0 1852 0 1 2525
box -3 -3 3 3
use M3_M2  M3_M2_6604
timestamp 1745462530
transform 1 0 1820 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_6605
timestamp 1745462530
transform 1 0 1684 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_6606
timestamp 1745462530
transform 1 0 1668 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_6607
timestamp 1745462530
transform 1 0 1668 0 1 1525
box -3 -3 3 3
use M3_M2  M3_M2_6608
timestamp 1745462530
transform 1 0 1548 0 1 1525
box -3 -3 3 3
use M3_M2  M3_M2_6609
timestamp 1745462530
transform 1 0 1924 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_6610
timestamp 1745462530
transform 1 0 1836 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_6611
timestamp 1745462530
transform 1 0 1828 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_6612
timestamp 1745462530
transform 1 0 1796 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_6613
timestamp 1745462530
transform 1 0 876 0 1 3215
box -3 -3 3 3
use M3_M2  M3_M2_6614
timestamp 1745462530
transform 1 0 796 0 1 3215
box -3 -3 3 3
use M3_M2  M3_M2_6615
timestamp 1745462530
transform 1 0 996 0 1 3205
box -3 -3 3 3
use M3_M2  M3_M2_6616
timestamp 1745462530
transform 1 0 924 0 1 3205
box -3 -3 3 3
use M3_M2  M3_M2_6617
timestamp 1745462530
transform 1 0 812 0 1 3205
box -3 -3 3 3
use M3_M2  M3_M2_6618
timestamp 1745462530
transform 1 0 940 0 1 3215
box -3 -3 3 3
use M3_M2  M3_M2_6619
timestamp 1745462530
transform 1 0 868 0 1 3225
box -3 -3 3 3
use M3_M2  M3_M2_6620
timestamp 1745462530
transform 1 0 700 0 1 3215
box -3 -3 3 3
use M3_M2  M3_M2_6621
timestamp 1745462530
transform 1 0 668 0 1 3215
box -3 -3 3 3
use M3_M2  M3_M2_6622
timestamp 1745462530
transform 1 0 3140 0 1 3615
box -3 -3 3 3
use M3_M2  M3_M2_6623
timestamp 1745462530
transform 1 0 3116 0 1 3615
box -3 -3 3 3
use M3_M2  M3_M2_6624
timestamp 1745462530
transform 1 0 3092 0 1 3615
box -3 -3 3 3
use M3_M2  M3_M2_6625
timestamp 1745462530
transform 1 0 2996 0 1 3615
box -3 -3 3 3
use M3_M2  M3_M2_6626
timestamp 1745462530
transform 1 0 3412 0 1 3745
box -3 -3 3 3
use M3_M2  M3_M2_6627
timestamp 1745462530
transform 1 0 3348 0 1 3745
box -3 -3 3 3
use M3_M2  M3_M2_6628
timestamp 1745462530
transform 1 0 3132 0 1 3745
box -3 -3 3 3
use M3_M2  M3_M2_6629
timestamp 1745462530
transform 1 0 3116 0 1 3635
box -3 -3 3 3
use M3_M2  M3_M2_6630
timestamp 1745462530
transform 1 0 2980 0 1 3635
box -3 -3 3 3
use M3_M2  M3_M2_6631
timestamp 1745462530
transform 1 0 2972 0 1 3575
box -3 -3 3 3
use M3_M2  M3_M2_6632
timestamp 1745462530
transform 1 0 2780 0 1 3575
box -3 -3 3 3
use M3_M2  M3_M2_6633
timestamp 1745462530
transform 1 0 2308 0 1 3585
box -3 -3 3 3
use M3_M2  M3_M2_6634
timestamp 1745462530
transform 1 0 2140 0 1 3585
box -3 -3 3 3
use M3_M2  M3_M2_6635
timestamp 1745462530
transform 1 0 1732 0 1 3585
box -3 -3 3 3
use M3_M2  M3_M2_6636
timestamp 1745462530
transform 1 0 3060 0 1 3745
box -3 -3 3 3
use M3_M2  M3_M2_6637
timestamp 1745462530
transform 1 0 2996 0 1 3745
box -3 -3 3 3
use M3_M2  M3_M2_6638
timestamp 1745462530
transform 1 0 2988 0 1 3665
box -3 -3 3 3
use M3_M2  M3_M2_6639
timestamp 1745462530
transform 1 0 2988 0 1 3415
box -3 -3 3 3
use M3_M2  M3_M2_6640
timestamp 1745462530
transform 1 0 2972 0 1 3665
box -3 -3 3 3
use M3_M2  M3_M2_6641
timestamp 1745462530
transform 1 0 2916 0 1 3665
box -3 -3 3 3
use M3_M2  M3_M2_6642
timestamp 1745462530
transform 1 0 2036 0 1 3415
box -3 -3 3 3
use M3_M2  M3_M2_6643
timestamp 1745462530
transform 1 0 2036 0 1 3355
box -3 -3 3 3
use M3_M2  M3_M2_6644
timestamp 1745462530
transform 1 0 1948 0 1 3355
box -3 -3 3 3
use M3_M2  M3_M2_6645
timestamp 1745462530
transform 1 0 1844 0 1 3355
box -3 -3 3 3
use M3_M2  M3_M2_6646
timestamp 1745462530
transform 1 0 1692 0 1 3355
box -3 -3 3 3
use M3_M2  M3_M2_6647
timestamp 1745462530
transform 1 0 2204 0 1 3135
box -3 -3 3 3
use M3_M2  M3_M2_6648
timestamp 1745462530
transform 1 0 2108 0 1 3135
box -3 -3 3 3
use M3_M2  M3_M2_6649
timestamp 1745462530
transform 1 0 3308 0 1 3345
box -3 -3 3 3
use M3_M2  M3_M2_6650
timestamp 1745462530
transform 1 0 3268 0 1 3345
box -3 -3 3 3
use M3_M2  M3_M2_6651
timestamp 1745462530
transform 1 0 3260 0 1 3395
box -3 -3 3 3
use M3_M2  M3_M2_6652
timestamp 1745462530
transform 1 0 3228 0 1 3395
box -3 -3 3 3
use M3_M2  M3_M2_6653
timestamp 1745462530
transform 1 0 3156 0 1 3395
box -3 -3 3 3
use M3_M2  M3_M2_6654
timestamp 1745462530
transform 1 0 3068 0 1 3395
box -3 -3 3 3
use M3_M2  M3_M2_6655
timestamp 1745462530
transform 1 0 2836 0 1 3395
box -3 -3 3 3
use M3_M2  M3_M2_6656
timestamp 1745462530
transform 1 0 2388 0 1 3395
box -3 -3 3 3
use M3_M2  M3_M2_6657
timestamp 1745462530
transform 1 0 2356 0 1 3395
box -3 -3 3 3
use M3_M2  M3_M2_6658
timestamp 1745462530
transform 1 0 3076 0 1 3345
box -3 -3 3 3
use M3_M2  M3_M2_6659
timestamp 1745462530
transform 1 0 3052 0 1 3585
box -3 -3 3 3
use M3_M2  M3_M2_6660
timestamp 1745462530
transform 1 0 3020 0 1 3345
box -3 -3 3 3
use M3_M2  M3_M2_6661
timestamp 1745462530
transform 1 0 3004 0 1 3585
box -3 -3 3 3
use M3_M2  M3_M2_6662
timestamp 1745462530
transform 1 0 2972 0 1 3345
box -3 -3 3 3
use M3_M2  M3_M2_6663
timestamp 1745462530
transform 1 0 2932 0 1 3345
box -3 -3 3 3
use M3_M2  M3_M2_6664
timestamp 1745462530
transform 1 0 2924 0 1 3585
box -3 -3 3 3
use M3_M2  M3_M2_6665
timestamp 1745462530
transform 1 0 2828 0 1 3335
box -3 -3 3 3
use M3_M2  M3_M2_6666
timestamp 1745462530
transform 1 0 3100 0 1 3415
box -3 -3 3 3
use M3_M2  M3_M2_6667
timestamp 1745462530
transform 1 0 3060 0 1 3415
box -3 -3 3 3
use M3_M2  M3_M2_6668
timestamp 1745462530
transform 1 0 2004 0 1 3165
box -3 -3 3 3
use M3_M2  M3_M2_6669
timestamp 1745462530
transform 1 0 1948 0 1 3165
box -3 -3 3 3
use M3_M2  M3_M2_6670
timestamp 1745462530
transform 1 0 3220 0 1 3415
box -3 -3 3 3
use M3_M2  M3_M2_6671
timestamp 1745462530
transform 1 0 3180 0 1 3415
box -3 -3 3 3
use M3_M2  M3_M2_6672
timestamp 1745462530
transform 1 0 3140 0 1 3415
box -3 -3 3 3
use M3_M2  M3_M2_6673
timestamp 1745462530
transform 1 0 3140 0 1 3385
box -3 -3 3 3
use M3_M2  M3_M2_6674
timestamp 1745462530
transform 1 0 3060 0 1 3385
box -3 -3 3 3
use M3_M2  M3_M2_6675
timestamp 1745462530
transform 1 0 2892 0 1 3385
box -3 -3 3 3
use M3_M2  M3_M2_6676
timestamp 1745462530
transform 1 0 2692 0 1 3665
box -3 -3 3 3
use M3_M2  M3_M2_6677
timestamp 1745462530
transform 1 0 2668 0 1 3665
box -3 -3 3 3
use M3_M2  M3_M2_6678
timestamp 1745462530
transform 1 0 2668 0 1 3385
box -3 -3 3 3
use M3_M2  M3_M2_6679
timestamp 1745462530
transform 1 0 2660 0 1 3345
box -3 -3 3 3
use M3_M2  M3_M2_6680
timestamp 1745462530
transform 1 0 2612 0 1 3345
box -3 -3 3 3
use M3_M2  M3_M2_6681
timestamp 1745462530
transform 1 0 3404 0 1 3955
box -3 -3 3 3
use M3_M2  M3_M2_6682
timestamp 1745462530
transform 1 0 3372 0 1 3955
box -3 -3 3 3
use M3_M2  M3_M2_6683
timestamp 1745462530
transform 1 0 3436 0 1 3715
box -3 -3 3 3
use M3_M2  M3_M2_6684
timestamp 1745462530
transform 1 0 3412 0 1 3715
box -3 -3 3 3
use M3_M2  M3_M2_6685
timestamp 1745462530
transform 1 0 3884 0 1 3295
box -3 -3 3 3
use M3_M2  M3_M2_6686
timestamp 1745462530
transform 1 0 3868 0 1 3585
box -3 -3 3 3
use M3_M2  M3_M2_6687
timestamp 1745462530
transform 1 0 3812 0 1 3695
box -3 -3 3 3
use M3_M2  M3_M2_6688
timestamp 1745462530
transform 1 0 3804 0 1 3585
box -3 -3 3 3
use M3_M2  M3_M2_6689
timestamp 1745462530
transform 1 0 3764 0 1 3295
box -3 -3 3 3
use M3_M2  M3_M2_6690
timestamp 1745462530
transform 1 0 3724 0 1 3585
box -3 -3 3 3
use M3_M2  M3_M2_6691
timestamp 1745462530
transform 1 0 3596 0 1 3585
box -3 -3 3 3
use M3_M2  M3_M2_6692
timestamp 1745462530
transform 1 0 3420 0 1 3695
box -3 -3 3 3
use M3_M2  M3_M2_6693
timestamp 1745462530
transform 1 0 3284 0 1 3735
box -3 -3 3 3
use M3_M2  M3_M2_6694
timestamp 1745462530
transform 1 0 3284 0 1 3695
box -3 -3 3 3
use M3_M2  M3_M2_6695
timestamp 1745462530
transform 1 0 3220 0 1 3735
box -3 -3 3 3
use M3_M2  M3_M2_6696
timestamp 1745462530
transform 1 0 1796 0 1 3735
box -3 -3 3 3
use M3_M2  M3_M2_6697
timestamp 1745462530
transform 1 0 3668 0 1 3315
box -3 -3 3 3
use M3_M2  M3_M2_6698
timestamp 1745462530
transform 1 0 3604 0 1 3335
box -3 -3 3 3
use M3_M2  M3_M2_6699
timestamp 1745462530
transform 1 0 3596 0 1 3315
box -3 -3 3 3
use M3_M2  M3_M2_6700
timestamp 1745462530
transform 1 0 3492 0 1 3405
box -3 -3 3 3
use M3_M2  M3_M2_6701
timestamp 1745462530
transform 1 0 3492 0 1 3335
box -3 -3 3 3
use M3_M2  M3_M2_6702
timestamp 1745462530
transform 1 0 3436 0 1 3415
box -3 -3 3 3
use M3_M2  M3_M2_6703
timestamp 1745462530
transform 1 0 3412 0 1 3565
box -3 -3 3 3
use M3_M2  M3_M2_6704
timestamp 1745462530
transform 1 0 3300 0 1 3565
box -3 -3 3 3
use M3_M2  M3_M2_6705
timestamp 1745462530
transform 1 0 3292 0 1 3335
box -3 -3 3 3
use M3_M2  M3_M2_6706
timestamp 1745462530
transform 1 0 3180 0 1 3335
box -3 -3 3 3
use M3_M2  M3_M2_6707
timestamp 1745462530
transform 1 0 3324 0 1 3315
box -3 -3 3 3
use M3_M2  M3_M2_6708
timestamp 1745462530
transform 1 0 3188 0 1 3315
box -3 -3 3 3
use M3_M2  M3_M2_6709
timestamp 1745462530
transform 1 0 2372 0 1 3095
box -3 -3 3 3
use M3_M2  M3_M2_6710
timestamp 1745462530
transform 1 0 2012 0 1 3095
box -3 -3 3 3
use M3_M2  M3_M2_6711
timestamp 1745462530
transform 1 0 3340 0 1 3935
box -3 -3 3 3
use M3_M2  M3_M2_6712
timestamp 1745462530
transform 1 0 3284 0 1 3935
box -3 -3 3 3
use M3_M2  M3_M2_6713
timestamp 1745462530
transform 1 0 3268 0 1 3645
box -3 -3 3 3
use M3_M2  M3_M2_6714
timestamp 1745462530
transform 1 0 3268 0 1 3525
box -3 -3 3 3
use M3_M2  M3_M2_6715
timestamp 1745462530
transform 1 0 3244 0 1 3525
box -3 -3 3 3
use M3_M2  M3_M2_6716
timestamp 1745462530
transform 1 0 3236 0 1 3645
box -3 -3 3 3
use M3_M2  M3_M2_6717
timestamp 1745462530
transform 1 0 3372 0 1 3755
box -3 -3 3 3
use M3_M2  M3_M2_6718
timestamp 1745462530
transform 1 0 3284 0 1 3755
box -3 -3 3 3
use M3_M2  M3_M2_6719
timestamp 1745462530
transform 1 0 3820 0 1 3325
box -3 -3 3 3
use M3_M2  M3_M2_6720
timestamp 1745462530
transform 1 0 3764 0 1 3495
box -3 -3 3 3
use M3_M2  M3_M2_6721
timestamp 1745462530
transform 1 0 3740 0 1 3325
box -3 -3 3 3
use M3_M2  M3_M2_6722
timestamp 1745462530
transform 1 0 3732 0 1 3355
box -3 -3 3 3
use M3_M2  M3_M2_6723
timestamp 1745462530
transform 1 0 3708 0 1 3745
box -3 -3 3 3
use M3_M2  M3_M2_6724
timestamp 1745462530
transform 1 0 3652 0 1 3355
box -3 -3 3 3
use M3_M2  M3_M2_6725
timestamp 1745462530
transform 1 0 3644 0 1 3745
box -3 -3 3 3
use M3_M2  M3_M2_6726
timestamp 1745462530
transform 1 0 3644 0 1 3715
box -3 -3 3 3
use M3_M2  M3_M2_6727
timestamp 1745462530
transform 1 0 3644 0 1 3495
box -3 -3 3 3
use M3_M2  M3_M2_6728
timestamp 1745462530
transform 1 0 3436 0 1 3705
box -3 -3 3 3
use M3_M2  M3_M2_6729
timestamp 1745462530
transform 1 0 3356 0 1 3775
box -3 -3 3 3
use M3_M2  M3_M2_6730
timestamp 1745462530
transform 1 0 3356 0 1 3705
box -3 -3 3 3
use M3_M2  M3_M2_6731
timestamp 1745462530
transform 1 0 3196 0 1 3775
box -3 -3 3 3
use M3_M2  M3_M2_6732
timestamp 1745462530
transform 1 0 3188 0 1 3915
box -3 -3 3 3
use M3_M2  M3_M2_6733
timestamp 1745462530
transform 1 0 2092 0 1 3915
box -3 -3 3 3
use M3_M2  M3_M2_6734
timestamp 1745462530
transform 1 0 2052 0 1 3625
box -3 -3 3 3
use M3_M2  M3_M2_6735
timestamp 1745462530
transform 1 0 1940 0 1 3625
box -3 -3 3 3
use M3_M2  M3_M2_6736
timestamp 1745462530
transform 1 0 1940 0 1 3495
box -3 -3 3 3
use M3_M2  M3_M2_6737
timestamp 1745462530
transform 1 0 1892 0 1 3495
box -3 -3 3 3
use M3_M2  M3_M2_6738
timestamp 1745462530
transform 1 0 1892 0 1 3335
box -3 -3 3 3
use M3_M2  M3_M2_6739
timestamp 1745462530
transform 1 0 1748 0 1 3335
box -3 -3 3 3
use M3_M2  M3_M2_6740
timestamp 1745462530
transform 1 0 3716 0 1 3565
box -3 -3 3 3
use M3_M2  M3_M2_6741
timestamp 1745462530
transform 1 0 3676 0 1 3245
box -3 -3 3 3
use M3_M2  M3_M2_6742
timestamp 1745462530
transform 1 0 3660 0 1 3625
box -3 -3 3 3
use M3_M2  M3_M2_6743
timestamp 1745462530
transform 1 0 3660 0 1 3565
box -3 -3 3 3
use M3_M2  M3_M2_6744
timestamp 1745462530
transform 1 0 3572 0 1 3245
box -3 -3 3 3
use M3_M2  M3_M2_6745
timestamp 1745462530
transform 1 0 3436 0 1 3365
box -3 -3 3 3
use M3_M2  M3_M2_6746
timestamp 1745462530
transform 1 0 3436 0 1 3245
box -3 -3 3 3
use M3_M2  M3_M2_6747
timestamp 1745462530
transform 1 0 3388 0 1 3615
box -3 -3 3 3
use M3_M2  M3_M2_6748
timestamp 1745462530
transform 1 0 3292 0 1 3615
box -3 -3 3 3
use M3_M2  M3_M2_6749
timestamp 1745462530
transform 1 0 3236 0 1 3385
box -3 -3 3 3
use M3_M2  M3_M2_6750
timestamp 1745462530
transform 1 0 3236 0 1 3365
box -3 -3 3 3
use M3_M2  M3_M2_6751
timestamp 1745462530
transform 1 0 3156 0 1 3385
box -3 -3 3 3
use M3_M2  M3_M2_6752
timestamp 1745462530
transform 1 0 3252 0 1 3405
box -3 -3 3 3
use M3_M2  M3_M2_6753
timestamp 1745462530
transform 1 0 3212 0 1 3405
box -3 -3 3 3
use M3_M2  M3_M2_6754
timestamp 1745462530
transform 1 0 3388 0 1 3645
box -3 -3 3 3
use M3_M2  M3_M2_6755
timestamp 1745462530
transform 1 0 3340 0 1 3645
box -3 -3 3 3
use M3_M2  M3_M2_6756
timestamp 1745462530
transform 1 0 3324 0 1 3405
box -3 -3 3 3
use M3_M2  M3_M2_6757
timestamp 1745462530
transform 1 0 3300 0 1 3405
box -3 -3 3 3
use M3_M2  M3_M2_6758
timestamp 1745462530
transform 1 0 3860 0 1 3565
box -3 -3 3 3
use M3_M2  M3_M2_6759
timestamp 1745462530
transform 1 0 3828 0 1 3225
box -3 -3 3 3
use M3_M2  M3_M2_6760
timestamp 1745462530
transform 1 0 3756 0 1 3605
box -3 -3 3 3
use M3_M2  M3_M2_6761
timestamp 1745462530
transform 1 0 3756 0 1 3565
box -3 -3 3 3
use M3_M2  M3_M2_6762
timestamp 1745462530
transform 1 0 3740 0 1 3565
box -3 -3 3 3
use M3_M2  M3_M2_6763
timestamp 1745462530
transform 1 0 3628 0 1 3225
box -3 -3 3 3
use M3_M2  M3_M2_6764
timestamp 1745462530
transform 1 0 3524 0 1 3605
box -3 -3 3 3
use M3_M2  M3_M2_6765
timestamp 1745462530
transform 1 0 3356 0 1 3625
box -3 -3 3 3
use M3_M2  M3_M2_6766
timestamp 1745462530
transform 1 0 3356 0 1 3605
box -3 -3 3 3
use M3_M2  M3_M2_6767
timestamp 1745462530
transform 1 0 3164 0 1 3605
box -3 -3 3 3
use M3_M2  M3_M2_6768
timestamp 1745462530
transform 1 0 1876 0 1 3595
box -3 -3 3 3
use M3_M2  M3_M2_6769
timestamp 1745462530
transform 1 0 1876 0 1 3495
box -3 -3 3 3
use M3_M2  M3_M2_6770
timestamp 1745462530
transform 1 0 1724 0 1 3495
box -3 -3 3 3
use M3_M2  M3_M2_6771
timestamp 1745462530
transform 1 0 3556 0 1 3345
box -3 -3 3 3
use M3_M2  M3_M2_6772
timestamp 1745462530
transform 1 0 3540 0 1 3035
box -3 -3 3 3
use M3_M2  M3_M2_6773
timestamp 1745462530
transform 1 0 3532 0 1 3345
box -3 -3 3 3
use M3_M2  M3_M2_6774
timestamp 1745462530
transform 1 0 3532 0 1 3285
box -3 -3 3 3
use M3_M2  M3_M2_6775
timestamp 1745462530
transform 1 0 3396 0 1 3285
box -3 -3 3 3
use M3_M2  M3_M2_6776
timestamp 1745462530
transform 1 0 3316 0 1 3395
box -3 -3 3 3
use M3_M2  M3_M2_6777
timestamp 1745462530
transform 1 0 3276 0 1 3395
box -3 -3 3 3
use M3_M2  M3_M2_6778
timestamp 1745462530
transform 1 0 3276 0 1 3285
box -3 -3 3 3
use M3_M2  M3_M2_6779
timestamp 1745462530
transform 1 0 3116 0 1 3035
box -3 -3 3 3
use M3_M2  M3_M2_6780
timestamp 1745462530
transform 1 0 3292 0 1 3295
box -3 -3 3 3
use M3_M2  M3_M2_6781
timestamp 1745462530
transform 1 0 3236 0 1 3295
box -3 -3 3 3
use M3_M2  M3_M2_6782
timestamp 1745462530
transform 1 0 3196 0 1 3955
box -3 -3 3 3
use M3_M2  M3_M2_6783
timestamp 1745462530
transform 1 0 3164 0 1 3955
box -3 -3 3 3
use M3_M2  M3_M2_6784
timestamp 1745462530
transform 1 0 3164 0 1 3635
box -3 -3 3 3
use M3_M2  M3_M2_6785
timestamp 1745462530
transform 1 0 3132 0 1 3635
box -3 -3 3 3
use M3_M2  M3_M2_6786
timestamp 1745462530
transform 1 0 3780 0 1 3385
box -3 -3 3 3
use M3_M2  M3_M2_6787
timestamp 1745462530
transform 1 0 3772 0 1 3655
box -3 -3 3 3
use M3_M2  M3_M2_6788
timestamp 1745462530
transform 1 0 3740 0 1 3385
box -3 -3 3 3
use M3_M2  M3_M2_6789
timestamp 1745462530
transform 1 0 3660 0 1 3675
box -3 -3 3 3
use M3_M2  M3_M2_6790
timestamp 1745462530
transform 1 0 3660 0 1 3655
box -3 -3 3 3
use M3_M2  M3_M2_6791
timestamp 1745462530
transform 1 0 3556 0 1 3675
box -3 -3 3 3
use M3_M2  M3_M2_6792
timestamp 1745462530
transform 1 0 3540 0 1 3715
box -3 -3 3 3
use M3_M2  M3_M2_6793
timestamp 1745462530
transform 1 0 3332 0 1 3785
box -3 -3 3 3
use M3_M2  M3_M2_6794
timestamp 1745462530
transform 1 0 3332 0 1 3725
box -3 -3 3 3
use M3_M2  M3_M2_6795
timestamp 1745462530
transform 1 0 3156 0 1 3755
box -3 -3 3 3
use M3_M2  M3_M2_6796
timestamp 1745462530
transform 1 0 3108 0 1 3875
box -3 -3 3 3
use M3_M2  M3_M2_6797
timestamp 1745462530
transform 1 0 3108 0 1 3795
box -3 -3 3 3
use M3_M2  M3_M2_6798
timestamp 1745462530
transform 1 0 3108 0 1 3755
box -3 -3 3 3
use M3_M2  M3_M2_6799
timestamp 1745462530
transform 1 0 1652 0 1 3875
box -3 -3 3 3
use M3_M2  M3_M2_6800
timestamp 1745462530
transform 1 0 1652 0 1 3355
box -3 -3 3 3
use M3_M2  M3_M2_6801
timestamp 1745462530
transform 1 0 1636 0 1 3635
box -3 -3 3 3
use M3_M2  M3_M2_6802
timestamp 1745462530
transform 1 0 1572 0 1 3355
box -3 -3 3 3
use M3_M2  M3_M2_6803
timestamp 1745462530
transform 1 0 1564 0 1 3635
box -3 -3 3 3
use M3_M2  M3_M2_6804
timestamp 1745462530
transform 1 0 3580 0 1 3255
box -3 -3 3 3
use M3_M2  M3_M2_6805
timestamp 1745462530
transform 1 0 3524 0 1 3255
box -3 -3 3 3
use M3_M2  M3_M2_6806
timestamp 1745462530
transform 1 0 3220 0 1 3275
box -3 -3 3 3
use M3_M2  M3_M2_6807
timestamp 1745462530
transform 1 0 3212 0 1 3545
box -3 -3 3 3
use M3_M2  M3_M2_6808
timestamp 1745462530
transform 1 0 3172 0 1 3295
box -3 -3 3 3
use M3_M2  M3_M2_6809
timestamp 1745462530
transform 1 0 3148 0 1 3545
box -3 -3 3 3
use M3_M2  M3_M2_6810
timestamp 1745462530
transform 1 0 3092 0 1 3295
box -3 -3 3 3
use M3_M2  M3_M2_6811
timestamp 1745462530
transform 1 0 3180 0 1 3345
box -3 -3 3 3
use M3_M2  M3_M2_6812
timestamp 1745462530
transform 1 0 3132 0 1 3345
box -3 -3 3 3
use M3_M2  M3_M2_6813
timestamp 1745462530
transform 1 0 2044 0 1 3135
box -3 -3 3 3
use M3_M2  M3_M2_6814
timestamp 1745462530
transform 1 0 1932 0 1 3135
box -3 -3 3 3
use M3_M2  M3_M2_6815
timestamp 1745462530
transform 1 0 2428 0 1 3935
box -3 -3 3 3
use M3_M2  M3_M2_6816
timestamp 1745462530
transform 1 0 2388 0 1 3935
box -3 -3 3 3
use M3_M2  M3_M2_6817
timestamp 1745462530
transform 1 0 2420 0 1 3475
box -3 -3 3 3
use M3_M2  M3_M2_6818
timestamp 1745462530
transform 1 0 2364 0 1 3475
box -3 -3 3 3
use M3_M2  M3_M2_6819
timestamp 1745462530
transform 1 0 2460 0 1 3665
box -3 -3 3 3
use M3_M2  M3_M2_6820
timestamp 1745462530
transform 1 0 2412 0 1 3695
box -3 -3 3 3
use M3_M2  M3_M2_6821
timestamp 1745462530
transform 1 0 2412 0 1 3665
box -3 -3 3 3
use M3_M2  M3_M2_6822
timestamp 1745462530
transform 1 0 2356 0 1 3695
box -3 -3 3 3
use M3_M2  M3_M2_6823
timestamp 1745462530
transform 1 0 2356 0 1 3665
box -3 -3 3 3
use M3_M2  M3_M2_6824
timestamp 1745462530
transform 1 0 2356 0 1 3625
box -3 -3 3 3
use M3_M2  M3_M2_6825
timestamp 1745462530
transform 1 0 2340 0 1 3625
box -3 -3 3 3
use M3_M2  M3_M2_6826
timestamp 1745462530
transform 1 0 2108 0 1 3665
box -3 -3 3 3
use M3_M2  M3_M2_6827
timestamp 1745462530
transform 1 0 2108 0 1 3465
box -3 -3 3 3
use M3_M2  M3_M2_6828
timestamp 1745462530
transform 1 0 2108 0 1 3195
box -3 -3 3 3
use M3_M2  M3_M2_6829
timestamp 1745462530
transform 1 0 1980 0 1 3495
box -3 -3 3 3
use M3_M2  M3_M2_6830
timestamp 1745462530
transform 1 0 1980 0 1 3465
box -3 -3 3 3
use M3_M2  M3_M2_6831
timestamp 1745462530
transform 1 0 1964 0 1 3195
box -3 -3 3 3
use M3_M2  M3_M2_6832
timestamp 1745462530
transform 1 0 1908 0 1 3515
box -3 -3 3 3
use M3_M2  M3_M2_6833
timestamp 1745462530
transform 1 0 1884 0 1 3195
box -3 -3 3 3
use M3_M2  M3_M2_6834
timestamp 1745462530
transform 1 0 1796 0 1 3205
box -3 -3 3 3
use M3_M2  M3_M2_6835
timestamp 1745462530
transform 1 0 1796 0 1 3155
box -3 -3 3 3
use M3_M2  M3_M2_6836
timestamp 1745462530
transform 1 0 1684 0 1 3155
box -3 -3 3 3
use M3_M2  M3_M2_6837
timestamp 1745462530
transform 1 0 2956 0 1 3265
box -3 -3 3 3
use M3_M2  M3_M2_6838
timestamp 1745462530
transform 1 0 2588 0 1 3635
box -3 -3 3 3
use M3_M2  M3_M2_6839
timestamp 1745462530
transform 1 0 2500 0 1 3635
box -3 -3 3 3
use M3_M2  M3_M2_6840
timestamp 1745462530
transform 1 0 2500 0 1 3615
box -3 -3 3 3
use M3_M2  M3_M2_6841
timestamp 1745462530
transform 1 0 2460 0 1 3265
box -3 -3 3 3
use M3_M2  M3_M2_6842
timestamp 1745462530
transform 1 0 2436 0 1 3265
box -3 -3 3 3
use M3_M2  M3_M2_6843
timestamp 1745462530
transform 1 0 2412 0 1 3615
box -3 -3 3 3
use M3_M2  M3_M2_6844
timestamp 1745462530
transform 1 0 2404 0 1 3265
box -3 -3 3 3
use M3_M2  M3_M2_6845
timestamp 1745462530
transform 1 0 2364 0 1 3265
box -3 -3 3 3
use M3_M2  M3_M2_6846
timestamp 1745462530
transform 1 0 2644 0 1 3375
box -3 -3 3 3
use M3_M2  M3_M2_6847
timestamp 1745462530
transform 1 0 2428 0 1 3375
box -3 -3 3 3
use M3_M2  M3_M2_6848
timestamp 1745462530
transform 1 0 2260 0 1 3225
box -3 -3 3 3
use M3_M2  M3_M2_6849
timestamp 1745462530
transform 1 0 1980 0 1 3225
box -3 -3 3 3
use M3_M2  M3_M2_6850
timestamp 1745462530
transform 1 0 2148 0 1 3905
box -3 -3 3 3
use M3_M2  M3_M2_6851
timestamp 1745462530
transform 1 0 2108 0 1 3955
box -3 -3 3 3
use M3_M2  M3_M2_6852
timestamp 1745462530
transform 1 0 2076 0 1 3955
box -3 -3 3 3
use M3_M2  M3_M2_6853
timestamp 1745462530
transform 1 0 2076 0 1 3905
box -3 -3 3 3
use M3_M2  M3_M2_6854
timestamp 1745462530
transform 1 0 2380 0 1 3565
box -3 -3 3 3
use M3_M2  M3_M2_6855
timestamp 1745462530
transform 1 0 2100 0 1 3565
box -3 -3 3 3
use M3_M2  M3_M2_6856
timestamp 1745462530
transform 1 0 2260 0 1 3765
box -3 -3 3 3
use M3_M2  M3_M2_6857
timestamp 1745462530
transform 1 0 2260 0 1 3655
box -3 -3 3 3
use M3_M2  M3_M2_6858
timestamp 1745462530
transform 1 0 2236 0 1 3655
box -3 -3 3 3
use M3_M2  M3_M2_6859
timestamp 1745462530
transform 1 0 2236 0 1 3605
box -3 -3 3 3
use M3_M2  M3_M2_6860
timestamp 1745462530
transform 1 0 2228 0 1 3765
box -3 -3 3 3
use M3_M2  M3_M2_6861
timestamp 1745462530
transform 1 0 2180 0 1 3475
box -3 -3 3 3
use M3_M2  M3_M2_6862
timestamp 1745462530
transform 1 0 2148 0 1 3605
box -3 -3 3 3
use M3_M2  M3_M2_6863
timestamp 1745462530
transform 1 0 2148 0 1 3515
box -3 -3 3 3
use M3_M2  M3_M2_6864
timestamp 1745462530
transform 1 0 2148 0 1 3475
box -3 -3 3 3
use M3_M2  M3_M2_6865
timestamp 1745462530
transform 1 0 1996 0 1 3515
box -3 -3 3 3
use M3_M2  M3_M2_6866
timestamp 1745462530
transform 1 0 1996 0 1 3415
box -3 -3 3 3
use M3_M2  M3_M2_6867
timestamp 1745462530
transform 1 0 1884 0 1 3415
box -3 -3 3 3
use M3_M2  M3_M2_6868
timestamp 1745462530
transform 1 0 1852 0 1 3415
box -3 -3 3 3
use M3_M2  M3_M2_6869
timestamp 1745462530
transform 1 0 1852 0 1 3295
box -3 -3 3 3
use M3_M2  M3_M2_6870
timestamp 1745462530
transform 1 0 1804 0 1 3295
box -3 -3 3 3
use M3_M2  M3_M2_6871
timestamp 1745462530
transform 1 0 1692 0 1 3415
box -3 -3 3 3
use M3_M2  M3_M2_6872
timestamp 1745462530
transform 1 0 2364 0 1 3455
box -3 -3 3 3
use M3_M2  M3_M2_6873
timestamp 1745462530
transform 1 0 2316 0 1 3475
box -3 -3 3 3
use M3_M2  M3_M2_6874
timestamp 1745462530
transform 1 0 2316 0 1 3455
box -3 -3 3 3
use M3_M2  M3_M2_6875
timestamp 1745462530
transform 1 0 2316 0 1 3085
box -3 -3 3 3
use M3_M2  M3_M2_6876
timestamp 1745462530
transform 1 0 2284 0 1 3475
box -3 -3 3 3
use M3_M2  M3_M2_6877
timestamp 1745462530
transform 1 0 2276 0 1 3555
box -3 -3 3 3
use M3_M2  M3_M2_6878
timestamp 1745462530
transform 1 0 2276 0 1 3085
box -3 -3 3 3
use M3_M2  M3_M2_6879
timestamp 1745462530
transform 1 0 2236 0 1 3555
box -3 -3 3 3
use M3_M2  M3_M2_6880
timestamp 1745462530
transform 1 0 2604 0 1 3455
box -3 -3 3 3
use M3_M2  M3_M2_6881
timestamp 1745462530
transform 1 0 2380 0 1 3455
box -3 -3 3 3
use M3_M2  M3_M2_6882
timestamp 1745462530
transform 1 0 2876 0 1 3955
box -3 -3 3 3
use M3_M2  M3_M2_6883
timestamp 1745462530
transform 1 0 2844 0 1 3955
box -3 -3 3 3
use M3_M2  M3_M2_6884
timestamp 1745462530
transform 1 0 3604 0 1 3685
box -3 -3 3 3
use M3_M2  M3_M2_6885
timestamp 1745462530
transform 1 0 3532 0 1 3685
box -3 -3 3 3
use M3_M2  M3_M2_6886
timestamp 1745462530
transform 1 0 3428 0 1 3685
box -3 -3 3 3
use M3_M2  M3_M2_6887
timestamp 1745462530
transform 1 0 3124 0 1 3685
box -3 -3 3 3
use M3_M2  M3_M2_6888
timestamp 1745462530
transform 1 0 3052 0 1 3685
box -3 -3 3 3
use M3_M2  M3_M2_6889
timestamp 1745462530
transform 1 0 2828 0 1 3715
box -3 -3 3 3
use M3_M2  M3_M2_6890
timestamp 1745462530
transform 1 0 2820 0 1 3685
box -3 -3 3 3
use M3_M2  M3_M2_6891
timestamp 1745462530
transform 1 0 2636 0 1 3725
box -3 -3 3 3
use M3_M2  M3_M2_6892
timestamp 1745462530
transform 1 0 2636 0 1 3655
box -3 -3 3 3
use M3_M2  M3_M2_6893
timestamp 1745462530
transform 1 0 2492 0 1 3655
box -3 -3 3 3
use M3_M2  M3_M2_6894
timestamp 1745462530
transform 1 0 2468 0 1 3715
box -3 -3 3 3
use M3_M2  M3_M2_6895
timestamp 1745462530
transform 1 0 2404 0 1 3715
box -3 -3 3 3
use M3_M2  M3_M2_6896
timestamp 1745462530
transform 1 0 2276 0 1 3715
box -3 -3 3 3
use M3_M2  M3_M2_6897
timestamp 1745462530
transform 1 0 1900 0 1 3575
box -3 -3 3 3
use M3_M2  M3_M2_6898
timestamp 1745462530
transform 1 0 1868 0 1 3715
box -3 -3 3 3
use M3_M2  M3_M2_6899
timestamp 1745462530
transform 1 0 1860 0 1 3575
box -3 -3 3 3
use M3_M2  M3_M2_6900
timestamp 1745462530
transform 1 0 2836 0 1 3635
box -3 -3 3 3
use M3_M2  M3_M2_6901
timestamp 1745462530
transform 1 0 2764 0 1 3635
box -3 -3 3 3
use M3_M2  M3_M2_6902
timestamp 1745462530
transform 1 0 2764 0 1 3405
box -3 -3 3 3
use M3_M2  M3_M2_6903
timestamp 1745462530
transform 1 0 2724 0 1 3635
box -3 -3 3 3
use M3_M2  M3_M2_6904
timestamp 1745462530
transform 1 0 2604 0 1 3405
box -3 -3 3 3
use M3_M2  M3_M2_6905
timestamp 1745462530
transform 1 0 2580 0 1 3465
box -3 -3 3 3
use M3_M2  M3_M2_6906
timestamp 1745462530
transform 1 0 2580 0 1 3405
box -3 -3 3 3
use M3_M2  M3_M2_6907
timestamp 1745462530
transform 1 0 2172 0 1 3465
box -3 -3 3 3
use M3_M2  M3_M2_6908
timestamp 1745462530
transform 1 0 2172 0 1 3255
box -3 -3 3 3
use M3_M2  M3_M2_6909
timestamp 1745462530
transform 1 0 1956 0 1 3245
box -3 -3 3 3
use M3_M2  M3_M2_6910
timestamp 1745462530
transform 1 0 1756 0 1 3245
box -3 -3 3 3
use M3_M2  M3_M2_6911
timestamp 1745462530
transform 1 0 3428 0 1 3515
box -3 -3 3 3
use M3_M2  M3_M2_6912
timestamp 1745462530
transform 1 0 3396 0 1 3515
box -3 -3 3 3
use M3_M2  M3_M2_6913
timestamp 1745462530
transform 1 0 3148 0 1 3515
box -3 -3 3 3
use M3_M2  M3_M2_6914
timestamp 1745462530
transform 1 0 3060 0 1 3515
box -3 -3 3 3
use M3_M2  M3_M2_6915
timestamp 1745462530
transform 1 0 2844 0 1 3515
box -3 -3 3 3
use M3_M2  M3_M2_6916
timestamp 1745462530
transform 1 0 2500 0 1 3515
box -3 -3 3 3
use M3_M2  M3_M2_6917
timestamp 1745462530
transform 1 0 2316 0 1 3515
box -3 -3 3 3
use M3_M2  M3_M2_6918
timestamp 1745462530
transform 1 0 3020 0 1 3285
box -3 -3 3 3
use M3_M2  M3_M2_6919
timestamp 1745462530
transform 1 0 2836 0 1 3495
box -3 -3 3 3
use M3_M2  M3_M2_6920
timestamp 1745462530
transform 1 0 2836 0 1 3285
box -3 -3 3 3
use M3_M2  M3_M2_6921
timestamp 1745462530
transform 1 0 2740 0 1 3505
box -3 -3 3 3
use M3_M2  M3_M2_6922
timestamp 1745462530
transform 1 0 2708 0 1 3245
box -3 -3 3 3
use M3_M2  M3_M2_6923
timestamp 1745462530
transform 1 0 2684 0 1 3505
box -3 -3 3 3
use M3_M2  M3_M2_6924
timestamp 1745462530
transform 1 0 2652 0 1 3505
box -3 -3 3 3
use M3_M2  M3_M2_6925
timestamp 1745462530
transform 1 0 2636 0 1 3245
box -3 -3 3 3
use M3_M2  M3_M2_6926
timestamp 1745462530
transform 1 0 3412 0 1 3495
box -3 -3 3 3
use M3_M2  M3_M2_6927
timestamp 1745462530
transform 1 0 3388 0 1 3495
box -3 -3 3 3
use M3_M2  M3_M2_6928
timestamp 1745462530
transform 1 0 3364 0 1 3495
box -3 -3 3 3
use M3_M2  M3_M2_6929
timestamp 1745462530
transform 1 0 3132 0 1 3505
box -3 -3 3 3
use M3_M2  M3_M2_6930
timestamp 1745462530
transform 1 0 3084 0 1 3505
box -3 -3 3 3
use M3_M2  M3_M2_6931
timestamp 1745462530
transform 1 0 2908 0 1 3505
box -3 -3 3 3
use M3_M2  M3_M2_6932
timestamp 1745462530
transform 1 0 2884 0 1 3605
box -3 -3 3 3
use M3_M2  M3_M2_6933
timestamp 1745462530
transform 1 0 2580 0 1 3615
box -3 -3 3 3
use M3_M2  M3_M2_6934
timestamp 1745462530
transform 1 0 2532 0 1 3485
box -3 -3 3 3
use M3_M2  M3_M2_6935
timestamp 1745462530
transform 1 0 2484 0 1 3485
box -3 -3 3 3
use M3_M2  M3_M2_6936
timestamp 1745462530
transform 1 0 3628 0 1 3575
box -3 -3 3 3
use M3_M2  M3_M2_6937
timestamp 1745462530
transform 1 0 3460 0 1 3575
box -3 -3 3 3
use M3_M2  M3_M2_6938
timestamp 1745462530
transform 1 0 3444 0 1 3505
box -3 -3 3 3
use M3_M2  M3_M2_6939
timestamp 1745462530
transform 1 0 3348 0 1 3505
box -3 -3 3 3
use M3_M2  M3_M2_6940
timestamp 1745462530
transform 1 0 3644 0 1 3895
box -3 -3 3 3
use M3_M2  M3_M2_6941
timestamp 1745462530
transform 1 0 3588 0 1 3895
box -3 -3 3 3
use M3_M2  M3_M2_6942
timestamp 1745462530
transform 1 0 3500 0 1 3895
box -3 -3 3 3
use M3_M2  M3_M2_6943
timestamp 1745462530
transform 1 0 3628 0 1 3745
box -3 -3 3 3
use M3_M2  M3_M2_6944
timestamp 1745462530
transform 1 0 3596 0 1 3745
box -3 -3 3 3
use M3_M2  M3_M2_6945
timestamp 1745462530
transform 1 0 3596 0 1 3615
box -3 -3 3 3
use M3_M2  M3_M2_6946
timestamp 1745462530
transform 1 0 3508 0 1 3615
box -3 -3 3 3
use M3_M2  M3_M2_6947
timestamp 1745462530
transform 1 0 3452 0 1 3465
box -3 -3 3 3
use M3_M2  M3_M2_6948
timestamp 1745462530
transform 1 0 3412 0 1 3465
box -3 -3 3 3
use M3_M2  M3_M2_6949
timestamp 1745462530
transform 1 0 3532 0 1 3725
box -3 -3 3 3
use M3_M2  M3_M2_6950
timestamp 1745462530
transform 1 0 3516 0 1 3725
box -3 -3 3 3
use M3_M2  M3_M2_6951
timestamp 1745462530
transform 1 0 3420 0 1 3415
box -3 -3 3 3
use M3_M2  M3_M2_6952
timestamp 1745462530
transform 1 0 3380 0 1 3415
box -3 -3 3 3
use M3_M2  M3_M2_6953
timestamp 1745462530
transform 1 0 3268 0 1 4085
box -3 -3 3 3
use M3_M2  M3_M2_6954
timestamp 1745462530
transform 1 0 3252 0 1 3875
box -3 -3 3 3
use M3_M2  M3_M2_6955
timestamp 1745462530
transform 1 0 3236 0 1 4085
box -3 -3 3 3
use M3_M2  M3_M2_6956
timestamp 1745462530
transform 1 0 3196 0 1 3875
box -3 -3 3 3
use M3_M2  M3_M2_6957
timestamp 1745462530
transform 1 0 3196 0 1 3575
box -3 -3 3 3
use M3_M2  M3_M2_6958
timestamp 1745462530
transform 1 0 3164 0 1 3575
box -3 -3 3 3
use M3_M2  M3_M2_6959
timestamp 1745462530
transform 1 0 3204 0 1 3785
box -3 -3 3 3
use M3_M2  M3_M2_6960
timestamp 1745462530
transform 1 0 3148 0 1 3785
box -3 -3 3 3
use M3_M2  M3_M2_6961
timestamp 1745462530
transform 1 0 3172 0 1 3585
box -3 -3 3 3
use M3_M2  M3_M2_6962
timestamp 1745462530
transform 1 0 3116 0 1 3585
box -3 -3 3 3
use M3_M2  M3_M2_6963
timestamp 1745462530
transform 1 0 2540 0 1 3695
box -3 -3 3 3
use M3_M2  M3_M2_6964
timestamp 1745462530
transform 1 0 2444 0 1 3695
box -3 -3 3 3
use M3_M2  M3_M2_6965
timestamp 1745462530
transform 1 0 2532 0 1 3545
box -3 -3 3 3
use M3_M2  M3_M2_6966
timestamp 1745462530
transform 1 0 2508 0 1 3545
box -3 -3 3 3
use M3_M2  M3_M2_6967
timestamp 1745462530
transform 1 0 2348 0 1 3885
box -3 -3 3 3
use M3_M2  M3_M2_6968
timestamp 1745462530
transform 1 0 2252 0 1 3895
box -3 -3 3 3
use M3_M2  M3_M2_6969
timestamp 1745462530
transform 1 0 2212 0 1 3895
box -3 -3 3 3
use M3_M2  M3_M2_6970
timestamp 1745462530
transform 1 0 2452 0 1 3495
box -3 -3 3 3
use M3_M2  M3_M2_6971
timestamp 1745462530
transform 1 0 2372 0 1 3495
box -3 -3 3 3
use M3_M2  M3_M2_6972
timestamp 1745462530
transform 1 0 2116 0 1 3745
box -3 -3 3 3
use M3_M2  M3_M2_6973
timestamp 1745462530
transform 1 0 1900 0 1 3745
box -3 -3 3 3
use M3_M2  M3_M2_6974
timestamp 1745462530
transform 1 0 2652 0 1 3675
box -3 -3 3 3
use M3_M2  M3_M2_6975
timestamp 1745462530
transform 1 0 2628 0 1 3675
box -3 -3 3 3
use M3_M2  M3_M2_6976
timestamp 1745462530
transform 1 0 2588 0 1 3675
box -3 -3 3 3
use M3_M2  M3_M2_6977
timestamp 1745462530
transform 1 0 2548 0 1 3675
box -3 -3 3 3
use M3_M2  M3_M2_6978
timestamp 1745462530
transform 1 0 2396 0 1 3675
box -3 -3 3 3
use M3_M2  M3_M2_6979
timestamp 1745462530
transform 1 0 1884 0 1 3675
box -3 -3 3 3
use M3_M2  M3_M2_6980
timestamp 1745462530
transform 1 0 1780 0 1 3675
box -3 -3 3 3
use M3_M2  M3_M2_6981
timestamp 1745462530
transform 1 0 1780 0 1 3595
box -3 -3 3 3
use M3_M2  M3_M2_6982
timestamp 1745462530
transform 1 0 1628 0 1 3595
box -3 -3 3 3
use M3_M2  M3_M2_6983
timestamp 1745462530
transform 1 0 2724 0 1 2965
box -3 -3 3 3
use M3_M2  M3_M2_6984
timestamp 1745462530
transform 1 0 2716 0 1 2565
box -3 -3 3 3
use M3_M2  M3_M2_6985
timestamp 1745462530
transform 1 0 2652 0 1 2565
box -3 -3 3 3
use M3_M2  M3_M2_6986
timestamp 1745462530
transform 1 0 2644 0 1 2285
box -3 -3 3 3
use M3_M2  M3_M2_6987
timestamp 1745462530
transform 1 0 2580 0 1 2965
box -3 -3 3 3
use M3_M2  M3_M2_6988
timestamp 1745462530
transform 1 0 2476 0 1 2965
box -3 -3 3 3
use M3_M2  M3_M2_6989
timestamp 1745462530
transform 1 0 2476 0 1 2285
box -3 -3 3 3
use M3_M2  M3_M2_6990
timestamp 1745462530
transform 1 0 2468 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_6991
timestamp 1745462530
transform 1 0 2412 0 1 2965
box -3 -3 3 3
use M3_M2  M3_M2_6992
timestamp 1745462530
transform 1 0 2412 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_6993
timestamp 1745462530
transform 1 0 2540 0 1 3025
box -3 -3 3 3
use M3_M2  M3_M2_6994
timestamp 1745462530
transform 1 0 2508 0 1 3025
box -3 -3 3 3
use M3_M2  M3_M2_6995
timestamp 1745462530
transform 1 0 2484 0 1 3025
box -3 -3 3 3
use M3_M2  M3_M2_6996
timestamp 1745462530
transform 1 0 2420 0 1 3025
box -3 -3 3 3
use M3_M2  M3_M2_6997
timestamp 1745462530
transform 1 0 2396 0 1 2565
box -3 -3 3 3
use M3_M2  M3_M2_6998
timestamp 1745462530
transform 1 0 2380 0 1 2565
box -3 -3 3 3
use M3_M2  M3_M2_6999
timestamp 1745462530
transform 1 0 2372 0 1 3025
box -3 -3 3 3
use M3_M2  M3_M2_7000
timestamp 1745462530
transform 1 0 2612 0 1 3015
box -3 -3 3 3
use M3_M2  M3_M2_7001
timestamp 1745462530
transform 1 0 2572 0 1 3015
box -3 -3 3 3
use M3_M2  M3_M2_7002
timestamp 1745462530
transform 1 0 2428 0 1 3015
box -3 -3 3 3
use M3_M2  M3_M2_7003
timestamp 1745462530
transform 1 0 2364 0 1 3015
box -3 -3 3 3
use M3_M2  M3_M2_7004
timestamp 1745462530
transform 1 0 2356 0 1 1865
box -3 -3 3 3
use M3_M2  M3_M2_7005
timestamp 1745462530
transform 1 0 2284 0 1 1865
box -3 -3 3 3
use M3_M2  M3_M2_7006
timestamp 1745462530
transform 1 0 2260 0 1 3365
box -3 -3 3 3
use M3_M2  M3_M2_7007
timestamp 1745462530
transform 1 0 2140 0 1 3365
box -3 -3 3 3
use M3_M2  M3_M2_7008
timestamp 1745462530
transform 1 0 2748 0 1 3945
box -3 -3 3 3
use M3_M2  M3_M2_7009
timestamp 1745462530
transform 1 0 2732 0 1 3945
box -3 -3 3 3
use M3_M2  M3_M2_7010
timestamp 1745462530
transform 1 0 2772 0 1 3565
box -3 -3 3 3
use M3_M2  M3_M2_7011
timestamp 1745462530
transform 1 0 2748 0 1 3565
box -3 -3 3 3
use M3_M2  M3_M2_7012
timestamp 1745462530
transform 1 0 2788 0 1 3625
box -3 -3 3 3
use M3_M2  M3_M2_7013
timestamp 1745462530
transform 1 0 2772 0 1 3625
box -3 -3 3 3
use M3_M2  M3_M2_7014
timestamp 1745462530
transform 1 0 3236 0 1 3695
box -3 -3 3 3
use M3_M2  M3_M2_7015
timestamp 1745462530
transform 1 0 3180 0 1 3695
box -3 -3 3 3
use M3_M2  M3_M2_7016
timestamp 1745462530
transform 1 0 3156 0 1 3695
box -3 -3 3 3
use M3_M2  M3_M2_7017
timestamp 1745462530
transform 1 0 2996 0 1 3695
box -3 -3 3 3
use M3_M2  M3_M2_7018
timestamp 1745462530
transform 1 0 2780 0 1 3685
box -3 -3 3 3
use M3_M2  M3_M2_7019
timestamp 1745462530
transform 1 0 2364 0 1 3685
box -3 -3 3 3
use M3_M2  M3_M2_7020
timestamp 1745462530
transform 1 0 2228 0 1 3685
box -3 -3 3 3
use M3_M2  M3_M2_7021
timestamp 1745462530
transform 1 0 2116 0 1 3685
box -3 -3 3 3
use M3_M2  M3_M2_7022
timestamp 1745462530
transform 1 0 2116 0 1 3615
box -3 -3 3 3
use M3_M2  M3_M2_7023
timestamp 1745462530
transform 1 0 1852 0 1 3615
box -3 -3 3 3
use M3_M2  M3_M2_7024
timestamp 1745462530
transform 1 0 3308 0 1 3505
box -3 -3 3 3
use M3_M2  M3_M2_7025
timestamp 1745462530
transform 1 0 3292 0 1 3575
box -3 -3 3 3
use M3_M2  M3_M2_7026
timestamp 1745462530
transform 1 0 3220 0 1 3585
box -3 -3 3 3
use M3_M2  M3_M2_7027
timestamp 1745462530
transform 1 0 3220 0 1 3505
box -3 -3 3 3
use M3_M2  M3_M2_7028
timestamp 1745462530
transform 1 0 3188 0 1 3615
box -3 -3 3 3
use M3_M2  M3_M2_7029
timestamp 1745462530
transform 1 0 3188 0 1 3585
box -3 -3 3 3
use M3_M2  M3_M2_7030
timestamp 1745462530
transform 1 0 3004 0 1 3625
box -3 -3 3 3
use M3_M2  M3_M2_7031
timestamp 1745462530
transform 1 0 2908 0 1 3625
box -3 -3 3 3
use M3_M2  M3_M2_7032
timestamp 1745462530
transform 1 0 2908 0 1 3585
box -3 -3 3 3
use M3_M2  M3_M2_7033
timestamp 1745462530
transform 1 0 2756 0 1 3585
box -3 -3 3 3
use M3_M2  M3_M2_7034
timestamp 1745462530
transform 1 0 2404 0 1 3585
box -3 -3 3 3
use M3_M2  M3_M2_7035
timestamp 1745462530
transform 1 0 2372 0 1 3535
box -3 -3 3 3
use M3_M2  M3_M2_7036
timestamp 1745462530
transform 1 0 2244 0 1 3535
box -3 -3 3 3
use M3_M2  M3_M2_7037
timestamp 1745462530
transform 1 0 3284 0 1 3565
box -3 -3 3 3
use M3_M2  M3_M2_7038
timestamp 1745462530
transform 1 0 3284 0 1 3415
box -3 -3 3 3
use M3_M2  M3_M2_7039
timestamp 1745462530
transform 1 0 3244 0 1 3415
box -3 -3 3 3
use M3_M2  M3_M2_7040
timestamp 1745462530
transform 1 0 3036 0 1 3565
box -3 -3 3 3
use M3_M2  M3_M2_7041
timestamp 1745462530
transform 1 0 2828 0 1 3565
box -3 -3 3 3
use M3_M2  M3_M2_7042
timestamp 1745462530
transform 1 0 2828 0 1 3555
box -3 -3 3 3
use M3_M2  M3_M2_7043
timestamp 1745462530
transform 1 0 2644 0 1 3555
box -3 -3 3 3
use M3_M2  M3_M2_7044
timestamp 1745462530
transform 1 0 2628 0 1 3665
box -3 -3 3 3
use M3_M2  M3_M2_7045
timestamp 1745462530
transform 1 0 2564 0 1 3665
box -3 -3 3 3
use M3_M2  M3_M2_7046
timestamp 1745462530
transform 1 0 2500 0 1 3665
box -3 -3 3 3
use M3_M2  M3_M2_7047
timestamp 1745462530
transform 1 0 2492 0 1 3545
box -3 -3 3 3
use M3_M2  M3_M2_7048
timestamp 1745462530
transform 1 0 2428 0 1 3545
box -3 -3 3 3
use M3_M2  M3_M2_7049
timestamp 1745462530
transform 1 0 3060 0 1 4135
box -3 -3 3 3
use M3_M2  M3_M2_7050
timestamp 1745462530
transform 1 0 3060 0 1 3985
box -3 -3 3 3
use M3_M2  M3_M2_7051
timestamp 1745462530
transform 1 0 3020 0 1 4135
box -3 -3 3 3
use M3_M2  M3_M2_7052
timestamp 1745462530
transform 1 0 3020 0 1 3985
box -3 -3 3 3
use M3_M2  M3_M2_7053
timestamp 1745462530
transform 1 0 3492 0 1 4105
box -3 -3 3 3
use M3_M2  M3_M2_7054
timestamp 1745462530
transform 1 0 3492 0 1 3955
box -3 -3 3 3
use M3_M2  M3_M2_7055
timestamp 1745462530
transform 1 0 3468 0 1 4105
box -3 -3 3 3
use M3_M2  M3_M2_7056
timestamp 1745462530
transform 1 0 3428 0 1 3955
box -3 -3 3 3
use M3_M2  M3_M2_7057
timestamp 1745462530
transform 1 0 3428 0 1 3785
box -3 -3 3 3
use M3_M2  M3_M2_7058
timestamp 1745462530
transform 1 0 3348 0 1 3785
box -3 -3 3 3
use M3_M2  M3_M2_7059
timestamp 1745462530
transform 1 0 3332 0 1 3575
box -3 -3 3 3
use M3_M2  M3_M2_7060
timestamp 1745462530
transform 1 0 3308 0 1 3575
box -3 -3 3 3
use M3_M2  M3_M2_7061
timestamp 1745462530
transform 1 0 3340 0 1 3705
box -3 -3 3 3
use M3_M2  M3_M2_7062
timestamp 1745462530
transform 1 0 3260 0 1 3695
box -3 -3 3 3
use M3_M2  M3_M2_7063
timestamp 1745462530
transform 1 0 3324 0 1 3525
box -3 -3 3 3
use M3_M2  M3_M2_7064
timestamp 1745462530
transform 1 0 3284 0 1 3525
box -3 -3 3 3
use M3_M2  M3_M2_7065
timestamp 1745462530
transform 1 0 3388 0 1 4145
box -3 -3 3 3
use M3_M2  M3_M2_7066
timestamp 1745462530
transform 1 0 3364 0 1 4145
box -3 -3 3 3
use M3_M2  M3_M2_7067
timestamp 1745462530
transform 1 0 3324 0 1 3645
box -3 -3 3 3
use M3_M2  M3_M2_7068
timestamp 1745462530
transform 1 0 3292 0 1 3645
box -3 -3 3 3
use M3_M2  M3_M2_7069
timestamp 1745462530
transform 1 0 3308 0 1 3715
box -3 -3 3 3
use M3_M2  M3_M2_7070
timestamp 1745462530
transform 1 0 3228 0 1 3715
box -3 -3 3 3
use M3_M2  M3_M2_7071
timestamp 1745462530
transform 1 0 3316 0 1 3605
box -3 -3 3 3
use M3_M2  M3_M2_7072
timestamp 1745462530
transform 1 0 3268 0 1 3605
box -3 -3 3 3
use M3_M2  M3_M2_7073
timestamp 1745462530
transform 1 0 3508 0 1 3975
box -3 -3 3 3
use M3_M2  M3_M2_7074
timestamp 1745462530
transform 1 0 3476 0 1 3975
box -3 -3 3 3
use M3_M2  M3_M2_7075
timestamp 1745462530
transform 1 0 3292 0 1 3785
box -3 -3 3 3
use M3_M2  M3_M2_7076
timestamp 1745462530
transform 1 0 3284 0 1 3975
box -3 -3 3 3
use M3_M2  M3_M2_7077
timestamp 1745462530
transform 1 0 3220 0 1 3785
box -3 -3 3 3
use M3_M2  M3_M2_7078
timestamp 1745462530
transform 1 0 3332 0 1 3475
box -3 -3 3 3
use M3_M2  M3_M2_7079
timestamp 1745462530
transform 1 0 3252 0 1 3575
box -3 -3 3 3
use M3_M2  M3_M2_7080
timestamp 1745462530
transform 1 0 3252 0 1 3475
box -3 -3 3 3
use M3_M2  M3_M2_7081
timestamp 1745462530
transform 1 0 3212 0 1 3575
box -3 -3 3 3
use M3_M2  M3_M2_7082
timestamp 1745462530
transform 1 0 3224 0 1 3615
box -3 -3 3 3
use M3_M2  M3_M2_7083
timestamp 1745462530
transform 1 0 3204 0 1 3615
box -3 -3 3 3
use M3_M2  M3_M2_7084
timestamp 1745462530
transform 1 0 3340 0 1 3415
box -3 -3 3 3
use M3_M2  M3_M2_7085
timestamp 1745462530
transform 1 0 3300 0 1 3415
box -3 -3 3 3
use M3_M2  M3_M2_7086
timestamp 1745462530
transform 1 0 3228 0 1 3825
box -3 -3 3 3
use M3_M2  M3_M2_7087
timestamp 1745462530
transform 1 0 3188 0 1 3755
box -3 -3 3 3
use M3_M2  M3_M2_7088
timestamp 1745462530
transform 1 0 3172 0 1 3825
box -3 -3 3 3
use M3_M2  M3_M2_7089
timestamp 1745462530
transform 1 0 3172 0 1 3755
box -3 -3 3 3
use M3_M2  M3_M2_7090
timestamp 1745462530
transform 1 0 3236 0 1 3475
box -3 -3 3 3
use M3_M2  M3_M2_7091
timestamp 1745462530
transform 1 0 3196 0 1 3475
box -3 -3 3 3
use M3_M2  M3_M2_7092
timestamp 1745462530
transform 1 0 2444 0 1 3795
box -3 -3 3 3
use M3_M2  M3_M2_7093
timestamp 1745462530
transform 1 0 2412 0 1 3795
box -3 -3 3 3
use M3_M2  M3_M2_7094
timestamp 1745462530
transform 1 0 2268 0 1 3695
box -3 -3 3 3
use M3_M2  M3_M2_7095
timestamp 1745462530
transform 1 0 2188 0 1 3695
box -3 -3 3 3
use M3_M2  M3_M2_7096
timestamp 1745462530
transform 1 0 1812 0 1 3425
box -3 -3 3 3
use M3_M2  M3_M2_7097
timestamp 1745462530
transform 1 0 1804 0 1 3625
box -3 -3 3 3
use M3_M2  M3_M2_7098
timestamp 1745462530
transform 1 0 1748 0 1 3625
box -3 -3 3 3
use M3_M2  M3_M2_7099
timestamp 1745462530
transform 1 0 1740 0 1 3425
box -3 -3 3 3
use M3_M2  M3_M2_7100
timestamp 1745462530
transform 1 0 2396 0 1 3525
box -3 -3 3 3
use M3_M2  M3_M2_7101
timestamp 1745462530
transform 1 0 2276 0 1 3525
box -3 -3 3 3
use M3_M2  M3_M2_7102
timestamp 1745462530
transform 1 0 2140 0 1 3725
box -3 -3 3 3
use M3_M2  M3_M2_7103
timestamp 1745462530
transform 1 0 1812 0 1 3725
box -3 -3 3 3
use M3_M2  M3_M2_7104
timestamp 1745462530
transform 1 0 2180 0 1 3355
box -3 -3 3 3
use M3_M2  M3_M2_7105
timestamp 1745462530
transform 1 0 2172 0 1 3525
box -3 -3 3 3
use M3_M2  M3_M2_7106
timestamp 1745462530
transform 1 0 2156 0 1 3355
box -3 -3 3 3
use M3_M2  M3_M2_7107
timestamp 1745462530
transform 1 0 2140 0 1 3355
box -3 -3 3 3
use M3_M2  M3_M2_7108
timestamp 1745462530
transform 1 0 2124 0 1 3355
box -3 -3 3 3
use M3_M2  M3_M2_7109
timestamp 1745462530
transform 1 0 2108 0 1 3365
box -3 -3 3 3
use M3_M2  M3_M2_7110
timestamp 1745462530
transform 1 0 2092 0 1 3525
box -3 -3 3 3
use M3_M2  M3_M2_7111
timestamp 1745462530
transform 1 0 2044 0 1 3365
box -3 -3 3 3
use M3_M2  M3_M2_7112
timestamp 1745462530
transform 1 0 1844 0 1 3525
box -3 -3 3 3
use M3_M2  M3_M2_7113
timestamp 1745462530
transform 1 0 1836 0 1 3575
box -3 -3 3 3
use M3_M2  M3_M2_7114
timestamp 1745462530
transform 1 0 1764 0 1 3565
box -3 -3 3 3
use M3_M2  M3_M2_7115
timestamp 1745462530
transform 1 0 1716 0 1 3335
box -3 -3 3 3
use M3_M2  M3_M2_7116
timestamp 1745462530
transform 1 0 1708 0 1 3495
box -3 -3 3 3
use M3_M2  M3_M2_7117
timestamp 1745462530
transform 1 0 1692 0 1 3565
box -3 -3 3 3
use M3_M2  M3_M2_7118
timestamp 1745462530
transform 1 0 1692 0 1 3495
box -3 -3 3 3
use M3_M2  M3_M2_7119
timestamp 1745462530
transform 1 0 1116 0 1 3335
box -3 -3 3 3
use M3_M2  M3_M2_7120
timestamp 1745462530
transform 1 0 2708 0 1 4115
box -3 -3 3 3
use M3_M2  M3_M2_7121
timestamp 1745462530
transform 1 0 2652 0 1 4115
box -3 -3 3 3
use M3_M2  M3_M2_7122
timestamp 1745462530
transform 1 0 2764 0 1 3765
box -3 -3 3 3
use M3_M2  M3_M2_7123
timestamp 1745462530
transform 1 0 2740 0 1 3765
box -3 -3 3 3
use M3_M2  M3_M2_7124
timestamp 1745462530
transform 1 0 3724 0 1 3735
box -3 -3 3 3
use M3_M2  M3_M2_7125
timestamp 1745462530
transform 1 0 3668 0 1 3735
box -3 -3 3 3
use M3_M2  M3_M2_7126
timestamp 1745462530
transform 1 0 2940 0 1 3725
box -3 -3 3 3
use M3_M2  M3_M2_7127
timestamp 1745462530
transform 1 0 2932 0 1 3745
box -3 -3 3 3
use M3_M2  M3_M2_7128
timestamp 1745462530
transform 1 0 2748 0 1 3745
box -3 -3 3 3
use M3_M2  M3_M2_7129
timestamp 1745462530
transform 1 0 2476 0 1 3725
box -3 -3 3 3
use M3_M2  M3_M2_7130
timestamp 1745462530
transform 1 0 2468 0 1 3745
box -3 -3 3 3
use M3_M2  M3_M2_7131
timestamp 1745462530
transform 1 0 2420 0 1 3725
box -3 -3 3 3
use M3_M2  M3_M2_7132
timestamp 1745462530
transform 1 0 2420 0 1 3635
box -3 -3 3 3
use M3_M2  M3_M2_7133
timestamp 1745462530
transform 1 0 2260 0 1 3635
box -3 -3 3 3
use M3_M2  M3_M2_7134
timestamp 1745462530
transform 1 0 1756 0 1 3635
box -3 -3 3 3
use M3_M2  M3_M2_7135
timestamp 1745462530
transform 1 0 3668 0 1 3665
box -3 -3 3 3
use M3_M2  M3_M2_7136
timestamp 1745462530
transform 1 0 3612 0 1 3665
box -3 -3 3 3
use M3_M2  M3_M2_7137
timestamp 1745462530
transform 1 0 3068 0 1 3775
box -3 -3 3 3
use M3_M2  M3_M2_7138
timestamp 1745462530
transform 1 0 3068 0 1 3665
box -3 -3 3 3
use M3_M2  M3_M2_7139
timestamp 1745462530
transform 1 0 2940 0 1 3555
box -3 -3 3 3
use M3_M2  M3_M2_7140
timestamp 1745462530
transform 1 0 2852 0 1 3885
box -3 -3 3 3
use M3_M2  M3_M2_7141
timestamp 1745462530
transform 1 0 2852 0 1 3775
box -3 -3 3 3
use M3_M2  M3_M2_7142
timestamp 1745462530
transform 1 0 2844 0 1 3555
box -3 -3 3 3
use M3_M2  M3_M2_7143
timestamp 1745462530
transform 1 0 2636 0 1 3565
box -3 -3 3 3
use M3_M2  M3_M2_7144
timestamp 1745462530
transform 1 0 2596 0 1 3565
box -3 -3 3 3
use M3_M2  M3_M2_7145
timestamp 1745462530
transform 1 0 2572 0 1 3765
box -3 -3 3 3
use M3_M2  M3_M2_7146
timestamp 1745462530
transform 1 0 2372 0 1 3885
box -3 -3 3 3
use M3_M2  M3_M2_7147
timestamp 1745462530
transform 1 0 2372 0 1 3765
box -3 -3 3 3
use M3_M2  M3_M2_7148
timestamp 1745462530
transform 1 0 2292 0 1 3765
box -3 -3 3 3
use M3_M2  M3_M2_7149
timestamp 1745462530
transform 1 0 2292 0 1 3515
box -3 -3 3 3
use M3_M2  M3_M2_7150
timestamp 1745462530
transform 1 0 2180 0 1 3515
box -3 -3 3 3
use M3_M2  M3_M2_7151
timestamp 1745462530
transform 1 0 2708 0 1 3495
box -3 -3 3 3
use M3_M2  M3_M2_7152
timestamp 1745462530
transform 1 0 2692 0 1 3495
box -3 -3 3 3
use M3_M2  M3_M2_7153
timestamp 1745462530
transform 1 0 3580 0 1 3485
box -3 -3 3 3
use M3_M2  M3_M2_7154
timestamp 1745462530
transform 1 0 3532 0 1 3485
box -3 -3 3 3
use M3_M2  M3_M2_7155
timestamp 1745462530
transform 1 0 3492 0 1 3485
box -3 -3 3 3
use M3_M2  M3_M2_7156
timestamp 1745462530
transform 1 0 2996 0 1 3475
box -3 -3 3 3
use M3_M2  M3_M2_7157
timestamp 1745462530
transform 1 0 2724 0 1 3475
box -3 -3 3 3
use M3_M2  M3_M2_7158
timestamp 1745462530
transform 1 0 2644 0 1 3475
box -3 -3 3 3
use M3_M2  M3_M2_7159
timestamp 1745462530
transform 1 0 2636 0 1 3505
box -3 -3 3 3
use M3_M2  M3_M2_7160
timestamp 1745462530
transform 1 0 2580 0 1 3505
box -3 -3 3 3
use M3_M2  M3_M2_7161
timestamp 1745462530
transform 1 0 2980 0 1 3745
box -3 -3 3 3
use M3_M2  M3_M2_7162
timestamp 1745462530
transform 1 0 2956 0 1 3755
box -3 -3 3 3
use M3_M2  M3_M2_7163
timestamp 1745462530
transform 1 0 3764 0 1 4005
box -3 -3 3 3
use M3_M2  M3_M2_7164
timestamp 1745462530
transform 1 0 3748 0 1 4005
box -3 -3 3 3
use M3_M2  M3_M2_7165
timestamp 1745462530
transform 1 0 3748 0 1 3595
box -3 -3 3 3
use M3_M2  M3_M2_7166
timestamp 1745462530
transform 1 0 3716 0 1 3595
box -3 -3 3 3
use M3_M2  M3_M2_7167
timestamp 1745462530
transform 1 0 3700 0 1 3525
box -3 -3 3 3
use M3_M2  M3_M2_7168
timestamp 1745462530
transform 1 0 3572 0 1 3525
box -3 -3 3 3
use M3_M2  M3_M2_7169
timestamp 1745462530
transform 1 0 3892 0 1 3965
box -3 -3 3 3
use M3_M2  M3_M2_7170
timestamp 1745462530
transform 1 0 3796 0 1 3965
box -3 -3 3 3
use M3_M2  M3_M2_7171
timestamp 1745462530
transform 1 0 3748 0 1 3675
box -3 -3 3 3
use M3_M2  M3_M2_7172
timestamp 1745462530
transform 1 0 3700 0 1 3675
box -3 -3 3 3
use M3_M2  M3_M2_7173
timestamp 1745462530
transform 1 0 3684 0 1 3635
box -3 -3 3 3
use M3_M2  M3_M2_7174
timestamp 1745462530
transform 1 0 3572 0 1 3635
box -3 -3 3 3
use M3_M2  M3_M2_7175
timestamp 1745462530
transform 1 0 3788 0 1 3835
box -3 -3 3 3
use M3_M2  M3_M2_7176
timestamp 1745462530
transform 1 0 3788 0 1 3575
box -3 -3 3 3
use M3_M2  M3_M2_7177
timestamp 1745462530
transform 1 0 3724 0 1 3575
box -3 -3 3 3
use M3_M2  M3_M2_7178
timestamp 1745462530
transform 1 0 3684 0 1 3835
box -3 -3 3 3
use M3_M2  M3_M2_7179
timestamp 1745462530
transform 1 0 3708 0 1 3535
box -3 -3 3 3
use M3_M2  M3_M2_7180
timestamp 1745462530
transform 1 0 3628 0 1 3545
box -3 -3 3 3
use M3_M2  M3_M2_7181
timestamp 1745462530
transform 1 0 3772 0 1 3545
box -3 -3 3 3
use M3_M2  M3_M2_7182
timestamp 1745462530
transform 1 0 3732 0 1 3545
box -3 -3 3 3
use M3_M2  M3_M2_7183
timestamp 1745462530
transform 1 0 3620 0 1 3505
box -3 -3 3 3
use M3_M2  M3_M2_7184
timestamp 1745462530
transform 1 0 3516 0 1 3505
box -3 -3 3 3
use M3_M2  M3_M2_7185
timestamp 1745462530
transform 1 0 3652 0 1 3515
box -3 -3 3 3
use M3_M2  M3_M2_7186
timestamp 1745462530
transform 1 0 3476 0 1 3515
box -3 -3 3 3
use M3_M2  M3_M2_7187
timestamp 1745462530
transform 1 0 2516 0 1 3795
box -3 -3 3 3
use M3_M2  M3_M2_7188
timestamp 1745462530
transform 1 0 2508 0 1 3865
box -3 -3 3 3
use M3_M2  M3_M2_7189
timestamp 1745462530
transform 1 0 2460 0 1 3865
box -3 -3 3 3
use M3_M2  M3_M2_7190
timestamp 1745462530
transform 1 0 2460 0 1 3795
box -3 -3 3 3
use M3_M2  M3_M2_7191
timestamp 1745462530
transform 1 0 2612 0 1 3725
box -3 -3 3 3
use M3_M2  M3_M2_7192
timestamp 1745462530
transform 1 0 2500 0 1 3725
box -3 -3 3 3
use M3_M2  M3_M2_7193
timestamp 1745462530
transform 1 0 2324 0 1 4145
box -3 -3 3 3
use M3_M2  M3_M2_7194
timestamp 1745462530
transform 1 0 2316 0 1 3825
box -3 -3 3 3
use M3_M2  M3_M2_7195
timestamp 1745462530
transform 1 0 2292 0 1 4145
box -3 -3 3 3
use M3_M2  M3_M2_7196
timestamp 1745462530
transform 1 0 2292 0 1 4045
box -3 -3 3 3
use M3_M2  M3_M2_7197
timestamp 1745462530
transform 1 0 2284 0 1 3825
box -3 -3 3 3
use M3_M2  M3_M2_7198
timestamp 1745462530
transform 1 0 2276 0 1 4045
box -3 -3 3 3
use M3_M2  M3_M2_7199
timestamp 1745462530
transform 1 0 2316 0 1 3545
box -3 -3 3 3
use M3_M2  M3_M2_7200
timestamp 1745462530
transform 1 0 2284 0 1 3545
box -3 -3 3 3
use M3_M2  M3_M2_7201
timestamp 1745462530
transform 1 0 2308 0 1 3625
box -3 -3 3 3
use M3_M2  M3_M2_7202
timestamp 1745462530
transform 1 0 2284 0 1 3625
box -3 -3 3 3
use M3_M2  M3_M2_7203
timestamp 1745462530
transform 1 0 2564 0 1 3555
box -3 -3 3 3
use M3_M2  M3_M2_7204
timestamp 1745462530
transform 1 0 2324 0 1 3555
box -3 -3 3 3
use M3_M2  M3_M2_7205
timestamp 1745462530
transform 1 0 2684 0 1 3015
box -3 -3 3 3
use M3_M2  M3_M2_7206
timestamp 1745462530
transform 1 0 2628 0 1 3015
box -3 -3 3 3
use M3_M2  M3_M2_7207
timestamp 1745462530
transform 1 0 2684 0 1 3705
box -3 -3 3 3
use M3_M2  M3_M2_7208
timestamp 1745462530
transform 1 0 2636 0 1 3995
box -3 -3 3 3
use M3_M2  M3_M2_7209
timestamp 1745462530
transform 1 0 2596 0 1 3995
box -3 -3 3 3
use M3_M2  M3_M2_7210
timestamp 1745462530
transform 1 0 2596 0 1 3705
box -3 -3 3 3
use M3_M2  M3_M2_7211
timestamp 1745462530
transform 1 0 2716 0 1 3565
box -3 -3 3 3
use M3_M2  M3_M2_7212
timestamp 1745462530
transform 1 0 2668 0 1 3565
box -3 -3 3 3
use M3_M2  M3_M2_7213
timestamp 1745462530
transform 1 0 2748 0 1 3625
box -3 -3 3 3
use M3_M2  M3_M2_7214
timestamp 1745462530
transform 1 0 2708 0 1 3625
box -3 -3 3 3
use M3_M2  M3_M2_7215
timestamp 1745462530
transform 1 0 3852 0 1 3515
box -3 -3 3 3
use M3_M2  M3_M2_7216
timestamp 1745462530
transform 1 0 3804 0 1 3625
box -3 -3 3 3
use M3_M2  M3_M2_7217
timestamp 1745462530
transform 1 0 3780 0 1 3625
box -3 -3 3 3
use M3_M2  M3_M2_7218
timestamp 1745462530
transform 1 0 3780 0 1 3515
box -3 -3 3 3
use M3_M2  M3_M2_7219
timestamp 1745462530
transform 1 0 2884 0 1 3645
box -3 -3 3 3
use M3_M2  M3_M2_7220
timestamp 1745462530
transform 1 0 2716 0 1 3645
box -3 -3 3 3
use M3_M2  M3_M2_7221
timestamp 1745462530
transform 1 0 2004 0 1 3485
box -3 -3 3 3
use M3_M2  M3_M2_7222
timestamp 1745462530
transform 1 0 1884 0 1 3645
box -3 -3 3 3
use M3_M2  M3_M2_7223
timestamp 1745462530
transform 1 0 1884 0 1 3505
box -3 -3 3 3
use M3_M2  M3_M2_7224
timestamp 1745462530
transform 1 0 1884 0 1 3485
box -3 -3 3 3
use M3_M2  M3_M2_7225
timestamp 1745462530
transform 1 0 1812 0 1 3505
box -3 -3 3 3
use M3_M2  M3_M2_7226
timestamp 1745462530
transform 1 0 3676 0 1 3405
box -3 -3 3 3
use M3_M2  M3_M2_7227
timestamp 1745462530
transform 1 0 3636 0 1 3405
box -3 -3 3 3
use M3_M2  M3_M2_7228
timestamp 1745462530
transform 1 0 3636 0 1 3355
box -3 -3 3 3
use M3_M2  M3_M2_7229
timestamp 1745462530
transform 1 0 3604 0 1 3405
box -3 -3 3 3
use M3_M2  M3_M2_7230
timestamp 1745462530
transform 1 0 2940 0 1 3355
box -3 -3 3 3
use M3_M2  M3_M2_7231
timestamp 1745462530
transform 1 0 2692 0 1 3355
box -3 -3 3 3
use M3_M2  M3_M2_7232
timestamp 1745462530
transform 1 0 2444 0 1 3355
box -3 -3 3 3
use M3_M2  M3_M2_7233
timestamp 1745462530
transform 1 0 2324 0 1 3355
box -3 -3 3 3
use M3_M2  M3_M2_7234
timestamp 1745462530
transform 1 0 2300 0 1 3435
box -3 -3 3 3
use M3_M2  M3_M2_7235
timestamp 1745462530
transform 1 0 2180 0 1 3435
box -3 -3 3 3
use M3_M2  M3_M2_7236
timestamp 1745462530
transform 1 0 2740 0 1 3465
box -3 -3 3 3
use M3_M2  M3_M2_7237
timestamp 1745462530
transform 1 0 2716 0 1 3465
box -3 -3 3 3
use M3_M2  M3_M2_7238
timestamp 1745462530
transform 1 0 3588 0 1 3465
box -3 -3 3 3
use M3_M2  M3_M2_7239
timestamp 1745462530
transform 1 0 3556 0 1 3465
box -3 -3 3 3
use M3_M2  M3_M2_7240
timestamp 1745462530
transform 1 0 3548 0 1 3445
box -3 -3 3 3
use M3_M2  M3_M2_7241
timestamp 1745462530
transform 1 0 3508 0 1 3445
box -3 -3 3 3
use M3_M2  M3_M2_7242
timestamp 1745462530
transform 1 0 3460 0 1 3445
box -3 -3 3 3
use M3_M2  M3_M2_7243
timestamp 1745462530
transform 1 0 3460 0 1 3375
box -3 -3 3 3
use M3_M2  M3_M2_7244
timestamp 1745462530
transform 1 0 2916 0 1 3375
box -3 -3 3 3
use M3_M2  M3_M2_7245
timestamp 1745462530
transform 1 0 2756 0 1 3485
box -3 -3 3 3
use M3_M2  M3_M2_7246
timestamp 1745462530
transform 1 0 2756 0 1 3375
box -3 -3 3 3
use M3_M2  M3_M2_7247
timestamp 1745462530
transform 1 0 2596 0 1 3485
box -3 -3 3 3
use M3_M2  M3_M2_7248
timestamp 1745462530
transform 1 0 2564 0 1 3505
box -3 -3 3 3
use M3_M2  M3_M2_7249
timestamp 1745462530
transform 1 0 2524 0 1 3505
box -3 -3 3 3
use M3_M2  M3_M2_7250
timestamp 1745462530
transform 1 0 2956 0 1 3435
box -3 -3 3 3
use M3_M2  M3_M2_7251
timestamp 1745462530
transform 1 0 2908 0 1 3435
box -3 -3 3 3
use M3_M2  M3_M2_7252
timestamp 1745462530
transform 1 0 4268 0 1 3725
box -3 -3 3 3
use M3_M2  M3_M2_7253
timestamp 1745462530
transform 1 0 3876 0 1 3725
box -3 -3 3 3
use M3_M2  M3_M2_7254
timestamp 1745462530
transform 1 0 3844 0 1 3425
box -3 -3 3 3
use M3_M2  M3_M2_7255
timestamp 1745462530
transform 1 0 3700 0 1 3425
box -3 -3 3 3
use M3_M2  M3_M2_7256
timestamp 1745462530
transform 1 0 3692 0 1 3395
box -3 -3 3 3
use M3_M2  M3_M2_7257
timestamp 1745462530
transform 1 0 3532 0 1 3395
box -3 -3 3 3
use M3_M2  M3_M2_7258
timestamp 1745462530
transform 1 0 4196 0 1 3765
box -3 -3 3 3
use M3_M2  M3_M2_7259
timestamp 1745462530
transform 1 0 3892 0 1 3765
box -3 -3 3 3
use M3_M2  M3_M2_7260
timestamp 1745462530
transform 1 0 3876 0 1 3555
box -3 -3 3 3
use M3_M2  M3_M2_7261
timestamp 1745462530
transform 1 0 3756 0 1 3555
box -3 -3 3 3
use M3_M2  M3_M2_7262
timestamp 1745462530
transform 1 0 3884 0 1 3615
box -3 -3 3 3
use M3_M2  M3_M2_7263
timestamp 1745462530
transform 1 0 3796 0 1 3615
box -3 -3 3 3
use M3_M2  M3_M2_7264
timestamp 1745462530
transform 1 0 3724 0 1 3445
box -3 -3 3 3
use M3_M2  M3_M2_7265
timestamp 1745462530
transform 1 0 3572 0 1 3445
box -3 -3 3 3
use M3_M2  M3_M2_7266
timestamp 1745462530
transform 1 0 4228 0 1 3625
box -3 -3 3 3
use M3_M2  M3_M2_7267
timestamp 1745462530
transform 1 0 4204 0 1 3625
box -3 -3 3 3
use M3_M2  M3_M2_7268
timestamp 1745462530
transform 1 0 4204 0 1 3555
box -3 -3 3 3
use M3_M2  M3_M2_7269
timestamp 1745462530
transform 1 0 3900 0 1 3555
box -3 -3 3 3
use M3_M2  M3_M2_7270
timestamp 1745462530
transform 1 0 3924 0 1 3505
box -3 -3 3 3
use M3_M2  M3_M2_7271
timestamp 1745462530
transform 1 0 3884 0 1 3505
box -3 -3 3 3
use M3_M2  M3_M2_7272
timestamp 1745462530
transform 1 0 3884 0 1 3415
box -3 -3 3 3
use M3_M2  M3_M2_7273
timestamp 1745462530
transform 1 0 3620 0 1 3415
box -3 -3 3 3
use M3_M2  M3_M2_7274
timestamp 1745462530
transform 1 0 3612 0 1 3425
box -3 -3 3 3
use M3_M2  M3_M2_7275
timestamp 1745462530
transform 1 0 3492 0 1 3425
box -3 -3 3 3
use M3_M2  M3_M2_7276
timestamp 1745462530
transform 1 0 3964 0 1 3545
box -3 -3 3 3
use M3_M2  M3_M2_7277
timestamp 1745462530
transform 1 0 3908 0 1 3545
box -3 -3 3 3
use M3_M2  M3_M2_7278
timestamp 1745462530
transform 1 0 3852 0 1 3545
box -3 -3 3 3
use M3_M2  M3_M2_7279
timestamp 1745462530
transform 1 0 3804 0 1 3505
box -3 -3 3 3
use M3_M2  M3_M2_7280
timestamp 1745462530
transform 1 0 3652 0 1 3505
box -3 -3 3 3
use M3_M2  M3_M2_7281
timestamp 1745462530
transform 1 0 3660 0 1 3385
box -3 -3 3 3
use M3_M2  M3_M2_7282
timestamp 1745462530
transform 1 0 3572 0 1 3405
box -3 -3 3 3
use M3_M2  M3_M2_7283
timestamp 1745462530
transform 1 0 3572 0 1 3385
box -3 -3 3 3
use M3_M2  M3_M2_7284
timestamp 1745462530
transform 1 0 3452 0 1 3425
box -3 -3 3 3
use M3_M2  M3_M2_7285
timestamp 1745462530
transform 1 0 2452 0 1 3405
box -3 -3 3 3
use M3_M2  M3_M2_7286
timestamp 1745462530
transform 1 0 1956 0 1 3405
box -3 -3 3 3
use M3_M2  M3_M2_7287
timestamp 1745462530
transform 1 0 1972 0 1 3515
box -3 -3 3 3
use M3_M2  M3_M2_7288
timestamp 1745462530
transform 1 0 1948 0 1 3515
box -3 -3 3 3
use M3_M2  M3_M2_7289
timestamp 1745462530
transform 1 0 2500 0 1 3425
box -3 -3 3 3
use M3_M2  M3_M2_7290
timestamp 1745462530
transform 1 0 2484 0 1 3425
box -3 -3 3 3
use M3_M2  M3_M2_7291
timestamp 1745462530
transform 1 0 2060 0 1 3685
box -3 -3 3 3
use M3_M2  M3_M2_7292
timestamp 1745462530
transform 1 0 2052 0 1 3815
box -3 -3 3 3
use M3_M2  M3_M2_7293
timestamp 1745462530
transform 1 0 2044 0 1 3685
box -3 -3 3 3
use M3_M2  M3_M2_7294
timestamp 1745462530
transform 1 0 2020 0 1 3905
box -3 -3 3 3
use M3_M2  M3_M2_7295
timestamp 1745462530
transform 1 0 1996 0 1 3905
box -3 -3 3 3
use M3_M2  M3_M2_7296
timestamp 1745462530
transform 1 0 1996 0 1 3815
box -3 -3 3 3
use M3_M2  M3_M2_7297
timestamp 1745462530
transform 1 0 2340 0 1 3495
box -3 -3 3 3
use M3_M2  M3_M2_7298
timestamp 1745462530
transform 1 0 2044 0 1 3495
box -3 -3 3 3
use M3_M2  M3_M2_7299
timestamp 1745462530
transform 1 0 2548 0 1 3475
box -3 -3 3 3
use M3_M2  M3_M2_7300
timestamp 1745462530
transform 1 0 2452 0 1 3475
box -3 -3 3 3
use M3_M2  M3_M2_7301
timestamp 1745462530
transform 1 0 2452 0 1 3425
box -3 -3 3 3
use M3_M2  M3_M2_7302
timestamp 1745462530
transform 1 0 2356 0 1 3425
box -3 -3 3 3
use M3_M2  M3_M2_7303
timestamp 1745462530
transform 1 0 2740 0 1 3375
box -3 -3 3 3
use M3_M2  M3_M2_7304
timestamp 1745462530
transform 1 0 2668 0 1 3375
box -3 -3 3 3
use M3_M2  M3_M2_7305
timestamp 1745462530
transform 1 0 3820 0 1 3435
box -3 -3 3 3
use M3_M2  M3_M2_7306
timestamp 1745462530
transform 1 0 3740 0 1 3435
box -3 -3 3 3
use M3_M2  M3_M2_7307
timestamp 1745462530
transform 1 0 3004 0 1 3435
box -3 -3 3 3
use M3_M2  M3_M2_7308
timestamp 1745462530
transform 1 0 3004 0 1 3315
box -3 -3 3 3
use M3_M2  M3_M2_7309
timestamp 1745462530
transform 1 0 2868 0 1 3315
box -3 -3 3 3
use M3_M2  M3_M2_7310
timestamp 1745462530
transform 1 0 2868 0 1 3025
box -3 -3 3 3
use M3_M2  M3_M2_7311
timestamp 1745462530
transform 1 0 2668 0 1 3225
box -3 -3 3 3
use M3_M2  M3_M2_7312
timestamp 1745462530
transform 1 0 2668 0 1 3005
box -3 -3 3 3
use M3_M2  M3_M2_7313
timestamp 1745462530
transform 1 0 2620 0 1 3225
box -3 -3 3 3
use M3_M2  M3_M2_7314
timestamp 1745462530
transform 1 0 2540 0 1 3325
box -3 -3 3 3
use M3_M2  M3_M2_7315
timestamp 1745462530
transform 1 0 2540 0 1 3225
box -3 -3 3 3
use M3_M2  M3_M2_7316
timestamp 1745462530
transform 1 0 2508 0 1 3505
box -3 -3 3 3
use M3_M2  M3_M2_7317
timestamp 1745462530
transform 1 0 2508 0 1 3325
box -3 -3 3 3
use M3_M2  M3_M2_7318
timestamp 1745462530
transform 1 0 1972 0 1 3505
box -3 -3 3 3
use M3_M2  M3_M2_7319
timestamp 1745462530
transform 1 0 1972 0 1 3425
box -3 -3 3 3
use M3_M2  M3_M2_7320
timestamp 1745462530
transform 1 0 1900 0 1 3425
box -3 -3 3 3
use M3_M2  M3_M2_7321
timestamp 1745462530
transform 1 0 3628 0 1 3305
box -3 -3 3 3
use M3_M2  M3_M2_7322
timestamp 1745462530
transform 1 0 3588 0 1 3305
box -3 -3 3 3
use M3_M2  M3_M2_7323
timestamp 1745462530
transform 1 0 3572 0 1 3045
box -3 -3 3 3
use M3_M2  M3_M2_7324
timestamp 1745462530
transform 1 0 2940 0 1 3055
box -3 -3 3 3
use M3_M2  M3_M2_7325
timestamp 1745462530
transform 1 0 2700 0 1 3055
box -3 -3 3 3
use M3_M2  M3_M2_7326
timestamp 1745462530
transform 1 0 2460 0 1 3325
box -3 -3 3 3
use M3_M2  M3_M2_7327
timestamp 1745462530
transform 1 0 2380 0 1 3055
box -3 -3 3 3
use M3_M2  M3_M2_7328
timestamp 1745462530
transform 1 0 2364 0 1 3305
box -3 -3 3 3
use M3_M2  M3_M2_7329
timestamp 1745462530
transform 1 0 2356 0 1 3325
box -3 -3 3 3
use M3_M2  M3_M2_7330
timestamp 1745462530
transform 1 0 2116 0 1 3305
box -3 -3 3 3
use M3_M2  M3_M2_7331
timestamp 1745462530
transform 1 0 3500 0 1 3325
box -3 -3 3 3
use M3_M2  M3_M2_7332
timestamp 1745462530
transform 1 0 3468 0 1 3325
box -3 -3 3 3
use M3_M2  M3_M2_7333
timestamp 1745462530
transform 1 0 3420 0 1 3325
box -3 -3 3 3
use M3_M2  M3_M2_7334
timestamp 1745462530
transform 1 0 3420 0 1 3265
box -3 -3 3 3
use M3_M2  M3_M2_7335
timestamp 1745462530
transform 1 0 3388 0 1 3265
box -3 -3 3 3
use M3_M2  M3_M2_7336
timestamp 1745462530
transform 1 0 2956 0 1 3325
box -3 -3 3 3
use M3_M2  M3_M2_7337
timestamp 1745462530
transform 1 0 2780 0 1 3325
box -3 -3 3 3
use M3_M2  M3_M2_7338
timestamp 1745462530
transform 1 0 2660 0 1 3765
box -3 -3 3 3
use M3_M2  M3_M2_7339
timestamp 1745462530
transform 1 0 2620 0 1 3765
box -3 -3 3 3
use M3_M2  M3_M2_7340
timestamp 1745462530
transform 1 0 2612 0 1 3475
box -3 -3 3 3
use M3_M2  M3_M2_7341
timestamp 1745462530
transform 1 0 2588 0 1 3325
box -3 -3 3 3
use M3_M2  M3_M2_7342
timestamp 1745462530
transform 1 0 2572 0 1 3475
box -3 -3 3 3
use M3_M2  M3_M2_7343
timestamp 1745462530
transform 1 0 2964 0 1 3485
box -3 -3 3 3
use M3_M2  M3_M2_7344
timestamp 1745462530
transform 1 0 2916 0 1 3635
box -3 -3 3 3
use M3_M2  M3_M2_7345
timestamp 1745462530
transform 1 0 2916 0 1 3485
box -3 -3 3 3
use M3_M2  M3_M2_7346
timestamp 1745462530
transform 1 0 2900 0 1 3725
box -3 -3 3 3
use M3_M2  M3_M2_7347
timestamp 1745462530
transform 1 0 2868 0 1 3725
box -3 -3 3 3
use M3_M2  M3_M2_7348
timestamp 1745462530
transform 1 0 2860 0 1 3635
box -3 -3 3 3
use M3_M2  M3_M2_7349
timestamp 1745462530
transform 1 0 2988 0 1 3295
box -3 -3 3 3
use M3_M2  M3_M2_7350
timestamp 1745462530
transform 1 0 2948 0 1 3295
box -3 -3 3 3
use M3_M2  M3_M2_7351
timestamp 1745462530
transform 1 0 4076 0 1 3505
box -3 -3 3 3
use M3_M2  M3_M2_7352
timestamp 1745462530
transform 1 0 3996 0 1 3515
box -3 -3 3 3
use M3_M2  M3_M2_7353
timestamp 1745462530
transform 1 0 3892 0 1 3515
box -3 -3 3 3
use M3_M2  M3_M2_7354
timestamp 1745462530
transform 1 0 3868 0 1 3335
box -3 -3 3 3
use M3_M2  M3_M2_7355
timestamp 1745462530
transform 1 0 3636 0 1 3335
box -3 -3 3 3
use M3_M2  M3_M2_7356
timestamp 1745462530
transform 1 0 3892 0 1 3315
box -3 -3 3 3
use M3_M2  M3_M2_7357
timestamp 1745462530
transform 1 0 3804 0 1 3315
box -3 -3 3 3
use M3_M2  M3_M2_7358
timestamp 1745462530
transform 1 0 3644 0 1 3295
box -3 -3 3 3
use M3_M2  M3_M2_7359
timestamp 1745462530
transform 1 0 3460 0 1 3295
box -3 -3 3 3
use M3_M2  M3_M2_7360
timestamp 1745462530
transform 1 0 4020 0 1 3495
box -3 -3 3 3
use M3_M2  M3_M2_7361
timestamp 1745462530
transform 1 0 3924 0 1 3495
box -3 -3 3 3
use M3_M2  M3_M2_7362
timestamp 1745462530
transform 1 0 3876 0 1 3375
box -3 -3 3 3
use M3_M2  M3_M2_7363
timestamp 1745462530
transform 1 0 3692 0 1 3375
box -3 -3 3 3
use M3_M2  M3_M2_7364
timestamp 1745462530
transform 1 0 3916 0 1 3395
box -3 -3 3 3
use M3_M2  M3_M2_7365
timestamp 1745462530
transform 1 0 3836 0 1 3395
box -3 -3 3 3
use M3_M2  M3_M2_7366
timestamp 1745462530
transform 1 0 3676 0 1 3325
box -3 -3 3 3
use M3_M2  M3_M2_7367
timestamp 1745462530
transform 1 0 3516 0 1 3325
box -3 -3 3 3
use M3_M2  M3_M2_7368
timestamp 1745462530
transform 1 0 4172 0 1 3395
box -3 -3 3 3
use M3_M2  M3_M2_7369
timestamp 1745462530
transform 1 0 4140 0 1 3395
box -3 -3 3 3
use M3_M2  M3_M2_7370
timestamp 1745462530
transform 1 0 3932 0 1 3395
box -3 -3 3 3
use M3_M2  M3_M2_7371
timestamp 1745462530
transform 1 0 3924 0 1 3345
box -3 -3 3 3
use M3_M2  M3_M2_7372
timestamp 1745462530
transform 1 0 3572 0 1 3345
box -3 -3 3 3
use M3_M2  M3_M2_7373
timestamp 1745462530
transform 1 0 3940 0 1 3445
box -3 -3 3 3
use M3_M2  M3_M2_7374
timestamp 1745462530
transform 1 0 3900 0 1 3445
box -3 -3 3 3
use M3_M2  M3_M2_7375
timestamp 1745462530
transform 1 0 3556 0 1 3315
box -3 -3 3 3
use M3_M2  M3_M2_7376
timestamp 1745462530
transform 1 0 3412 0 1 3315
box -3 -3 3 3
use M3_M2  M3_M2_7377
timestamp 1745462530
transform 1 0 3940 0 1 3385
box -3 -3 3 3
use M3_M2  M3_M2_7378
timestamp 1745462530
transform 1 0 3804 0 1 3385
box -3 -3 3 3
use M3_M2  M3_M2_7379
timestamp 1745462530
transform 1 0 3772 0 1 3365
box -3 -3 3 3
use M3_M2  M3_M2_7380
timestamp 1745462530
transform 1 0 3612 0 1 3365
box -3 -3 3 3
use M3_M2  M3_M2_7381
timestamp 1745462530
transform 1 0 3804 0 1 3445
box -3 -3 3 3
use M3_M2  M3_M2_7382
timestamp 1745462530
transform 1 0 3772 0 1 3445
box -3 -3 3 3
use M3_M2  M3_M2_7383
timestamp 1745462530
transform 1 0 3604 0 1 3275
box -3 -3 3 3
use M3_M2  M3_M2_7384
timestamp 1745462530
transform 1 0 3364 0 1 3275
box -3 -3 3 3
use M3_M2  M3_M2_7385
timestamp 1745462530
transform 1 0 2052 0 1 3565
box -3 -3 3 3
use M3_M2  M3_M2_7386
timestamp 1745462530
transform 1 0 2004 0 1 3565
box -3 -3 3 3
use M3_M2  M3_M2_7387
timestamp 1745462530
transform 1 0 2460 0 1 3335
box -3 -3 3 3
use M3_M2  M3_M2_7388
timestamp 1745462530
transform 1 0 2020 0 1 3335
box -3 -3 3 3
use M3_M2  M3_M2_7389
timestamp 1745462530
transform 1 0 2044 0 1 3425
box -3 -3 3 3
use M3_M2  M3_M2_7390
timestamp 1745462530
transform 1 0 2020 0 1 3425
box -3 -3 3 3
use M3_M2  M3_M2_7391
timestamp 1745462530
transform 1 0 1964 0 1 3925
box -3 -3 3 3
use M3_M2  M3_M2_7392
timestamp 1745462530
transform 1 0 1940 0 1 3925
box -3 -3 3 3
use M3_M2  M3_M2_7393
timestamp 1745462530
transform 1 0 2412 0 1 3375
box -3 -3 3 3
use M3_M2  M3_M2_7394
timestamp 1745462530
transform 1 0 1932 0 1 3375
box -3 -3 3 3
use M3_M2  M3_M2_7395
timestamp 1745462530
transform 1 0 2580 0 1 3365
box -3 -3 3 3
use M3_M2  M3_M2_7396
timestamp 1745462530
transform 1 0 2428 0 1 3365
box -3 -3 3 3
use M3_M2  M3_M2_7397
timestamp 1745462530
transform 1 0 2796 0 1 2975
box -3 -3 3 3
use M3_M2  M3_M2_7398
timestamp 1745462530
transform 1 0 2756 0 1 2975
box -3 -3 3 3
use M3_M2  M3_M2_7399
timestamp 1745462530
transform 1 0 2036 0 1 3605
box -3 -3 3 3
use M3_M2  M3_M2_7400
timestamp 1745462530
transform 1 0 1884 0 1 3745
box -3 -3 3 3
use M3_M2  M3_M2_7401
timestamp 1745462530
transform 1 0 1844 0 1 3745
box -3 -3 3 3
use M3_M2  M3_M2_7402
timestamp 1745462530
transform 1 0 1844 0 1 3605
box -3 -3 3 3
use M3_M2  M3_M2_7403
timestamp 1745462530
transform 1 0 2684 0 1 3175
box -3 -3 3 3
use M3_M2  M3_M2_7404
timestamp 1745462530
transform 1 0 2020 0 1 3175
box -3 -3 3 3
use M3_M2  M3_M2_7405
timestamp 1745462530
transform 1 0 3812 0 1 3305
box -3 -3 3 3
use M3_M2  M3_M2_7406
timestamp 1745462530
transform 1 0 3796 0 1 3115
box -3 -3 3 3
use M3_M2  M3_M2_7407
timestamp 1745462530
transform 1 0 3708 0 1 3305
box -3 -3 3 3
use M3_M2  M3_M2_7408
timestamp 1745462530
transform 1 0 2020 0 1 3145
box -3 -3 3 3
use M3_M2  M3_M2_7409
timestamp 1745462530
transform 1 0 2020 0 1 3115
box -3 -3 3 3
use M3_M2  M3_M2_7410
timestamp 1745462530
transform 1 0 1948 0 1 3225
box -3 -3 3 3
use M3_M2  M3_M2_7411
timestamp 1745462530
transform 1 0 1940 0 1 3145
box -3 -3 3 3
use M3_M2  M3_M2_7412
timestamp 1745462530
transform 1 0 1828 0 1 3365
box -3 -3 3 3
use M3_M2  M3_M2_7413
timestamp 1745462530
transform 1 0 1812 0 1 3365
box -3 -3 3 3
use M3_M2  M3_M2_7414
timestamp 1745462530
transform 1 0 1812 0 1 3225
box -3 -3 3 3
use M3_M2  M3_M2_7415
timestamp 1745462530
transform 1 0 3564 0 1 3135
box -3 -3 3 3
use M3_M2  M3_M2_7416
timestamp 1745462530
transform 1 0 3532 0 1 3135
box -3 -3 3 3
use M3_M2  M3_M2_7417
timestamp 1745462530
transform 1 0 2812 0 1 3335
box -3 -3 3 3
use M3_M2  M3_M2_7418
timestamp 1745462530
transform 1 0 2812 0 1 3135
box -3 -3 3 3
use M3_M2  M3_M2_7419
timestamp 1745462530
transform 1 0 2692 0 1 3345
box -3 -3 3 3
use M3_M2  M3_M2_7420
timestamp 1745462530
transform 1 0 2660 0 1 3195
box -3 -3 3 3
use M3_M2  M3_M2_7421
timestamp 1745462530
transform 1 0 2476 0 1 3195
box -3 -3 3 3
use M3_M2  M3_M2_7422
timestamp 1745462530
transform 1 0 2308 0 1 3195
box -3 -3 3 3
use M3_M2  M3_M2_7423
timestamp 1745462530
transform 1 0 2276 0 1 3195
box -3 -3 3 3
use M3_M2  M3_M2_7424
timestamp 1745462530
transform 1 0 2780 0 1 3225
box -3 -3 3 3
use M3_M2  M3_M2_7425
timestamp 1745462530
transform 1 0 2708 0 1 3225
box -3 -3 3 3
use M3_M2  M3_M2_7426
timestamp 1745462530
transform 1 0 3516 0 1 3065
box -3 -3 3 3
use M3_M2  M3_M2_7427
timestamp 1745462530
transform 1 0 3500 0 1 3215
box -3 -3 3 3
use M3_M2  M3_M2_7428
timestamp 1745462530
transform 1 0 3460 0 1 3065
box -3 -3 3 3
use M3_M2  M3_M2_7429
timestamp 1745462530
transform 1 0 3404 0 1 3065
box -3 -3 3 3
use M3_M2  M3_M2_7430
timestamp 1745462530
transform 1 0 3388 0 1 3215
box -3 -3 3 3
use M3_M2  M3_M2_7431
timestamp 1745462530
transform 1 0 2876 0 1 3195
box -3 -3 3 3
use M3_M2  M3_M2_7432
timestamp 1745462530
transform 1 0 2804 0 1 3225
box -3 -3 3 3
use M3_M2  M3_M2_7433
timestamp 1745462530
transform 1 0 2572 0 1 3205
box -3 -3 3 3
use M3_M2  M3_M2_7434
timestamp 1745462530
transform 1 0 2468 0 1 3315
box -3 -3 3 3
use M3_M2  M3_M2_7435
timestamp 1745462530
transform 1 0 2468 0 1 3215
box -3 -3 3 3
use M3_M2  M3_M2_7436
timestamp 1745462530
transform 1 0 1908 0 1 3565
box -3 -3 3 3
use M3_M2  M3_M2_7437
timestamp 1745462530
transform 1 0 1868 0 1 3565
box -3 -3 3 3
use M3_M2  M3_M2_7438
timestamp 1745462530
transform 1 0 1868 0 1 3315
box -3 -3 3 3
use M3_M2  M3_M2_7439
timestamp 1745462530
transform 1 0 1948 0 1 3575
box -3 -3 3 3
use M3_M2  M3_M2_7440
timestamp 1745462530
transform 1 0 1940 0 1 3905
box -3 -3 3 3
use M3_M2  M3_M2_7441
timestamp 1745462530
transform 1 0 1916 0 1 3575
box -3 -3 3 3
use M3_M2  M3_M2_7442
timestamp 1745462530
transform 1 0 1820 0 1 3965
box -3 -3 3 3
use M3_M2  M3_M2_7443
timestamp 1745462530
transform 1 0 1788 0 1 3965
box -3 -3 3 3
use M3_M2  M3_M2_7444
timestamp 1745462530
transform 1 0 1788 0 1 3905
box -3 -3 3 3
use M3_M2  M3_M2_7445
timestamp 1745462530
transform 1 0 2844 0 1 3295
box -3 -3 3 3
use M3_M2  M3_M2_7446
timestamp 1745462530
transform 1 0 1932 0 1 3305
box -3 -3 3 3
use M3_M2  M3_M2_7447
timestamp 1745462530
transform 1 0 2004 0 1 3365
box -3 -3 3 3
use M3_M2  M3_M2_7448
timestamp 1745462530
transform 1 0 1980 0 1 3365
box -3 -3 3 3
use M3_M2  M3_M2_7449
timestamp 1745462530
transform 1 0 4204 0 1 3325
box -3 -3 3 3
use M3_M2  M3_M2_7450
timestamp 1745462530
transform 1 0 3900 0 1 3325
box -3 -3 3 3
use M3_M2  M3_M2_7451
timestamp 1745462530
transform 1 0 3860 0 1 3155
box -3 -3 3 3
use M3_M2  M3_M2_7452
timestamp 1745462530
transform 1 0 3636 0 1 3155
box -3 -3 3 3
use M3_M2  M3_M2_7453
timestamp 1745462530
transform 1 0 3884 0 1 3215
box -3 -3 3 3
use M3_M2  M3_M2_7454
timestamp 1745462530
transform 1 0 3820 0 1 3215
box -3 -3 3 3
use M3_M2  M3_M2_7455
timestamp 1745462530
transform 1 0 3612 0 1 3105
box -3 -3 3 3
use M3_M2  M3_M2_7456
timestamp 1745462530
transform 1 0 3500 0 1 3105
box -3 -3 3 3
use M3_M2  M3_M2_7457
timestamp 1745462530
transform 1 0 4188 0 1 3365
box -3 -3 3 3
use M3_M2  M3_M2_7458
timestamp 1745462530
transform 1 0 3876 0 1 3365
box -3 -3 3 3
use M3_M2  M3_M2_7459
timestamp 1745462530
transform 1 0 3844 0 1 3255
box -3 -3 3 3
use M3_M2  M3_M2_7460
timestamp 1745462530
transform 1 0 3612 0 1 3255
box -3 -3 3 3
use M3_M2  M3_M2_7461
timestamp 1745462530
transform 1 0 3596 0 1 3095
box -3 -3 3 3
use M3_M2  M3_M2_7462
timestamp 1745462530
transform 1 0 3484 0 1 3095
box -3 -3 3 3
use M3_M2  M3_M2_7463
timestamp 1745462530
transform 1 0 4036 0 1 3225
box -3 -3 3 3
use M3_M2  M3_M2_7464
timestamp 1745462530
transform 1 0 3988 0 1 3215
box -3 -3 3 3
use M3_M2  M3_M2_7465
timestamp 1745462530
transform 1 0 3924 0 1 3215
box -3 -3 3 3
use M3_M2  M3_M2_7466
timestamp 1745462530
transform 1 0 3892 0 1 3175
box -3 -3 3 3
use M3_M2  M3_M2_7467
timestamp 1745462530
transform 1 0 3580 0 1 3175
box -3 -3 3 3
use M3_M2  M3_M2_7468
timestamp 1745462530
transform 1 0 3916 0 1 3195
box -3 -3 3 3
use M3_M2  M3_M2_7469
timestamp 1745462530
transform 1 0 3852 0 1 3195
box -3 -3 3 3
use M3_M2  M3_M2_7470
timestamp 1745462530
transform 1 0 3564 0 1 3085
box -3 -3 3 3
use M3_M2  M3_M2_7471
timestamp 1745462530
transform 1 0 3444 0 1 3085
box -3 -3 3 3
use M3_M2  M3_M2_7472
timestamp 1745462530
transform 1 0 3932 0 1 3165
box -3 -3 3 3
use M3_M2  M3_M2_7473
timestamp 1745462530
transform 1 0 3708 0 1 3165
box -3 -3 3 3
use M3_M2  M3_M2_7474
timestamp 1745462530
transform 1 0 3668 0 1 3195
box -3 -3 3 3
use M3_M2  M3_M2_7475
timestamp 1745462530
transform 1 0 3556 0 1 3195
box -3 -3 3 3
use M3_M2  M3_M2_7476
timestamp 1745462530
transform 1 0 3564 0 1 3155
box -3 -3 3 3
use M3_M2  M3_M2_7477
timestamp 1745462530
transform 1 0 3396 0 1 3155
box -3 -3 3 3
use M3_M2  M3_M2_7478
timestamp 1745462530
transform 1 0 1876 0 1 3465
box -3 -3 3 3
use M3_M2  M3_M2_7479
timestamp 1745462530
transform 1 0 1700 0 1 3795
box -3 -3 3 3
use M3_M2  M3_M2_7480
timestamp 1745462530
transform 1 0 1668 0 1 3795
box -3 -3 3 3
use M3_M2  M3_M2_7481
timestamp 1745462530
transform 1 0 1668 0 1 3465
box -3 -3 3 3
use M3_M2  M3_M2_7482
timestamp 1745462530
transform 1 0 2508 0 1 3185
box -3 -3 3 3
use M3_M2  M3_M2_7483
timestamp 1745462530
transform 1 0 1868 0 1 3185
box -3 -3 3 3
use M3_M2  M3_M2_7484
timestamp 1745462530
transform 1 0 2556 0 1 3205
box -3 -3 3 3
use M3_M2  M3_M2_7485
timestamp 1745462530
transform 1 0 2532 0 1 3205
box -3 -3 3 3
use M3_M2  M3_M2_7486
timestamp 1745462530
transform 1 0 1828 0 1 3305
box -3 -3 3 3
use M3_M2  M3_M2_7487
timestamp 1745462530
transform 1 0 1740 0 1 3405
box -3 -3 3 3
use M3_M2  M3_M2_7488
timestamp 1745462530
transform 1 0 1740 0 1 3305
box -3 -3 3 3
use M3_M2  M3_M2_7489
timestamp 1745462530
transform 1 0 1716 0 1 3825
box -3 -3 3 3
use M3_M2  M3_M2_7490
timestamp 1745462530
transform 1 0 1716 0 1 3585
box -3 -3 3 3
use M3_M2  M3_M2_7491
timestamp 1745462530
transform 1 0 1692 0 1 3925
box -3 -3 3 3
use M3_M2  M3_M2_7492
timestamp 1745462530
transform 1 0 1692 0 1 3825
box -3 -3 3 3
use M3_M2  M3_M2_7493
timestamp 1745462530
transform 1 0 1660 0 1 3925
box -3 -3 3 3
use M3_M2  M3_M2_7494
timestamp 1745462530
transform 1 0 1660 0 1 3585
box -3 -3 3 3
use M3_M2  M3_M2_7495
timestamp 1745462530
transform 1 0 1660 0 1 3405
box -3 -3 3 3
use M3_M2  M3_M2_7496
timestamp 1745462530
transform 1 0 2316 0 1 3155
box -3 -3 3 3
use M3_M2  M3_M2_7497
timestamp 1745462530
transform 1 0 1812 0 1 3155
box -3 -3 3 3
use M3_M2  M3_M2_7498
timestamp 1745462530
transform 1 0 2524 0 1 3085
box -3 -3 3 3
use M3_M2  M3_M2_7499
timestamp 1745462530
transform 1 0 2364 0 1 3085
box -3 -3 3 3
use M3_M2  M3_M2_7500
timestamp 1745462530
transform 1 0 2756 0 1 3085
box -3 -3 3 3
use M3_M2  M3_M2_7501
timestamp 1745462530
transform 1 0 2724 0 1 3085
box -3 -3 3 3
use M3_M2  M3_M2_7502
timestamp 1745462530
transform 1 0 2308 0 1 3325
box -3 -3 3 3
use M3_M2  M3_M2_7503
timestamp 1745462530
transform 1 0 2212 0 1 3325
box -3 -3 3 3
use M3_M2  M3_M2_7504
timestamp 1745462530
transform 1 0 2156 0 1 3325
box -3 -3 3 3
use M3_M2  M3_M2_7505
timestamp 1745462530
transform 1 0 1764 0 1 3515
box -3 -3 3 3
use M3_M2  M3_M2_7506
timestamp 1745462530
transform 1 0 1756 0 1 3935
box -3 -3 3 3
use M3_M2  M3_M2_7507
timestamp 1745462530
transform 1 0 1748 0 1 3505
box -3 -3 3 3
use M3_M2  M3_M2_7508
timestamp 1745462530
transform 1 0 1716 0 1 3935
box -3 -3 3 3
use M3_M2  M3_M2_7509
timestamp 1745462530
transform 1 0 2628 0 1 3285
box -3 -3 3 3
use M3_M2  M3_M2_7510
timestamp 1745462530
transform 1 0 1756 0 1 3285
box -3 -3 3 3
use M3_M2  M3_M2_7511
timestamp 1745462530
transform 1 0 1828 0 1 3345
box -3 -3 3 3
use M3_M2  M3_M2_7512
timestamp 1745462530
transform 1 0 1780 0 1 3345
box -3 -3 3 3
use M3_M2  M3_M2_7513
timestamp 1745462530
transform 1 0 3756 0 1 3195
box -3 -3 3 3
use M3_M2  M3_M2_7514
timestamp 1745462530
transform 1 0 3732 0 1 3195
box -3 -3 3 3
use M3_M2  M3_M2_7515
timestamp 1745462530
transform 1 0 3652 0 1 3185
box -3 -3 3 3
use M3_M2  M3_M2_7516
timestamp 1745462530
transform 1 0 3628 0 1 3075
box -3 -3 3 3
use M3_M2  M3_M2_7517
timestamp 1745462530
transform 1 0 3188 0 1 3235
box -3 -3 3 3
use M3_M2  M3_M2_7518
timestamp 1745462530
transform 1 0 3180 0 1 3075
box -3 -3 3 3
use M3_M2  M3_M2_7519
timestamp 1745462530
transform 1 0 3180 0 1 2965
box -3 -3 3 3
use M3_M2  M3_M2_7520
timestamp 1745462530
transform 1 0 3084 0 1 3235
box -3 -3 3 3
use M3_M2  M3_M2_7521
timestamp 1745462530
transform 1 0 2164 0 1 2945
box -3 -3 3 3
use M3_M2  M3_M2_7522
timestamp 1745462530
transform 1 0 2140 0 1 3245
box -3 -3 3 3
use M3_M2  M3_M2_7523
timestamp 1745462530
transform 1 0 2092 0 1 3245
box -3 -3 3 3
use M3_M2  M3_M2_7524
timestamp 1745462530
transform 1 0 2084 0 1 3295
box -3 -3 3 3
use M3_M2  M3_M2_7525
timestamp 1745462530
transform 1 0 1860 0 1 3405
box -3 -3 3 3
use M3_M2  M3_M2_7526
timestamp 1745462530
transform 1 0 1860 0 1 3305
box -3 -3 3 3
use M3_M2  M3_M2_7527
timestamp 1745462530
transform 1 0 1804 0 1 3405
box -3 -3 3 3
use M3_M2  M3_M2_7528
timestamp 1745462530
transform 1 0 1756 0 1 3405
box -3 -3 3 3
use M3_M2  M3_M2_7529
timestamp 1745462530
transform 1 0 3420 0 1 3245
box -3 -3 3 3
use M3_M2  M3_M2_7530
timestamp 1745462530
transform 1 0 3404 0 1 3245
box -3 -3 3 3
use M3_M2  M3_M2_7531
timestamp 1745462530
transform 1 0 3340 0 1 3245
box -3 -3 3 3
use M3_M2  M3_M2_7532
timestamp 1745462530
transform 1 0 3228 0 1 3245
box -3 -3 3 3
use M3_M2  M3_M2_7533
timestamp 1745462530
transform 1 0 2828 0 1 3245
box -3 -3 3 3
use M3_M2  M3_M2_7534
timestamp 1745462530
transform 1 0 2740 0 1 3285
box -3 -3 3 3
use M3_M2  M3_M2_7535
timestamp 1745462530
transform 1 0 2740 0 1 3245
box -3 -3 3 3
use M3_M2  M3_M2_7536
timestamp 1745462530
transform 1 0 2652 0 1 3305
box -3 -3 3 3
use M3_M2  M3_M2_7537
timestamp 1745462530
transform 1 0 2652 0 1 3285
box -3 -3 3 3
use M3_M2  M3_M2_7538
timestamp 1745462530
transform 1 0 2580 0 1 3305
box -3 -3 3 3
use M3_M2  M3_M2_7539
timestamp 1745462530
transform 1 0 2380 0 1 3305
box -3 -3 3 3
use M3_M2  M3_M2_7540
timestamp 1745462530
transform 1 0 2372 0 1 3225
box -3 -3 3 3
use M3_M2  M3_M2_7541
timestamp 1745462530
transform 1 0 2300 0 1 3225
box -3 -3 3 3
use M3_M2  M3_M2_7542
timestamp 1745462530
transform 1 0 2724 0 1 3205
box -3 -3 3 3
use M3_M2  M3_M2_7543
timestamp 1745462530
transform 1 0 2652 0 1 3205
box -3 -3 3 3
use M3_M2  M3_M2_7544
timestamp 1745462530
transform 1 0 3356 0 1 3225
box -3 -3 3 3
use M3_M2  M3_M2_7545
timestamp 1745462530
transform 1 0 3324 0 1 3225
box -3 -3 3 3
use M3_M2  M3_M2_7546
timestamp 1745462530
transform 1 0 3276 0 1 3225
box -3 -3 3 3
use M3_M2  M3_M2_7547
timestamp 1745462530
transform 1 0 2908 0 1 3225
box -3 -3 3 3
use M3_M2  M3_M2_7548
timestamp 1745462530
transform 1 0 2828 0 1 3225
box -3 -3 3 3
use M3_M2  M3_M2_7549
timestamp 1745462530
transform 1 0 2828 0 1 3205
box -3 -3 3 3
use M3_M2  M3_M2_7550
timestamp 1745462530
transform 1 0 2828 0 1 3065
box -3 -3 3 3
use M3_M2  M3_M2_7551
timestamp 1745462530
transform 1 0 2740 0 1 3205
box -3 -3 3 3
use M3_M2  M3_M2_7552
timestamp 1745462530
transform 1 0 2620 0 1 3065
box -3 -3 3 3
use M3_M2  M3_M2_7553
timestamp 1745462530
transform 1 0 2620 0 1 3045
box -3 -3 3 3
use M3_M2  M3_M2_7554
timestamp 1745462530
transform 1 0 2460 0 1 3045
box -3 -3 3 3
use M3_M2  M3_M2_7555
timestamp 1745462530
transform 1 0 2452 0 1 3225
box -3 -3 3 3
use M3_M2  M3_M2_7556
timestamp 1745462530
transform 1 0 1836 0 1 3215
box -3 -3 3 3
use M3_M2  M3_M2_7557
timestamp 1745462530
transform 1 0 1828 0 1 3595
box -3 -3 3 3
use M3_M2  M3_M2_7558
timestamp 1745462530
transform 1 0 1804 0 1 3595
box -3 -3 3 3
use M3_M2  M3_M2_7559
timestamp 1745462530
transform 1 0 1924 0 1 3755
box -3 -3 3 3
use M3_M2  M3_M2_7560
timestamp 1745462530
transform 1 0 1924 0 1 3685
box -3 -3 3 3
use M3_M2  M3_M2_7561
timestamp 1745462530
transform 1 0 1892 0 1 3685
box -3 -3 3 3
use M3_M2  M3_M2_7562
timestamp 1745462530
transform 1 0 1780 0 1 3985
box -3 -3 3 3
use M3_M2  M3_M2_7563
timestamp 1745462530
transform 1 0 1780 0 1 3755
box -3 -3 3 3
use M3_M2  M3_M2_7564
timestamp 1745462530
transform 1 0 1740 0 1 3985
box -3 -3 3 3
use M3_M2  M3_M2_7565
timestamp 1745462530
transform 1 0 1692 0 1 3985
box -3 -3 3 3
use M3_M2  M3_M2_7566
timestamp 1745462530
transform 1 0 2844 0 1 3315
box -3 -3 3 3
use M3_M2  M3_M2_7567
timestamp 1745462530
transform 1 0 1956 0 1 3365
box -3 -3 3 3
use M3_M2  M3_M2_7568
timestamp 1745462530
transform 1 0 1956 0 1 3345
box -3 -3 3 3
use M3_M2  M3_M2_7569
timestamp 1745462530
transform 1 0 1900 0 1 3365
box -3 -3 3 3
use M3_M2  M3_M2_7570
timestamp 1745462530
transform 1 0 2892 0 1 3255
box -3 -3 3 3
use M3_M2  M3_M2_7571
timestamp 1745462530
transform 1 0 2860 0 1 3255
box -3 -3 3 3
use M3_M2  M3_M2_7572
timestamp 1745462530
transform 1 0 3084 0 1 3015
box -3 -3 3 3
use M3_M2  M3_M2_7573
timestamp 1745462530
transform 1 0 3036 0 1 3015
box -3 -3 3 3
use M3_M2  M3_M2_7574
timestamp 1745462530
transform 1 0 2980 0 1 3015
box -3 -3 3 3
use M3_M2  M3_M2_7575
timestamp 1745462530
transform 1 0 2964 0 1 2405
box -3 -3 3 3
use M3_M2  M3_M2_7576
timestamp 1745462530
transform 1 0 2964 0 1 1815
box -3 -3 3 3
use M3_M2  M3_M2_7577
timestamp 1745462530
transform 1 0 2908 0 1 2405
box -3 -3 3 3
use M3_M2  M3_M2_7578
timestamp 1745462530
transform 1 0 2564 0 1 1815
box -3 -3 3 3
use M3_M2  M3_M2_7579
timestamp 1745462530
transform 1 0 2964 0 1 2885
box -3 -3 3 3
use M3_M2  M3_M2_7580
timestamp 1745462530
transform 1 0 2956 0 1 3015
box -3 -3 3 3
use M3_M2  M3_M2_7581
timestamp 1745462530
transform 1 0 2916 0 1 2845
box -3 -3 3 3
use M3_M2  M3_M2_7582
timestamp 1745462530
transform 1 0 2916 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_7583
timestamp 1745462530
transform 1 0 2900 0 1 3015
box -3 -3 3 3
use M3_M2  M3_M2_7584
timestamp 1745462530
transform 1 0 2876 0 1 2885
box -3 -3 3 3
use M3_M2  M3_M2_7585
timestamp 1745462530
transform 1 0 2876 0 1 2845
box -3 -3 3 3
use M3_M2  M3_M2_7586
timestamp 1745462530
transform 1 0 2868 0 1 2375
box -3 -3 3 3
use M3_M2  M3_M2_7587
timestamp 1745462530
transform 1 0 2860 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_7588
timestamp 1745462530
transform 1 0 2460 0 1 2375
box -3 -3 3 3
use M3_M2  M3_M2_7589
timestamp 1745462530
transform 1 0 4172 0 1 3145
box -3 -3 3 3
use M3_M2  M3_M2_7590
timestamp 1745462530
transform 1 0 3804 0 1 3145
box -3 -3 3 3
use M3_M2  M3_M2_7591
timestamp 1745462530
transform 1 0 3732 0 1 3145
box -3 -3 3 3
use M3_M2  M3_M2_7592
timestamp 1745462530
transform 1 0 3372 0 1 3145
box -3 -3 3 3
use M3_M2  M3_M2_7593
timestamp 1745462530
transform 1 0 3348 0 1 3085
box -3 -3 3 3
use M3_M2  M3_M2_7594
timestamp 1745462530
transform 1 0 3284 0 1 3085
box -3 -3 3 3
use M3_M2  M3_M2_7595
timestamp 1745462530
transform 1 0 3156 0 1 3055
box -3 -3 3 3
use M3_M2  M3_M2_7596
timestamp 1745462530
transform 1 0 3068 0 1 3055
box -3 -3 3 3
use M3_M2  M3_M2_7597
timestamp 1745462530
transform 1 0 3060 0 1 3035
box -3 -3 3 3
use M3_M2  M3_M2_7598
timestamp 1745462530
transform 1 0 2972 0 1 3035
box -3 -3 3 3
use M3_M2  M3_M2_7599
timestamp 1745462530
transform 1 0 2900 0 1 3035
box -3 -3 3 3
use M3_M2  M3_M2_7600
timestamp 1745462530
transform 1 0 2892 0 1 3065
box -3 -3 3 3
use M3_M2  M3_M2_7601
timestamp 1745462530
transform 1 0 2852 0 1 3065
box -3 -3 3 3
use M3_M2  M3_M2_7602
timestamp 1745462530
transform 1 0 2732 0 1 3035
box -3 -3 3 3
use M3_M2  M3_M2_7603
timestamp 1745462530
transform 1 0 2732 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_7604
timestamp 1745462530
transform 1 0 2620 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_7605
timestamp 1745462530
transform 1 0 2604 0 1 2055
box -3 -3 3 3
use M3_M2  M3_M2_7606
timestamp 1745462530
transform 1 0 2588 0 1 2055
box -3 -3 3 3
use M3_M2  M3_M2_7607
timestamp 1745462530
transform 1 0 4188 0 1 3185
box -3 -3 3 3
use M3_M2  M3_M2_7608
timestamp 1745462530
transform 1 0 3740 0 1 3185
box -3 -3 3 3
use M3_M2  M3_M2_7609
timestamp 1745462530
transform 1 0 3716 0 1 3205
box -3 -3 3 3
use M3_M2  M3_M2_7610
timestamp 1745462530
transform 1 0 3452 0 1 3185
box -3 -3 3 3
use M3_M2  M3_M2_7611
timestamp 1745462530
transform 1 0 3452 0 1 3225
box -3 -3 3 3
use M3_M2  M3_M2_7612
timestamp 1745462530
transform 1 0 3366 0 1 3225
box -3 -3 3 3
use M3_M2  M3_M2_7613
timestamp 1745462530
transform 1 0 3188 0 1 3195
box -3 -3 3 3
use M3_M2  M3_M2_7614
timestamp 1745462530
transform 1 0 3108 0 1 3195
box -3 -3 3 3
use M3_M2  M3_M2_7615
timestamp 1745462530
transform 1 0 4076 0 1 3345
box -3 -3 3 3
use M3_M2  M3_M2_7616
timestamp 1745462530
transform 1 0 4036 0 1 3345
box -3 -3 3 3
use M3_M2  M3_M2_7617
timestamp 1745462530
transform 1 0 4028 0 1 3275
box -3 -3 3 3
use M3_M2  M3_M2_7618
timestamp 1745462530
transform 1 0 3636 0 1 3275
box -3 -3 3 3
use M3_M2  M3_M2_7619
timestamp 1745462530
transform 1 0 3604 0 1 3265
box -3 -3 3 3
use M3_M2  M3_M2_7620
timestamp 1745462530
transform 1 0 3444 0 1 3265
box -3 -3 3 3
use M3_M2  M3_M2_7621
timestamp 1745462530
transform 1 0 3428 0 1 3205
box -3 -3 3 3
use M3_M2  M3_M2_7622
timestamp 1745462530
transform 1 0 3308 0 1 3205
box -3 -3 3 3
use M3_M2  M3_M2_7623
timestamp 1745462530
transform 1 0 3172 0 1 3085
box -3 -3 3 3
use M3_M2  M3_M2_7624
timestamp 1745462530
transform 1 0 3028 0 1 3085
box -3 -3 3 3
use M3_M2  M3_M2_7625
timestamp 1745462530
transform 1 0 3788 0 1 3235
box -3 -3 3 3
use M3_M2  M3_M2_7626
timestamp 1745462530
transform 1 0 3276 0 1 3235
box -3 -3 3 3
use M3_M2  M3_M2_7627
timestamp 1745462530
transform 1 0 3268 0 1 3255
box -3 -3 3 3
use M3_M2  M3_M2_7628
timestamp 1745462530
transform 1 0 3116 0 1 3265
box -3 -3 3 3
use M3_M2  M3_M2_7629
timestamp 1745462530
transform 1 0 2092 0 1 3655
box -3 -3 3 3
use M3_M2  M3_M2_7630
timestamp 1745462530
transform 1 0 1604 0 1 3655
box -3 -3 3 3
use M3_M2  M3_M2_7631
timestamp 1745462530
transform 1 0 1596 0 1 3755
box -3 -3 3 3
use M3_M2  M3_M2_7632
timestamp 1745462530
transform 1 0 1564 0 1 3755
box -3 -3 3 3
use M3_M2  M3_M2_7633
timestamp 1745462530
transform 1 0 2380 0 1 3205
box -3 -3 3 3
use M3_M2  M3_M2_7634
timestamp 1745462530
transform 1 0 2092 0 1 3205
box -3 -3 3 3
use M3_M2  M3_M2_7635
timestamp 1745462530
transform 1 0 2156 0 1 3195
box -3 -3 3 3
use M3_M2  M3_M2_7636
timestamp 1745462530
transform 1 0 2124 0 1 3195
box -3 -3 3 3
use M3_M2  M3_M2_7637
timestamp 1745462530
transform 1 0 2436 0 1 3225
box -3 -3 3 3
use M3_M2  M3_M2_7638
timestamp 1745462530
transform 1 0 2420 0 1 3225
box -3 -3 3 3
use M3_M2  M3_M2_7639
timestamp 1745462530
transform 1 0 2860 0 1 3045
box -3 -3 3 3
use M3_M2  M3_M2_7640
timestamp 1745462530
transform 1 0 2788 0 1 3045
box -3 -3 3 3
use M3_M2  M3_M2_7641
timestamp 1745462530
transform 1 0 2876 0 1 3345
box -3 -3 3 3
use M3_M2  M3_M2_7642
timestamp 1745462530
transform 1 0 2820 0 1 3345
box -3 -3 3 3
use M3_M2  M3_M2_7643
timestamp 1745462530
transform 1 0 2836 0 1 3435
box -3 -3 3 3
use M3_M2  M3_M2_7644
timestamp 1745462530
transform 1 0 2820 0 1 3435
box -3 -3 3 3
use M3_M2  M3_M2_7645
timestamp 1745462530
transform 1 0 2244 0 1 3885
box -3 -3 3 3
use M3_M2  M3_M2_7646
timestamp 1745462530
transform 1 0 1636 0 1 3895
box -3 -3 3 3
use M3_M2  M3_M2_7647
timestamp 1745462530
transform 1 0 1628 0 1 3795
box -3 -3 3 3
use M3_M2  M3_M2_7648
timestamp 1745462530
transform 1 0 1596 0 1 3795
box -3 -3 3 3
use M3_M2  M3_M2_7649
timestamp 1745462530
transform 1 0 2292 0 1 3135
box -3 -3 3 3
use M3_M2  M3_M2_7650
timestamp 1745462530
transform 1 0 2236 0 1 3135
box -3 -3 3 3
use M3_M2  M3_M2_7651
timestamp 1745462530
transform 1 0 2444 0 1 3065
box -3 -3 3 3
use M3_M2  M3_M2_7652
timestamp 1745462530
transform 1 0 2332 0 1 3065
box -3 -3 3 3
use M3_M2  M3_M2_7653
timestamp 1745462530
transform 1 0 2932 0 1 3095
box -3 -3 3 3
use M3_M2  M3_M2_7654
timestamp 1745462530
transform 1 0 2804 0 1 3085
box -3 -3 3 3
use M3_M2  M3_M2_7655
timestamp 1745462530
transform 1 0 3724 0 1 1615
box -3 -3 3 3
use M3_M2  M3_M2_7656
timestamp 1745462530
transform 1 0 2484 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_7657
timestamp 1745462530
transform 1 0 2492 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_7658
timestamp 1745462530
transform 1 0 2076 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_7659
timestamp 1745462530
transform 1 0 2028 0 1 1845
box -3 -3 3 3
use M3_M2  M3_M2_7660
timestamp 1745462530
transform 1 0 1012 0 1 1845
box -3 -3 3 3
use M3_M2  M3_M2_7661
timestamp 1745462530
transform 1 0 2060 0 1 1775
box -3 -3 3 3
use M3_M2  M3_M2_7662
timestamp 1745462530
transform 1 0 876 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_7663
timestamp 1745462530
transform 1 0 876 0 1 1775
box -3 -3 3 3
use M3_M2  M3_M2_7664
timestamp 1745462530
transform 1 0 828 0 1 2235
box -3 -3 3 3
use M3_M2  M3_M2_7665
timestamp 1745462530
transform 1 0 804 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_7666
timestamp 1745462530
transform 1 0 804 0 1 2015
box -3 -3 3 3
use M3_M2  M3_M2_7667
timestamp 1745462530
transform 1 0 804 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_7668
timestamp 1745462530
transform 1 0 804 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_7669
timestamp 1745462530
transform 1 0 764 0 1 2235
box -3 -3 3 3
use M3_M2  M3_M2_7670
timestamp 1745462530
transform 1 0 764 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_7671
timestamp 1745462530
transform 1 0 2532 0 1 2665
box -3 -3 3 3
use M3_M2  M3_M2_7672
timestamp 1745462530
transform 1 0 2460 0 1 2665
box -3 -3 3 3
use M3_M2  M3_M2_7673
timestamp 1745462530
transform 1 0 2548 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_7674
timestamp 1745462530
transform 1 0 2516 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_7675
timestamp 1745462530
transform 1 0 2484 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_7676
timestamp 1745462530
transform 1 0 2468 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_7677
timestamp 1745462530
transform 1 0 2436 0 1 2455
box -3 -3 3 3
use M3_M2  M3_M2_7678
timestamp 1745462530
transform 1 0 2412 0 1 2455
box -3 -3 3 3
use M3_M2  M3_M2_7679
timestamp 1745462530
transform 1 0 2412 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_7680
timestamp 1745462530
transform 1 0 2052 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_7681
timestamp 1745462530
transform 1 0 2020 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_7682
timestamp 1745462530
transform 1 0 2484 0 1 2705
box -3 -3 3 3
use M3_M2  M3_M2_7683
timestamp 1745462530
transform 1 0 2452 0 1 2705
box -3 -3 3 3
use M3_M2  M3_M2_7684
timestamp 1745462530
transform 1 0 2436 0 1 2705
box -3 -3 3 3
use M3_M2  M3_M2_7685
timestamp 1745462530
transform 1 0 2636 0 1 2695
box -3 -3 3 3
use M3_M2  M3_M2_7686
timestamp 1745462530
transform 1 0 2596 0 1 2695
box -3 -3 3 3
use M3_M2  M3_M2_7687
timestamp 1745462530
transform 1 0 2548 0 1 2565
box -3 -3 3 3
use M3_M2  M3_M2_7688
timestamp 1745462530
transform 1 0 2532 0 1 2565
box -3 -3 3 3
use M3_M2  M3_M2_7689
timestamp 1745462530
transform 1 0 2484 0 1 2055
box -3 -3 3 3
use M3_M2  M3_M2_7690
timestamp 1745462530
transform 1 0 2452 0 1 2055
box -3 -3 3 3
use M3_M2  M3_M2_7691
timestamp 1745462530
transform 1 0 2164 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_7692
timestamp 1745462530
transform 1 0 2092 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_7693
timestamp 1745462530
transform 1 0 2348 0 1 2085
box -3 -3 3 3
use M3_M2  M3_M2_7694
timestamp 1745462530
transform 1 0 2324 0 1 2085
box -3 -3 3 3
use M3_M2  M3_M2_7695
timestamp 1745462530
transform 1 0 2300 0 1 2085
box -3 -3 3 3
use M3_M2  M3_M2_7696
timestamp 1745462530
transform 1 0 2420 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_7697
timestamp 1745462530
transform 1 0 2404 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_7698
timestamp 1745462530
transform 1 0 2388 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_7699
timestamp 1745462530
transform 1 0 828 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_7700
timestamp 1745462530
transform 1 0 740 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_7701
timestamp 1745462530
transform 1 0 852 0 1 2445
box -3 -3 3 3
use M3_M2  M3_M2_7702
timestamp 1745462530
transform 1 0 844 0 1 2575
box -3 -3 3 3
use M3_M2  M3_M2_7703
timestamp 1745462530
transform 1 0 820 0 1 2575
box -3 -3 3 3
use M3_M2  M3_M2_7704
timestamp 1745462530
transform 1 0 812 0 1 2425
box -3 -3 3 3
use M3_M2  M3_M2_7705
timestamp 1745462530
transform 1 0 980 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_7706
timestamp 1745462530
transform 1 0 964 0 1 1815
box -3 -3 3 3
use M3_M2  M3_M2_7707
timestamp 1745462530
transform 1 0 2116 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_7708
timestamp 1745462530
transform 1 0 2068 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_7709
timestamp 1745462530
transform 1 0 3724 0 1 1575
box -3 -3 3 3
use M3_M2  M3_M2_7710
timestamp 1745462530
transform 1 0 3700 0 1 1575
box -3 -3 3 3
use M3_M2  M3_M2_7711
timestamp 1745462530
transform 1 0 3732 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_7712
timestamp 1745462530
transform 1 0 3692 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_7713
timestamp 1745462530
transform 1 0 3828 0 1 2235
box -3 -3 3 3
use M3_M2  M3_M2_7714
timestamp 1745462530
transform 1 0 3828 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_7715
timestamp 1745462530
transform 1 0 3788 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_7716
timestamp 1745462530
transform 1 0 3780 0 1 2235
box -3 -3 3 3
use M3_M2  M3_M2_7717
timestamp 1745462530
transform 1 0 3732 0 1 1885
box -3 -3 3 3
use M3_M2  M3_M2_7718
timestamp 1745462530
transform 1 0 3692 0 1 2015
box -3 -3 3 3
use M3_M2  M3_M2_7719
timestamp 1745462530
transform 1 0 3692 0 1 1885
box -3 -3 3 3
use M3_M2  M3_M2_7720
timestamp 1745462530
transform 1 0 3660 0 1 2015
box -3 -3 3 3
use M3_M2  M3_M2_7721
timestamp 1745462530
transform 1 0 3788 0 1 2545
box -3 -3 3 3
use M3_M2  M3_M2_7722
timestamp 1745462530
transform 1 0 3708 0 1 2555
box -3 -3 3 3
use M3_M2  M3_M2_7723
timestamp 1745462530
transform 1 0 3740 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_7724
timestamp 1745462530
transform 1 0 3684 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_7725
timestamp 1745462530
transform 1 0 3820 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_7726
timestamp 1745462530
transform 1 0 3780 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_7727
timestamp 1745462530
transform 1 0 3788 0 1 2355
box -3 -3 3 3
use M3_M2  M3_M2_7728
timestamp 1745462530
transform 1 0 3180 0 1 2385
box -3 -3 3 3
use M3_M2  M3_M2_7729
timestamp 1745462530
transform 1 0 3180 0 1 2355
box -3 -3 3 3
use M3_M2  M3_M2_7730
timestamp 1745462530
transform 1 0 3124 0 1 2385
box -3 -3 3 3
use M3_M2  M3_M2_7731
timestamp 1745462530
transform 1 0 3780 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_7732
timestamp 1745462530
transform 1 0 3700 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_7733
timestamp 1745462530
transform 1 0 3716 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_7734
timestamp 1745462530
transform 1 0 3660 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_7735
timestamp 1745462530
transform 1 0 3764 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_7736
timestamp 1745462530
transform 1 0 3692 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_7737
timestamp 1745462530
transform 1 0 3820 0 1 975
box -3 -3 3 3
use M3_M2  M3_M2_7738
timestamp 1745462530
transform 1 0 3772 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_7739
timestamp 1745462530
transform 1 0 3772 0 1 975
box -3 -3 3 3
use M3_M2  M3_M2_7740
timestamp 1745462530
transform 1 0 3716 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_7741
timestamp 1745462530
transform 1 0 3740 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_7742
timestamp 1745462530
transform 1 0 3716 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_7743
timestamp 1745462530
transform 1 0 2508 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_7744
timestamp 1745462530
transform 1 0 1908 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_7745
timestamp 1745462530
transform 1 0 2012 0 1 2265
box -3 -3 3 3
use M3_M2  M3_M2_7746
timestamp 1745462530
transform 1 0 2012 0 1 2065
box -3 -3 3 3
use M3_M2  M3_M2_7747
timestamp 1745462530
transform 1 0 1916 0 1 2265
box -3 -3 3 3
use M3_M2  M3_M2_7748
timestamp 1745462530
transform 1 0 1916 0 1 2065
box -3 -3 3 3
use M3_M2  M3_M2_7749
timestamp 1745462530
transform 1 0 1924 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_7750
timestamp 1745462530
transform 1 0 1148 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_7751
timestamp 1745462530
transform 1 0 1924 0 1 1465
box -3 -3 3 3
use M3_M2  M3_M2_7752
timestamp 1745462530
transform 1 0 796 0 1 1465
box -3 -3 3 3
use M3_M2  M3_M2_7753
timestamp 1745462530
transform 1 0 828 0 1 815
box -3 -3 3 3
use M3_M2  M3_M2_7754
timestamp 1745462530
transform 1 0 780 0 1 815
box -3 -3 3 3
use M3_M2  M3_M2_7755
timestamp 1745462530
transform 1 0 804 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_7756
timestamp 1745462530
transform 1 0 732 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_7757
timestamp 1745462530
transform 1 0 828 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_7758
timestamp 1745462530
transform 1 0 788 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_7759
timestamp 1745462530
transform 1 0 1116 0 1 1085
box -3 -3 3 3
use M3_M2  M3_M2_7760
timestamp 1745462530
transform 1 0 1004 0 1 1085
box -3 -3 3 3
use M3_M2  M3_M2_7761
timestamp 1745462530
transform 1 0 1124 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_7762
timestamp 1745462530
transform 1 0 1100 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_7763
timestamp 1745462530
transform 1 0 1972 0 1 2535
box -3 -3 3 3
use M3_M2  M3_M2_7764
timestamp 1745462530
transform 1 0 1924 0 1 2535
box -3 -3 3 3
use M3_M2  M3_M2_7765
timestamp 1745462530
transform 1 0 1884 0 1 2565
box -3 -3 3 3
use M3_M2  M3_M2_7766
timestamp 1745462530
transform 1 0 1852 0 1 2565
box -3 -3 3 3
use M3_M2  M3_M2_7767
timestamp 1745462530
transform 1 0 1924 0 1 1895
box -3 -3 3 3
use M3_M2  M3_M2_7768
timestamp 1745462530
transform 1 0 1868 0 1 1895
box -3 -3 3 3
use M3_M2  M3_M2_7769
timestamp 1745462530
transform 1 0 1956 0 1 1835
box -3 -3 3 3
use M3_M2  M3_M2_7770
timestamp 1745462530
transform 1 0 1924 0 1 1835
box -3 -3 3 3
use M3_M2  M3_M2_7771
timestamp 1745462530
transform 1 0 2628 0 1 1485
box -3 -3 3 3
use M3_M2  M3_M2_7772
timestamp 1745462530
transform 1 0 2548 0 1 1485
box -3 -3 3 3
use M3_M2  M3_M2_7773
timestamp 1745462530
transform 1 0 3148 0 1 1415
box -3 -3 3 3
use M3_M2  M3_M2_7774
timestamp 1745462530
transform 1 0 2548 0 1 1405
box -3 -3 3 3
use M3_M2  M3_M2_7775
timestamp 1745462530
transform 1 0 3740 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_7776
timestamp 1745462530
transform 1 0 3468 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_7777
timestamp 1745462530
transform 1 0 3468 0 1 1405
box -3 -3 3 3
use M3_M2  M3_M2_7778
timestamp 1745462530
transform 1 0 3132 0 1 1405
box -3 -3 3 3
use M3_M2  M3_M2_7779
timestamp 1745462530
transform 1 0 3212 0 1 1465
box -3 -3 3 3
use M3_M2  M3_M2_7780
timestamp 1745462530
transform 1 0 3172 0 1 1465
box -3 -3 3 3
use M3_M2  M3_M2_7781
timestamp 1745462530
transform 1 0 3748 0 1 1535
box -3 -3 3 3
use M3_M2  M3_M2_7782
timestamp 1745462530
transform 1 0 3740 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_7783
timestamp 1745462530
transform 1 0 3724 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_7784
timestamp 1745462530
transform 1 0 2620 0 1 1535
box -3 -3 3 3
use M3_M2  M3_M2_7785
timestamp 1745462530
transform 1 0 2564 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_7786
timestamp 1745462530
transform 1 0 2564 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_7787
timestamp 1745462530
transform 1 0 2548 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_7788
timestamp 1745462530
transform 1 0 2508 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_7789
timestamp 1745462530
transform 1 0 2564 0 1 1665
box -3 -3 3 3
use M3_M2  M3_M2_7790
timestamp 1745462530
transform 1 0 2492 0 1 1665
box -3 -3 3 3
use M3_M2  M3_M2_7791
timestamp 1745462530
transform 1 0 2588 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_7792
timestamp 1745462530
transform 1 0 2468 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_7793
timestamp 1745462530
transform 1 0 3516 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_7794
timestamp 1745462530
transform 1 0 2428 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_7795
timestamp 1745462530
transform 1 0 2420 0 1 1685
box -3 -3 3 3
use M3_M2  M3_M2_7796
timestamp 1745462530
transform 1 0 1060 0 1 1685
box -3 -3 3 3
use M3_M2  M3_M2_7797
timestamp 1745462530
transform 1 0 1068 0 1 2375
box -3 -3 3 3
use M3_M2  M3_M2_7798
timestamp 1745462530
transform 1 0 828 0 1 2375
box -3 -3 3 3
use M3_M2  M3_M2_7799
timestamp 1745462530
transform 1 0 1140 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_7800
timestamp 1745462530
transform 1 0 1100 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_7801
timestamp 1745462530
transform 1 0 1084 0 1 975
box -3 -3 3 3
use M3_M2  M3_M2_7802
timestamp 1745462530
transform 1 0 1036 0 1 975
box -3 -3 3 3
use M3_M2  M3_M2_7803
timestamp 1745462530
transform 1 0 1236 0 1 1535
box -3 -3 3 3
use M3_M2  M3_M2_7804
timestamp 1745462530
transform 1 0 1212 0 1 1535
box -3 -3 3 3
use M3_M2  M3_M2_7805
timestamp 1745462530
transform 1 0 820 0 1 2405
box -3 -3 3 3
use M3_M2  M3_M2_7806
timestamp 1745462530
transform 1 0 756 0 1 2405
box -3 -3 3 3
use M3_M2  M3_M2_7807
timestamp 1745462530
transform 1 0 996 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_7808
timestamp 1745462530
transform 1 0 940 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_7809
timestamp 1745462530
transform 1 0 956 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_7810
timestamp 1745462530
transform 1 0 916 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_7811
timestamp 1745462530
transform 1 0 3540 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_7812
timestamp 1745462530
transform 1 0 3508 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_7813
timestamp 1745462530
transform 1 0 3556 0 1 2485
box -3 -3 3 3
use M3_M2  M3_M2_7814
timestamp 1745462530
transform 1 0 3524 0 1 1935
box -3 -3 3 3
use M3_M2  M3_M2_7815
timestamp 1745462530
transform 1 0 3492 0 1 2485
box -3 -3 3 3
use M3_M2  M3_M2_7816
timestamp 1745462530
transform 1 0 3492 0 1 1935
box -3 -3 3 3
use M3_M2  M3_M2_7817
timestamp 1745462530
transform 1 0 3644 0 1 2555
box -3 -3 3 3
use M3_M2  M3_M2_7818
timestamp 1745462530
transform 1 0 3556 0 1 2555
box -3 -3 3 3
use M3_M2  M3_M2_7819
timestamp 1745462530
transform 1 0 3588 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_7820
timestamp 1745462530
transform 1 0 3516 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_7821
timestamp 1745462530
transform 1 0 3660 0 1 2695
box -3 -3 3 3
use M3_M2  M3_M2_7822
timestamp 1745462530
transform 1 0 3596 0 1 2695
box -3 -3 3 3
use M3_M2  M3_M2_7823
timestamp 1745462530
transform 1 0 3564 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_7824
timestamp 1745462530
transform 1 0 3524 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_7825
timestamp 1745462530
transform 1 0 3532 0 1 2295
box -3 -3 3 3
use M3_M2  M3_M2_7826
timestamp 1745462530
transform 1 0 3068 0 1 2295
box -3 -3 3 3
use M3_M2  M3_M2_7827
timestamp 1745462530
transform 1 0 3636 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_7828
timestamp 1745462530
transform 1 0 3540 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_7829
timestamp 1745462530
transform 1 0 3596 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_7830
timestamp 1745462530
transform 1 0 3572 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_7831
timestamp 1745462530
transform 1 0 3708 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_7832
timestamp 1745462530
transform 1 0 3524 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_7833
timestamp 1745462530
transform 1 0 3564 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_7834
timestamp 1745462530
transform 1 0 3524 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_7835
timestamp 1745462530
transform 1 0 2836 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_7836
timestamp 1745462530
transform 1 0 2428 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_7837
timestamp 1745462530
transform 1 0 2404 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_7838
timestamp 1745462530
transform 1 0 1396 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_7839
timestamp 1745462530
transform 1 0 1428 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_7840
timestamp 1745462530
transform 1 0 1388 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_7841
timestamp 1745462530
transform 1 0 1420 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_7842
timestamp 1745462530
transform 1 0 1188 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_7843
timestamp 1745462530
transform 1 0 1404 0 1 1275
box -3 -3 3 3
use M3_M2  M3_M2_7844
timestamp 1745462530
transform 1 0 932 0 1 1275
box -3 -3 3 3
use M3_M2  M3_M2_7845
timestamp 1745462530
transform 1 0 924 0 1 1085
box -3 -3 3 3
use M3_M2  M3_M2_7846
timestamp 1745462530
transform 1 0 788 0 1 1085
box -3 -3 3 3
use M3_M2  M3_M2_7847
timestamp 1745462530
transform 1 0 956 0 1 1205
box -3 -3 3 3
use M3_M2  M3_M2_7848
timestamp 1745462530
transform 1 0 924 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_7849
timestamp 1745462530
transform 1 0 924 0 1 1205
box -3 -3 3 3
use M3_M2  M3_M2_7850
timestamp 1745462530
transform 1 0 892 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_7851
timestamp 1745462530
transform 1 0 812 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_7852
timestamp 1745462530
transform 1 0 572 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_7853
timestamp 1745462530
transform 1 0 1156 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_7854
timestamp 1745462530
transform 1 0 1028 0 1 1065
box -3 -3 3 3
use M3_M2  M3_M2_7855
timestamp 1745462530
transform 1 0 1020 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_7856
timestamp 1745462530
transform 1 0 1012 0 1 1065
box -3 -3 3 3
use M3_M2  M3_M2_7857
timestamp 1745462530
transform 1 0 1500 0 1 2725
box -3 -3 3 3
use M3_M2  M3_M2_7858
timestamp 1745462530
transform 1 0 1412 0 1 2725
box -3 -3 3 3
use M3_M2  M3_M2_7859
timestamp 1745462530
transform 1 0 1476 0 1 2535
box -3 -3 3 3
use M3_M2  M3_M2_7860
timestamp 1745462530
transform 1 0 1452 0 1 2535
box -3 -3 3 3
use M3_M2  M3_M2_7861
timestamp 1745462530
transform 1 0 1532 0 1 2785
box -3 -3 3 3
use M3_M2  M3_M2_7862
timestamp 1745462530
transform 1 0 1516 0 1 2785
box -3 -3 3 3
use M3_M2  M3_M2_7863
timestamp 1745462530
transform 1 0 1460 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_7864
timestamp 1745462530
transform 1 0 1388 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_7865
timestamp 1745462530
transform 1 0 2820 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_7866
timestamp 1745462530
transform 1 0 2796 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_7867
timestamp 1745462530
transform 1 0 3244 0 1 1865
box -3 -3 3 3
use M3_M2  M3_M2_7868
timestamp 1745462530
transform 1 0 2812 0 1 1865
box -3 -3 3 3
use M3_M2  M3_M2_7869
timestamp 1745462530
transform 1 0 3412 0 1 1935
box -3 -3 3 3
use M3_M2  M3_M2_7870
timestamp 1745462530
transform 1 0 3252 0 1 1935
box -3 -3 3 3
use M3_M2  M3_M2_7871
timestamp 1745462530
transform 1 0 3268 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_7872
timestamp 1745462530
transform 1 0 3212 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_7873
timestamp 1745462530
transform 1 0 3588 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_7874
timestamp 1745462530
transform 1 0 3444 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_7875
timestamp 1745462530
transform 1 0 3388 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_7876
timestamp 1745462530
transform 1 0 2780 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_7877
timestamp 1745462530
transform 1 0 2812 0 1 875
box -3 -3 3 3
use M3_M2  M3_M2_7878
timestamp 1745462530
transform 1 0 2780 0 1 875
box -3 -3 3 3
use M3_M2  M3_M2_7879
timestamp 1745462530
transform 1 0 2796 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_7880
timestamp 1745462530
transform 1 0 2756 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_7881
timestamp 1745462530
transform 1 0 2812 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_7882
timestamp 1745462530
transform 1 0 2716 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_7883
timestamp 1745462530
transform 1 0 2812 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_7884
timestamp 1745462530
transform 1 0 2772 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_7885
timestamp 1745462530
transform 1 0 3380 0 1 1885
box -3 -3 3 3
use M3_M2  M3_M2_7886
timestamp 1745462530
transform 1 0 2468 0 1 1885
box -3 -3 3 3
use M3_M2  M3_M2_7887
timestamp 1745462530
transform 1 0 2444 0 1 1815
box -3 -3 3 3
use M3_M2  M3_M2_7888
timestamp 1745462530
transform 1 0 1116 0 1 1815
box -3 -3 3 3
use M3_M2  M3_M2_7889
timestamp 1745462530
transform 1 0 1100 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_7890
timestamp 1745462530
transform 1 0 892 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_7891
timestamp 1745462530
transform 1 0 1196 0 1 1645
box -3 -3 3 3
use M3_M2  M3_M2_7892
timestamp 1745462530
transform 1 0 1140 0 1 1645
box -3 -3 3 3
use M3_M2  M3_M2_7893
timestamp 1745462530
transform 1 0 1164 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_7894
timestamp 1745462530
transform 1 0 1108 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_7895
timestamp 1745462530
transform 1 0 1284 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_7896
timestamp 1745462530
transform 1 0 1252 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_7897
timestamp 1745462530
transform 1 0 916 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_7898
timestamp 1745462530
transform 1 0 868 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_7899
timestamp 1745462530
transform 1 0 876 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_7900
timestamp 1745462530
transform 1 0 852 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_7901
timestamp 1745462530
transform 1 0 3404 0 1 1865
box -3 -3 3 3
use M3_M2  M3_M2_7902
timestamp 1745462530
transform 1 0 3356 0 1 1865
box -3 -3 3 3
use M3_M2  M3_M2_7903
timestamp 1745462530
transform 1 0 3404 0 1 2155
box -3 -3 3 3
use M3_M2  M3_M2_7904
timestamp 1745462530
transform 1 0 3316 0 1 2155
box -3 -3 3 3
use M3_M2  M3_M2_7905
timestamp 1745462530
transform 1 0 3404 0 1 2245
box -3 -3 3 3
use M3_M2  M3_M2_7906
timestamp 1745462530
transform 1 0 3356 0 1 2555
box -3 -3 3 3
use M3_M2  M3_M2_7907
timestamp 1745462530
transform 1 0 3340 0 1 2555
box -3 -3 3 3
use M3_M2  M3_M2_7908
timestamp 1745462530
transform 1 0 3340 0 1 2245
box -3 -3 3 3
use M3_M2  M3_M2_7909
timestamp 1745462530
transform 1 0 3452 0 1 2565
box -3 -3 3 3
use M3_M2  M3_M2_7910
timestamp 1745462530
transform 1 0 3380 0 1 2565
box -3 -3 3 3
use M3_M2  M3_M2_7911
timestamp 1745462530
transform 1 0 3396 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_7912
timestamp 1745462530
transform 1 0 3284 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_7913
timestamp 1745462530
transform 1 0 3524 0 1 2725
box -3 -3 3 3
use M3_M2  M3_M2_7914
timestamp 1745462530
transform 1 0 3468 0 1 2725
box -3 -3 3 3
use M3_M2  M3_M2_7915
timestamp 1745462530
transform 1 0 3316 0 1 2245
box -3 -3 3 3
use M3_M2  M3_M2_7916
timestamp 1745462530
transform 1 0 3292 0 1 2245
box -3 -3 3 3
use M3_M2  M3_M2_7917
timestamp 1745462530
transform 1 0 3316 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_7918
timestamp 1745462530
transform 1 0 3236 0 1 2245
box -3 -3 3 3
use M3_M2  M3_M2_7919
timestamp 1745462530
transform 1 0 3236 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_7920
timestamp 1745462530
transform 1 0 2892 0 1 2235
box -3 -3 3 3
use M3_M2  M3_M2_7921
timestamp 1745462530
transform 1 0 3404 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_7922
timestamp 1745462530
transform 1 0 3356 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_7923
timestamp 1745462530
transform 1 0 3364 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_7924
timestamp 1745462530
transform 1 0 3308 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_7925
timestamp 1745462530
transform 1 0 3412 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_7926
timestamp 1745462530
transform 1 0 3380 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_7927
timestamp 1745462530
transform 1 0 3404 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_7928
timestamp 1745462530
transform 1 0 3380 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_7929
timestamp 1745462530
transform 1 0 2508 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_7930
timestamp 1745462530
transform 1 0 2396 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_7931
timestamp 1745462530
transform 1 0 2404 0 1 1875
box -3 -3 3 3
use M3_M2  M3_M2_7932
timestamp 1745462530
transform 1 0 1172 0 1 1875
box -3 -3 3 3
use M3_M2  M3_M2_7933
timestamp 1745462530
transform 1 0 1180 0 1 2405
box -3 -3 3 3
use M3_M2  M3_M2_7934
timestamp 1745462530
transform 1 0 1132 0 1 2405
box -3 -3 3 3
use M3_M2  M3_M2_7935
timestamp 1745462530
transform 1 0 1196 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_7936
timestamp 1745462530
transform 1 0 916 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_7937
timestamp 1745462530
transform 1 0 916 0 1 1135
box -3 -3 3 3
use M3_M2  M3_M2_7938
timestamp 1745462530
transform 1 0 860 0 1 1135
box -3 -3 3 3
use M3_M2  M3_M2_7939
timestamp 1745462530
transform 1 0 956 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_7940
timestamp 1745462530
transform 1 0 892 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_7941
timestamp 1745462530
transform 1 0 852 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_7942
timestamp 1745462530
transform 1 0 628 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_7943
timestamp 1745462530
transform 1 0 1188 0 1 1265
box -3 -3 3 3
use M3_M2  M3_M2_7944
timestamp 1745462530
transform 1 0 1156 0 1 1265
box -3 -3 3 3
use M3_M2  M3_M2_7945
timestamp 1745462530
transform 1 0 1156 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_7946
timestamp 1745462530
transform 1 0 964 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_7947
timestamp 1745462530
transform 1 0 1220 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_7948
timestamp 1745462530
transform 1 0 1188 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_7949
timestamp 1745462530
transform 1 0 1196 0 1 2725
box -3 -3 3 3
use M3_M2  M3_M2_7950
timestamp 1745462530
transform 1 0 1084 0 1 2705
box -3 -3 3 3
use M3_M2  M3_M2_7951
timestamp 1745462530
transform 1 0 1108 0 1 1865
box -3 -3 3 3
use M3_M2  M3_M2_7952
timestamp 1745462530
transform 1 0 1092 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_7953
timestamp 1745462530
transform 1 0 1012 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_7954
timestamp 1745462530
transform 1 0 1012 0 1 1865
box -3 -3 3 3
use M3_M2  M3_M2_7955
timestamp 1745462530
transform 1 0 1188 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_7956
timestamp 1745462530
transform 1 0 1164 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_7957
timestamp 1745462530
transform 1 0 2516 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_7958
timestamp 1745462530
transform 1 0 2468 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_7959
timestamp 1745462530
transform 1 0 2500 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_7960
timestamp 1745462530
transform 1 0 2452 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_7961
timestamp 1745462530
transform 1 0 3068 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_7962
timestamp 1745462530
transform 1 0 2516 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_7963
timestamp 1745462530
transform 1 0 3468 0 1 2045
box -3 -3 3 3
use M3_M2  M3_M2_7964
timestamp 1745462530
transform 1 0 3092 0 1 2055
box -3 -3 3 3
use M3_M2  M3_M2_7965
timestamp 1745462530
transform 1 0 3108 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_7966
timestamp 1745462530
transform 1 0 3068 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_7967
timestamp 1745462530
transform 1 0 3068 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_7968
timestamp 1745462530
transform 1 0 3044 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_7969
timestamp 1745462530
transform 1 0 3588 0 1 2045
box -3 -3 3 3
use M3_M2  M3_M2_7970
timestamp 1745462530
transform 1 0 3500 0 1 2045
box -3 -3 3 3
use M3_M2  M3_M2_7971
timestamp 1745462530
transform 1 0 3316 0 1 2045
box -3 -3 3 3
use M3_M2  M3_M2_7972
timestamp 1745462530
transform 1 0 2516 0 1 2045
box -3 -3 3 3
use M3_M2  M3_M2_7973
timestamp 1745462530
transform 1 0 2476 0 1 845
box -3 -3 3 3
use M3_M2  M3_M2_7974
timestamp 1745462530
transform 1 0 2452 0 1 845
box -3 -3 3 3
use M3_M2  M3_M2_7975
timestamp 1745462530
transform 1 0 2484 0 1 1005
box -3 -3 3 3
use M3_M2  M3_M2_7976
timestamp 1745462530
transform 1 0 2388 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_7977
timestamp 1745462530
transform 1 0 2484 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_7978
timestamp 1745462530
transform 1 0 2388 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_7979
timestamp 1745462530
transform 1 0 2476 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_7980
timestamp 1745462530
transform 1 0 2444 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_7981
timestamp 1745462530
transform 1 0 2532 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_7982
timestamp 1745462530
transform 1 0 2492 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_7983
timestamp 1745462530
transform 1 0 2628 0 1 3085
box -3 -3 3 3
use M3_M2  M3_M2_7984
timestamp 1745462530
transform 1 0 2588 0 1 3085
box -3 -3 3 3
use M3_M2  M3_M2_7985
timestamp 1745462530
transform 1 0 4060 0 1 1845
box -3 -3 3 3
use M3_M2  M3_M2_7986
timestamp 1745462530
transform 1 0 2356 0 1 1845
box -3 -3 3 3
use M3_M2  M3_M2_7987
timestamp 1745462530
transform 1 0 2332 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_7988
timestamp 1745462530
transform 1 0 1676 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_7989
timestamp 1745462530
transform 1 0 1644 0 1 1885
box -3 -3 3 3
use M3_M2  M3_M2_7990
timestamp 1745462530
transform 1 0 1084 0 1 1885
box -3 -3 3 3
use M3_M2  M3_M2_7991
timestamp 1745462530
transform 1 0 1636 0 1 1855
box -3 -3 3 3
use M3_M2  M3_M2_7992
timestamp 1745462530
transform 1 0 548 0 1 2155
box -3 -3 3 3
use M3_M2  M3_M2_7993
timestamp 1745462530
transform 1 0 508 0 1 2155
box -3 -3 3 3
use M3_M2  M3_M2_7994
timestamp 1745462530
transform 1 0 500 0 1 1855
box -3 -3 3 3
use M3_M2  M3_M2_7995
timestamp 1745462530
transform 1 0 1748 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_7996
timestamp 1745462530
transform 1 0 1708 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_7997
timestamp 1745462530
transform 1 0 1708 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_7998
timestamp 1745462530
transform 1 0 1676 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_7999
timestamp 1745462530
transform 1 0 1732 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_8000
timestamp 1745462530
transform 1 0 1708 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_8001
timestamp 1745462530
transform 1 0 1756 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_8002
timestamp 1745462530
transform 1 0 1716 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_8003
timestamp 1745462530
transform 1 0 580 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_8004
timestamp 1745462530
transform 1 0 524 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_8005
timestamp 1745462530
transform 1 0 660 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_8006
timestamp 1745462530
transform 1 0 564 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_8007
timestamp 1745462530
transform 1 0 1004 0 1 2155
box -3 -3 3 3
use M3_M2  M3_M2_8008
timestamp 1745462530
transform 1 0 924 0 1 2155
box -3 -3 3 3
use M3_M2  M3_M2_8009
timestamp 1745462530
transform 1 0 4036 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_8010
timestamp 1745462530
transform 1 0 3996 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_8011
timestamp 1745462530
transform 1 0 4044 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_8012
timestamp 1745462530
transform 1 0 4004 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_8013
timestamp 1745462530
transform 1 0 3932 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_8014
timestamp 1745462530
transform 1 0 3924 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_8015
timestamp 1745462530
transform 1 0 4172 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_8016
timestamp 1745462530
transform 1 0 4148 0 1 2245
box -3 -3 3 3
use M3_M2  M3_M2_8017
timestamp 1745462530
transform 1 0 4084 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_8018
timestamp 1745462530
transform 1 0 4076 0 1 2245
box -3 -3 3 3
use M3_M2  M3_M2_8019
timestamp 1745462530
transform 1 0 4148 0 1 2545
box -3 -3 3 3
use M3_M2  M3_M2_8020
timestamp 1745462530
transform 1 0 4092 0 1 2545
box -3 -3 3 3
use M3_M2  M3_M2_8021
timestamp 1745462530
transform 1 0 4100 0 1 2565
box -3 -3 3 3
use M3_M2  M3_M2_8022
timestamp 1745462530
transform 1 0 4020 0 1 2565
box -3 -3 3 3
use M3_M2  M3_M2_8023
timestamp 1745462530
transform 1 0 4116 0 1 2355
box -3 -3 3 3
use M3_M2  M3_M2_8024
timestamp 1745462530
transform 1 0 4076 0 1 2355
box -3 -3 3 3
use M3_M2  M3_M2_8025
timestamp 1745462530
transform 1 0 4092 0 1 2335
box -3 -3 3 3
use M3_M2  M3_M2_8026
timestamp 1745462530
transform 1 0 3012 0 1 2325
box -3 -3 3 3
use M3_M2  M3_M2_8027
timestamp 1745462530
transform 1 0 4052 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_8028
timestamp 1745462530
transform 1 0 3948 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_8029
timestamp 1745462530
transform 1 0 4004 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_8030
timestamp 1745462530
transform 1 0 3932 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_8031
timestamp 1745462530
transform 1 0 3996 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_8032
timestamp 1745462530
transform 1 0 3916 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_8033
timestamp 1745462530
transform 1 0 3148 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_8034
timestamp 1745462530
transform 1 0 2292 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_8035
timestamp 1745462530
transform 1 0 2284 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_8036
timestamp 1745462530
transform 1 0 2012 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_8037
timestamp 1745462530
transform 1 0 2028 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_8038
timestamp 1745462530
transform 1 0 1988 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_8039
timestamp 1745462530
transform 1 0 2068 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_8040
timestamp 1745462530
transform 1 0 1996 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_8041
timestamp 1745462530
transform 1 0 2068 0 1 1455
box -3 -3 3 3
use M3_M2  M3_M2_8042
timestamp 1745462530
transform 1 0 1012 0 1 1455
box -3 -3 3 3
use M3_M2  M3_M2_8043
timestamp 1745462530
transform 1 0 2012 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_8044
timestamp 1745462530
transform 1 0 1980 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_8045
timestamp 1745462530
transform 1 0 1980 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_8046
timestamp 1745462530
transform 1 0 596 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_8047
timestamp 1745462530
transform 1 0 684 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_8048
timestamp 1745462530
transform 1 0 588 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_8049
timestamp 1745462530
transform 1 0 588 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_8050
timestamp 1745462530
transform 1 0 524 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_8051
timestamp 1745462530
transform 1 0 660 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_8052
timestamp 1745462530
transform 1 0 588 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_8053
timestamp 1745462530
transform 1 0 956 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_8054
timestamp 1745462530
transform 1 0 884 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_8055
timestamp 1745462530
transform 1 0 988 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_8056
timestamp 1745462530
transform 1 0 964 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_8057
timestamp 1745462530
transform 1 0 2124 0 1 2375
box -3 -3 3 3
use M3_M2  M3_M2_8058
timestamp 1745462530
transform 1 0 2044 0 1 2375
box -3 -3 3 3
use M3_M2  M3_M2_8059
timestamp 1745462530
transform 1 0 2060 0 1 2625
box -3 -3 3 3
use M3_M2  M3_M2_8060
timestamp 1745462530
transform 1 0 1964 0 1 2625
box -3 -3 3 3
use M3_M2  M3_M2_8061
timestamp 1745462530
transform 1 0 3180 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_8062
timestamp 1745462530
transform 1 0 3124 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_8063
timestamp 1745462530
transform 1 0 3180 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_8064
timestamp 1745462530
transform 1 0 3156 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_8065
timestamp 1745462530
transform 1 0 3140 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_8066
timestamp 1745462530
transform 1 0 3140 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_8067
timestamp 1745462530
transform 1 0 3092 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_8068
timestamp 1745462530
transform 1 0 3084 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_8069
timestamp 1745462530
transform 1 0 3948 0 1 2075
box -3 -3 3 3
use M3_M2  M3_M2_8070
timestamp 1745462530
transform 1 0 3612 0 1 2075
box -3 -3 3 3
use M3_M2  M3_M2_8071
timestamp 1745462530
transform 1 0 3604 0 1 1895
box -3 -3 3 3
use M3_M2  M3_M2_8072
timestamp 1745462530
transform 1 0 3180 0 1 1895
box -3 -3 3 3
use M3_M2  M3_M2_8073
timestamp 1745462530
transform 1 0 4020 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_8074
timestamp 1745462530
transform 1 0 3996 0 1 2165
box -3 -3 3 3
use M3_M2  M3_M2_8075
timestamp 1745462530
transform 1 0 3996 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_8076
timestamp 1745462530
transform 1 0 3964 0 1 2165
box -3 -3 3 3
use M3_M2  M3_M2_8077
timestamp 1745462530
transform 1 0 3980 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_8078
timestamp 1745462530
transform 1 0 3924 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_8079
timestamp 1745462530
transform 1 0 3956 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_8080
timestamp 1745462530
transform 1 0 3092 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_8081
timestamp 1745462530
transform 1 0 3132 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_8082
timestamp 1745462530
transform 1 0 3116 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_8083
timestamp 1745462530
transform 1 0 3180 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_8084
timestamp 1745462530
transform 1 0 3148 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_8085
timestamp 1745462530
transform 1 0 3140 0 1 865
box -3 -3 3 3
use M3_M2  M3_M2_8086
timestamp 1745462530
transform 1 0 2972 0 1 865
box -3 -3 3 3
use M3_M2  M3_M2_8087
timestamp 1745462530
transform 1 0 3132 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_8088
timestamp 1745462530
transform 1 0 3060 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_8089
timestamp 1745462530
transform 1 0 4060 0 1 1835
box -3 -3 3 3
use M3_M2  M3_M2_8090
timestamp 1745462530
transform 1 0 2292 0 1 1835
box -3 -3 3 3
use M3_M2  M3_M2_8091
timestamp 1745462530
transform 1 0 2300 0 1 1845
box -3 -3 3 3
use M3_M2  M3_M2_8092
timestamp 1745462530
transform 1 0 2044 0 1 1845
box -3 -3 3 3
use M3_M2  M3_M2_8093
timestamp 1745462530
transform 1 0 2044 0 1 1665
box -3 -3 3 3
use M3_M2  M3_M2_8094
timestamp 1745462530
transform 1 0 1804 0 1 1665
box -3 -3 3 3
use M3_M2  M3_M2_8095
timestamp 1745462530
transform 1 0 1756 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_8096
timestamp 1745462530
transform 1 0 988 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_8097
timestamp 1745462530
transform 1 0 1812 0 1 1895
box -3 -3 3 3
use M3_M2  M3_M2_8098
timestamp 1745462530
transform 1 0 692 0 1 1895
box -3 -3 3 3
use M3_M2  M3_M2_8099
timestamp 1745462530
transform 1 0 1796 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_8100
timestamp 1745462530
transform 1 0 1772 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_8101
timestamp 1745462530
transform 1 0 1836 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_8102
timestamp 1745462530
transform 1 0 1812 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_8103
timestamp 1745462530
transform 1 0 1804 0 1 645
box -3 -3 3 3
use M3_M2  M3_M2_8104
timestamp 1745462530
transform 1 0 1756 0 1 645
box -3 -3 3 3
use M3_M2  M3_M2_8105
timestamp 1745462530
transform 1 0 668 0 1 2005
box -3 -3 3 3
use M3_M2  M3_M2_8106
timestamp 1745462530
transform 1 0 628 0 1 2165
box -3 -3 3 3
use M3_M2  M3_M2_8107
timestamp 1745462530
transform 1 0 580 0 1 2005
box -3 -3 3 3
use M3_M2  M3_M2_8108
timestamp 1745462530
transform 1 0 572 0 1 2165
box -3 -3 3 3
use M3_M2  M3_M2_8109
timestamp 1745462530
transform 1 0 684 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_8110
timestamp 1745462530
transform 1 0 596 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_8111
timestamp 1745462530
transform 1 0 956 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_8112
timestamp 1745462530
transform 1 0 908 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_8113
timestamp 1745462530
transform 1 0 1020 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_8114
timestamp 1745462530
transform 1 0 940 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_8115
timestamp 1745462530
transform 1 0 4156 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_8116
timestamp 1745462530
transform 1 0 4156 0 1 1455
box -3 -3 3 3
use M3_M2  M3_M2_8117
timestamp 1745462530
transform 1 0 4052 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_8118
timestamp 1745462530
transform 1 0 4052 0 1 1455
box -3 -3 3 3
use M3_M2  M3_M2_8119
timestamp 1745462530
transform 1 0 4084 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_8120
timestamp 1745462530
transform 1 0 4052 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_8121
timestamp 1745462530
transform 1 0 3996 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_8122
timestamp 1745462530
transform 1 0 3988 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_8123
timestamp 1745462530
transform 1 0 4356 0 1 2325
box -3 -3 3 3
use M3_M2  M3_M2_8124
timestamp 1745462530
transform 1 0 4348 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_8125
timestamp 1745462530
transform 1 0 4092 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_8126
timestamp 1745462530
transform 1 0 4068 0 1 2325
box -3 -3 3 3
use M3_M2  M3_M2_8127
timestamp 1745462530
transform 1 0 4108 0 1 2385
box -3 -3 3 3
use M3_M2  M3_M2_8128
timestamp 1745462530
transform 1 0 4052 0 1 2385
box -3 -3 3 3
use M3_M2  M3_M2_8129
timestamp 1745462530
transform 1 0 4068 0 1 2425
box -3 -3 3 3
use M3_M2  M3_M2_8130
timestamp 1745462530
transform 1 0 4004 0 1 2425
box -3 -3 3 3
use M3_M2  M3_M2_8131
timestamp 1745462530
transform 1 0 4108 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_8132
timestamp 1745462530
transform 1 0 4068 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_8133
timestamp 1745462530
transform 1 0 4052 0 1 2365
box -3 -3 3 3
use M3_M2  M3_M2_8134
timestamp 1745462530
transform 1 0 2948 0 1 2365
box -3 -3 3 3
use M3_M2  M3_M2_8135
timestamp 1745462530
transform 1 0 4084 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_8136
timestamp 1745462530
transform 1 0 3996 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_8137
timestamp 1745462530
transform 1 0 4060 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_8138
timestamp 1745462530
transform 1 0 3908 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_8139
timestamp 1745462530
transform 1 0 3900 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_8140
timestamp 1745462530
transform 1 0 3868 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_8141
timestamp 1745462530
transform 1 0 4060 0 1 1015
box -3 -3 3 3
use M3_M2  M3_M2_8142
timestamp 1745462530
transform 1 0 4036 0 1 1285
box -3 -3 3 3
use M3_M2  M3_M2_8143
timestamp 1745462530
transform 1 0 4036 0 1 1015
box -3 -3 3 3
use M3_M2  M3_M2_8144
timestamp 1745462530
transform 1 0 4012 0 1 1285
box -3 -3 3 3
use M3_M2  M3_M2_8145
timestamp 1745462530
transform 1 0 4028 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_8146
timestamp 1745462530
transform 1 0 3972 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_8147
timestamp 1745462530
transform 1 0 2276 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_8148
timestamp 1745462530
transform 1 0 1572 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_8149
timestamp 1745462530
transform 1 0 1636 0 1 2065
box -3 -3 3 3
use M3_M2  M3_M2_8150
timestamp 1745462530
transform 1 0 1572 0 1 2065
box -3 -3 3 3
use M3_M2  M3_M2_8151
timestamp 1745462530
transform 1 0 1572 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_8152
timestamp 1745462530
transform 1 0 1548 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_8153
timestamp 1745462530
transform 1 0 1548 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_8154
timestamp 1745462530
transform 1 0 1516 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_8155
timestamp 1745462530
transform 1 0 1588 0 1 1655
box -3 -3 3 3
use M3_M2  M3_M2_8156
timestamp 1745462530
transform 1 0 1012 0 1 1655
box -3 -3 3 3
use M3_M2  M3_M2_8157
timestamp 1745462530
transform 1 0 1580 0 1 1665
box -3 -3 3 3
use M3_M2  M3_M2_8158
timestamp 1745462530
transform 1 0 828 0 1 1665
box -3 -3 3 3
use M3_M2  M3_M2_8159
timestamp 1745462530
transform 1 0 828 0 1 1285
box -3 -3 3 3
use M3_M2  M3_M2_8160
timestamp 1745462530
transform 1 0 660 0 1 1285
box -3 -3 3 3
use M3_M2  M3_M2_8161
timestamp 1745462530
transform 1 0 644 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_8162
timestamp 1745462530
transform 1 0 580 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_8163
timestamp 1745462530
transform 1 0 596 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_8164
timestamp 1745462530
transform 1 0 524 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_8165
timestamp 1745462530
transform 1 0 1020 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_8166
timestamp 1745462530
transform 1 0 996 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_8167
timestamp 1745462530
transform 1 0 1652 0 1 2705
box -3 -3 3 3
use M3_M2  M3_M2_8168
timestamp 1745462530
transform 1 0 1596 0 1 2695
box -3 -3 3 3
use M3_M2  M3_M2_8169
timestamp 1745462530
transform 1 0 1644 0 1 2635
box -3 -3 3 3
use M3_M2  M3_M2_8170
timestamp 1745462530
transform 1 0 1620 0 1 2635
box -3 -3 3 3
use M3_M2  M3_M2_8171
timestamp 1745462530
transform 1 0 1652 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_8172
timestamp 1745462530
transform 1 0 1620 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_8173
timestamp 1745462530
transform 1 0 1612 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_8174
timestamp 1745462530
transform 1 0 1580 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_8175
timestamp 1745462530
transform 1 0 1604 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_8176
timestamp 1745462530
transform 1 0 1572 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_8177
timestamp 1745462530
transform 1 0 2612 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_8178
timestamp 1745462530
transform 1 0 2300 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_8179
timestamp 1745462530
transform 1 0 2916 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_8180
timestamp 1745462530
transform 1 0 2292 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_8181
timestamp 1745462530
transform 1 0 3268 0 1 1485
box -3 -3 3 3
use M3_M2  M3_M2_8182
timestamp 1745462530
transform 1 0 2948 0 1 1485
box -3 -3 3 3
use M3_M2  M3_M2_8183
timestamp 1745462530
transform 1 0 3404 0 1 1495
box -3 -3 3 3
use M3_M2  M3_M2_8184
timestamp 1745462530
transform 1 0 3300 0 1 1495
box -3 -3 3 3
use M3_M2  M3_M2_8185
timestamp 1745462530
transform 1 0 3212 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_8186
timestamp 1745462530
transform 1 0 2636 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_8187
timestamp 1745462530
transform 1 0 2636 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_8188
timestamp 1745462530
transform 1 0 2604 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_8189
timestamp 1745462530
transform 1 0 2276 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_8190
timestamp 1745462530
transform 1 0 2244 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_8191
timestamp 1745462530
transform 1 0 2276 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_8192
timestamp 1745462530
transform 1 0 2212 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_8193
timestamp 1745462530
transform 1 0 2340 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_8194
timestamp 1745462530
transform 1 0 2260 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_8195
timestamp 1745462530
transform 1 0 2348 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_8196
timestamp 1745462530
transform 1 0 2308 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_8197
timestamp 1745462530
transform 1 0 2412 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_8198
timestamp 1745462530
transform 1 0 2388 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_8199
timestamp 1745462530
transform 1 0 3148 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_8200
timestamp 1745462530
transform 1 0 2348 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_8201
timestamp 1745462530
transform 1 0 2324 0 1 1665
box -3 -3 3 3
use M3_M2  M3_M2_8202
timestamp 1745462530
transform 1 0 1460 0 1 1645
box -3 -3 3 3
use M3_M2  M3_M2_8203
timestamp 1745462530
transform 1 0 1436 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_8204
timestamp 1745462530
transform 1 0 1076 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_8205
timestamp 1745462530
transform 1 0 1452 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_8206
timestamp 1745462530
transform 1 0 1396 0 1 1835
box -3 -3 3 3
use M3_M2  M3_M2_8207
timestamp 1745462530
transform 1 0 1396 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_8208
timestamp 1745462530
transform 1 0 1076 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_8209
timestamp 1745462530
transform 1 0 1076 0 1 1835
box -3 -3 3 3
use M3_M2  M3_M2_8210
timestamp 1745462530
transform 1 0 1044 0 1 2125
box -3 -3 3 3
use M3_M2  M3_M2_8211
timestamp 1745462530
transform 1 0 1044 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_8212
timestamp 1745462530
transform 1 0 836 0 1 2175
box -3 -3 3 3
use M3_M2  M3_M2_8213
timestamp 1745462530
transform 1 0 836 0 1 2125
box -3 -3 3 3
use M3_M2  M3_M2_8214
timestamp 1745462530
transform 1 0 716 0 1 2275
box -3 -3 3 3
use M3_M2  M3_M2_8215
timestamp 1745462530
transform 1 0 676 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_8216
timestamp 1745462530
transform 1 0 676 0 1 2175
box -3 -3 3 3
use M3_M2  M3_M2_8217
timestamp 1745462530
transform 1 0 652 0 1 2275
box -3 -3 3 3
use M3_M2  M3_M2_8218
timestamp 1745462530
transform 1 0 652 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_8219
timestamp 1745462530
transform 1 0 1524 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_8220
timestamp 1745462530
transform 1 0 1508 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_8221
timestamp 1745462530
transform 1 0 1532 0 1 675
box -3 -3 3 3
use M3_M2  M3_M2_8222
timestamp 1745462530
transform 1 0 1380 0 1 675
box -3 -3 3 3
use M3_M2  M3_M2_8223
timestamp 1745462530
transform 1 0 1532 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_8224
timestamp 1745462530
transform 1 0 1492 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_8225
timestamp 1745462530
transform 1 0 668 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_8226
timestamp 1745462530
transform 1 0 644 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_8227
timestamp 1745462530
transform 1 0 700 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_8228
timestamp 1745462530
transform 1 0 644 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_8229
timestamp 1745462530
transform 1 0 676 0 1 2765
box -3 -3 3 3
use M3_M2  M3_M2_8230
timestamp 1745462530
transform 1 0 596 0 1 2765
box -3 -3 3 3
use M3_M2  M3_M2_8231
timestamp 1745462530
transform 1 0 1076 0 1 1815
box -3 -3 3 3
use M3_M2  M3_M2_8232
timestamp 1745462530
transform 1 0 1060 0 1 1815
box -3 -3 3 3
use M3_M2  M3_M2_8233
timestamp 1745462530
transform 1 0 3180 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_8234
timestamp 1745462530
transform 1 0 3132 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_8235
timestamp 1745462530
transform 1 0 3100 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_8236
timestamp 1745462530
transform 1 0 3092 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_8237
timestamp 1745462530
transform 1 0 3204 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_8238
timestamp 1745462530
transform 1 0 3164 0 1 1335
box -3 -3 3 3
use M3_M2  M3_M2_8239
timestamp 1745462530
transform 1 0 3164 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_8240
timestamp 1745462530
transform 1 0 3060 0 1 1335
box -3 -3 3 3
use M3_M2  M3_M2_8241
timestamp 1745462530
transform 1 0 3156 0 1 2135
box -3 -3 3 3
use M3_M2  M3_M2_8242
timestamp 1745462530
transform 1 0 3108 0 1 2135
box -3 -3 3 3
use M3_M2  M3_M2_8243
timestamp 1745462530
transform 1 0 3236 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_8244
timestamp 1745462530
transform 1 0 3132 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_8245
timestamp 1745462530
transform 1 0 3148 0 1 2545
box -3 -3 3 3
use M3_M2  M3_M2_8246
timestamp 1745462530
transform 1 0 3092 0 1 2545
box -3 -3 3 3
use M3_M2  M3_M2_8247
timestamp 1745462530
transform 1 0 3220 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_8248
timestamp 1745462530
transform 1 0 3172 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_8249
timestamp 1745462530
transform 1 0 3172 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_8250
timestamp 1745462530
transform 1 0 3148 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_8251
timestamp 1745462530
transform 1 0 3180 0 1 2065
box -3 -3 3 3
use M3_M2  M3_M2_8252
timestamp 1745462530
transform 1 0 2780 0 1 2065
box -3 -3 3 3
use M3_M2  M3_M2_8253
timestamp 1745462530
transform 1 0 3324 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_8254
timestamp 1745462530
transform 1 0 3204 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_8255
timestamp 1745462530
transform 1 0 3228 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_8256
timestamp 1745462530
transform 1 0 3116 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_8257
timestamp 1745462530
transform 1 0 3308 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_8258
timestamp 1745462530
transform 1 0 3220 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_8259
timestamp 1745462530
transform 1 0 3260 0 1 1055
box -3 -3 3 3
use M3_M2  M3_M2_8260
timestamp 1745462530
transform 1 0 3260 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_8261
timestamp 1745462530
transform 1 0 3220 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_8262
timestamp 1745462530
transform 1 0 3196 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_8263
timestamp 1745462530
transform 1 0 3196 0 1 1055
box -3 -3 3 3
use M3_M2  M3_M2_8264
timestamp 1745462530
transform 1 0 3148 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_8265
timestamp 1745462530
transform 1 0 3172 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_8266
timestamp 1745462530
transform 1 0 3148 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_8267
timestamp 1745462530
transform 1 0 3052 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_8268
timestamp 1745462530
transform 1 0 2372 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_8269
timestamp 1745462530
transform 1 0 2356 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_8270
timestamp 1745462530
transform 1 0 1172 0 1 1615
box -3 -3 3 3
use M3_M2  M3_M2_8271
timestamp 1745462530
transform 1 0 1244 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_8272
timestamp 1745462530
transform 1 0 1148 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_8273
timestamp 1745462530
transform 1 0 1356 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_8274
timestamp 1745462530
transform 1 0 1324 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_8275
timestamp 1745462530
transform 1 0 1324 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_8276
timestamp 1745462530
transform 1 0 1156 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_8277
timestamp 1745462530
transform 1 0 1188 0 1 1415
box -3 -3 3 3
use M3_M2  M3_M2_8278
timestamp 1745462530
transform 1 0 1100 0 1 1415
box -3 -3 3 3
use M3_M2  M3_M2_8279
timestamp 1745462530
transform 1 0 1172 0 1 1535
box -3 -3 3 3
use M3_M2  M3_M2_8280
timestamp 1745462530
transform 1 0 652 0 1 1535
box -3 -3 3 3
use M3_M2  M3_M2_8281
timestamp 1745462530
transform 1 0 652 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_8282
timestamp 1745462530
transform 1 0 628 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_8283
timestamp 1745462530
transform 1 0 652 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_8284
timestamp 1745462530
transform 1 0 588 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_8285
timestamp 1745462530
transform 1 0 644 0 1 685
box -3 -3 3 3
use M3_M2  M3_M2_8286
timestamp 1745462530
transform 1 0 588 0 1 685
box -3 -3 3 3
use M3_M2  M3_M2_8287
timestamp 1745462530
transform 1 0 1076 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_8288
timestamp 1745462530
transform 1 0 1052 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_8289
timestamp 1745462530
transform 1 0 1364 0 1 2685
box -3 -3 3 3
use M3_M2  M3_M2_8290
timestamp 1745462530
transform 1 0 1308 0 1 2685
box -3 -3 3 3
use M3_M2  M3_M2_8291
timestamp 1745462530
transform 1 0 1396 0 1 2805
box -3 -3 3 3
use M3_M2  M3_M2_8292
timestamp 1745462530
transform 1 0 1356 0 1 2805
box -3 -3 3 3
use M3_M2  M3_M2_8293
timestamp 1745462530
transform 1 0 1324 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_8294
timestamp 1745462530
transform 1 0 1260 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_8295
timestamp 1745462530
transform 1 0 3068 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_8296
timestamp 1745462530
transform 1 0 3012 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_8297
timestamp 1745462530
transform 1 0 2996 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_8298
timestamp 1745462530
transform 1 0 2996 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_8299
timestamp 1745462530
transform 1 0 3068 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_8300
timestamp 1745462530
transform 1 0 2972 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_8301
timestamp 1745462530
transform 1 0 3188 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_8302
timestamp 1745462530
transform 1 0 3108 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_8303
timestamp 1745462530
transform 1 0 3132 0 1 1495
box -3 -3 3 3
use M3_M2  M3_M2_8304
timestamp 1745462530
transform 1 0 3092 0 1 1495
box -3 -3 3 3
use M3_M2  M3_M2_8305
timestamp 1745462530
transform 1 0 3324 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_8306
timestamp 1745462530
transform 1 0 3212 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_8307
timestamp 1745462530
transform 1 0 3124 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_8308
timestamp 1745462530
transform 1 0 2956 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_8309
timestamp 1745462530
transform 1 0 3036 0 1 645
box -3 -3 3 3
use M3_M2  M3_M2_8310
timestamp 1745462530
transform 1 0 2916 0 1 645
box -3 -3 3 3
use M3_M2  M3_M2_8311
timestamp 1745462530
transform 1 0 2492 0 1 2475
box -3 -3 3 3
use M3_M2  M3_M2_8312
timestamp 1745462530
transform 1 0 2476 0 1 2475
box -3 -3 3 3
use M3_M2  M3_M2_8313
timestamp 1745462530
transform 1 0 2476 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_8314
timestamp 1745462530
transform 1 0 2428 0 1 2475
box -3 -3 3 3
use M3_M2  M3_M2_8315
timestamp 1745462530
transform 1 0 2412 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_8316
timestamp 1745462530
transform 1 0 3116 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_8317
timestamp 1745462530
transform 1 0 3116 0 1 1085
box -3 -3 3 3
use M3_M2  M3_M2_8318
timestamp 1745462530
transform 1 0 3116 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_8319
timestamp 1745462530
transform 1 0 3092 0 1 1085
box -3 -3 3 3
use M3_M2  M3_M2_8320
timestamp 1745462530
transform 1 0 3092 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_8321
timestamp 1745462530
transform 1 0 3052 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_8322
timestamp 1745462530
transform 1 0 3060 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_8323
timestamp 1745462530
transform 1 0 3044 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_8324
timestamp 1745462530
transform 1 0 2228 0 1 3835
box -3 -3 3 3
use M3_M2  M3_M2_8325
timestamp 1745462530
transform 1 0 2172 0 1 3835
box -3 -3 3 3
use M3_M2  M3_M2_8326
timestamp 1745462530
transform 1 0 2380 0 1 3795
box -3 -3 3 3
use M3_M2  M3_M2_8327
timestamp 1745462530
transform 1 0 2212 0 1 3795
box -3 -3 3 3
use M3_M2  M3_M2_8328
timestamp 1745462530
transform 1 0 2724 0 1 3825
box -3 -3 3 3
use M3_M2  M3_M2_8329
timestamp 1745462530
transform 1 0 2356 0 1 3825
box -3 -3 3 3
use M3_M2  M3_M2_8330
timestamp 1745462530
transform 1 0 2004 0 1 3045
box -3 -3 3 3
use M3_M2  M3_M2_8331
timestamp 1745462530
transform 1 0 1668 0 1 3145
box -3 -3 3 3
use M3_M2  M3_M2_8332
timestamp 1745462530
transform 1 0 1668 0 1 3045
box -3 -3 3 3
use M3_M2  M3_M2_8333
timestamp 1745462530
transform 1 0 1588 0 1 3145
box -3 -3 3 3
use M3_M2  M3_M2_8334
timestamp 1745462530
transform 1 0 1164 0 1 3145
box -3 -3 3 3
use M3_M2  M3_M2_8335
timestamp 1745462530
transform 1 0 2308 0 1 3845
box -3 -3 3 3
use M3_M2  M3_M2_8336
timestamp 1745462530
transform 1 0 2132 0 1 3845
box -3 -3 3 3
use M3_M2  M3_M2_8337
timestamp 1745462530
transform 1 0 3460 0 1 3835
box -3 -3 3 3
use M3_M2  M3_M2_8338
timestamp 1745462530
transform 1 0 2340 0 1 3835
box -3 -3 3 3
use M3_M2  M3_M2_8339
timestamp 1745462530
transform 1 0 3580 0 1 3745
box -3 -3 3 3
use M3_M2  M3_M2_8340
timestamp 1745462530
transform 1 0 3468 0 1 3745
box -3 -3 3 3
use M3_M2  M3_M2_8341
timestamp 1745462530
transform 1 0 3444 0 1 3895
box -3 -3 3 3
use M3_M2  M3_M2_8342
timestamp 1745462530
transform 1 0 3260 0 1 3895
box -3 -3 3 3
use M3_M2  M3_M2_8343
timestamp 1745462530
transform 1 0 3916 0 1 3805
box -3 -3 3 3
use M3_M2  M3_M2_8344
timestamp 1745462530
transform 1 0 3452 0 1 3805
box -3 -3 3 3
use M3_M2  M3_M2_8345
timestamp 1745462530
transform 1 0 3988 0 1 3785
box -3 -3 3 3
use M3_M2  M3_M2_8346
timestamp 1745462530
transform 1 0 3940 0 1 3785
box -3 -3 3 3
use M3_M2  M3_M2_8347
timestamp 1745462530
transform 1 0 4044 0 1 3795
box -3 -3 3 3
use M3_M2  M3_M2_8348
timestamp 1745462530
transform 1 0 3964 0 1 3795
box -3 -3 3 3
use M3_M2  M3_M2_8349
timestamp 1745462530
transform 1 0 4276 0 1 3885
box -3 -3 3 3
use M3_M2  M3_M2_8350
timestamp 1745462530
transform 1 0 4276 0 1 3765
box -3 -3 3 3
use M3_M2  M3_M2_8351
timestamp 1745462530
transform 1 0 4236 0 1 3765
box -3 -3 3 3
use M3_M2  M3_M2_8352
timestamp 1745462530
transform 1 0 4228 0 1 3635
box -3 -3 3 3
use M3_M2  M3_M2_8353
timestamp 1745462530
transform 1 0 4164 0 1 3885
box -3 -3 3 3
use M3_M2  M3_M2_8354
timestamp 1745462530
transform 1 0 4164 0 1 3635
box -3 -3 3 3
use M3_M2  M3_M2_8355
timestamp 1745462530
transform 1 0 4028 0 1 4025
box -3 -3 3 3
use M3_M2  M3_M2_8356
timestamp 1745462530
transform 1 0 4028 0 1 3885
box -3 -3 3 3
use M3_M2  M3_M2_8357
timestamp 1745462530
transform 1 0 1780 0 1 4025
box -3 -3 3 3
use M3_M2  M3_M2_8358
timestamp 1745462530
transform 1 0 1772 0 1 3845
box -3 -3 3 3
use M3_M2  M3_M2_8359
timestamp 1745462530
transform 1 0 1732 0 1 3775
box -3 -3 3 3
use M3_M2  M3_M2_8360
timestamp 1745462530
transform 1 0 1660 0 1 3845
box -3 -3 3 3
use M3_M2  M3_M2_8361
timestamp 1745462530
transform 1 0 1660 0 1 3775
box -3 -3 3 3
use M3_M2  M3_M2_8362
timestamp 1745462530
transform 1 0 4252 0 1 3665
box -3 -3 3 3
use M3_M2  M3_M2_8363
timestamp 1745462530
transform 1 0 4180 0 1 3955
box -3 -3 3 3
use M3_M2  M3_M2_8364
timestamp 1745462530
transform 1 0 4172 0 1 3665
box -3 -3 3 3
use M3_M2  M3_M2_8365
timestamp 1745462530
transform 1 0 4052 0 1 4085
box -3 -3 3 3
use M3_M2  M3_M2_8366
timestamp 1745462530
transform 1 0 4052 0 1 3955
box -3 -3 3 3
use M3_M2  M3_M2_8367
timestamp 1745462530
transform 1 0 4028 0 1 4085
box -3 -3 3 3
use M3_M2  M3_M2_8368
timestamp 1745462530
transform 1 0 4020 0 1 4245
box -3 -3 3 3
use M3_M2  M3_M2_8369
timestamp 1745462530
transform 1 0 2108 0 1 4245
box -3 -3 3 3
use M3_M2  M3_M2_8370
timestamp 1745462530
transform 1 0 2108 0 1 4045
box -3 -3 3 3
use M3_M2  M3_M2_8371
timestamp 1745462530
transform 1 0 1852 0 1 4045
box -3 -3 3 3
use M3_M2  M3_M2_8372
timestamp 1745462530
transform 1 0 4084 0 1 3855
box -3 -3 3 3
use M3_M2  M3_M2_8373
timestamp 1745462530
transform 1 0 4084 0 1 3715
box -3 -3 3 3
use M3_M2  M3_M2_8374
timestamp 1745462530
transform 1 0 4052 0 1 3715
box -3 -3 3 3
use M3_M2  M3_M2_8375
timestamp 1745462530
transform 1 0 3980 0 1 3845
box -3 -3 3 3
use M3_M2  M3_M2_8376
timestamp 1745462530
transform 1 0 3812 0 1 3945
box -3 -3 3 3
use M3_M2  M3_M2_8377
timestamp 1745462530
transform 1 0 3812 0 1 3845
box -3 -3 3 3
use M3_M2  M3_M2_8378
timestamp 1745462530
transform 1 0 3156 0 1 4065
box -3 -3 3 3
use M3_M2  M3_M2_8379
timestamp 1745462530
transform 1 0 3156 0 1 3945
box -3 -3 3 3
use M3_M2  M3_M2_8380
timestamp 1745462530
transform 1 0 2852 0 1 4195
box -3 -3 3 3
use M3_M2  M3_M2_8381
timestamp 1745462530
transform 1 0 2852 0 1 4065
box -3 -3 3 3
use M3_M2  M3_M2_8382
timestamp 1745462530
transform 1 0 2604 0 1 4195
box -3 -3 3 3
use M3_M2  M3_M2_8383
timestamp 1745462530
transform 1 0 2596 0 1 4085
box -3 -3 3 3
use M3_M2  M3_M2_8384
timestamp 1745462530
transform 1 0 2532 0 1 4085
box -3 -3 3 3
use M3_M2  M3_M2_8385
timestamp 1745462530
transform 1 0 2532 0 1 3995
box -3 -3 3 3
use M3_M2  M3_M2_8386
timestamp 1745462530
transform 1 0 2532 0 1 3935
box -3 -3 3 3
use M3_M2  M3_M2_8387
timestamp 1745462530
transform 1 0 2500 0 1 3935
box -3 -3 3 3
use M3_M2  M3_M2_8388
timestamp 1745462530
transform 1 0 1924 0 1 3995
box -3 -3 3 3
use M3_M2  M3_M2_8389
timestamp 1745462530
transform 1 0 4124 0 1 3685
box -3 -3 3 3
use M3_M2  M3_M2_8390
timestamp 1745462530
transform 1 0 4100 0 1 3825
box -3 -3 3 3
use M3_M2  M3_M2_8391
timestamp 1745462530
transform 1 0 4068 0 1 3685
box -3 -3 3 3
use M3_M2  M3_M2_8392
timestamp 1745462530
transform 1 0 3996 0 1 3855
box -3 -3 3 3
use M3_M2  M3_M2_8393
timestamp 1745462530
transform 1 0 3996 0 1 3825
box -3 -3 3 3
use M3_M2  M3_M2_8394
timestamp 1745462530
transform 1 0 3948 0 1 3855
box -3 -3 3 3
use M3_M2  M3_M2_8395
timestamp 1745462530
transform 1 0 3948 0 1 3685
box -3 -3 3 3
use M3_M2  M3_M2_8396
timestamp 1745462530
transform 1 0 2484 0 1 3855
box -3 -3 3 3
use M3_M2  M3_M2_8397
timestamp 1745462530
transform 1 0 1708 0 1 3855
box -3 -3 3 3
use M3_M2  M3_M2_8398
timestamp 1745462530
transform 1 0 1708 0 1 3755
box -3 -3 3 3
use M3_M2  M3_M2_8399
timestamp 1745462530
transform 1 0 1684 0 1 3755
box -3 -3 3 3
use M3_M2  M3_M2_8400
timestamp 1745462530
transform 1 0 1908 0 1 3165
box -3 -3 3 3
use M3_M2  M3_M2_8401
timestamp 1745462530
transform 1 0 1868 0 1 3165
box -3 -3 3 3
use M3_M2  M3_M2_8402
timestamp 1745462530
transform 1 0 1652 0 1 3165
box -3 -3 3 3
use M3_M2  M3_M2_8403
timestamp 1745462530
transform 1 0 1636 0 1 3165
box -3 -3 3 3
use M3_M2  M3_M2_8404
timestamp 1745462530
transform 1 0 3564 0 1 3755
box -3 -3 3 3
use M3_M2  M3_M2_8405
timestamp 1745462530
transform 1 0 3540 0 1 3755
box -3 -3 3 3
use M3_M2  M3_M2_8406
timestamp 1745462530
transform 1 0 3996 0 1 3705
box -3 -3 3 3
use M3_M2  M3_M2_8407
timestamp 1745462530
transform 1 0 3580 0 1 3705
box -3 -3 3 3
use M3_M2  M3_M2_8408
timestamp 1745462530
transform 1 0 4164 0 1 3705
box -3 -3 3 3
use M3_M2  M3_M2_8409
timestamp 1745462530
transform 1 0 4044 0 1 3705
box -3 -3 3 3
use M3_M2  M3_M2_8410
timestamp 1745462530
transform 1 0 3124 0 1 3105
box -3 -3 3 3
use M3_M2  M3_M2_8411
timestamp 1745462530
transform 1 0 1708 0 1 3105
box -3 -3 3 3
use M3_M2  M3_M2_8412
timestamp 1745462530
transform 1 0 2276 0 1 3865
box -3 -3 3 3
use M3_M2  M3_M2_8413
timestamp 1745462530
transform 1 0 2164 0 1 3865
box -3 -3 3 3
use M3_M2  M3_M2_8414
timestamp 1745462530
transform 1 0 2164 0 1 3795
box -3 -3 3 3
use M3_M2  M3_M2_8415
timestamp 1745462530
transform 1 0 2100 0 1 3795
box -3 -3 3 3
use M3_M2  M3_M2_8416
timestamp 1745462530
transform 1 0 1956 0 1 3175
box -3 -3 3 3
use M3_M2  M3_M2_8417
timestamp 1745462530
transform 1 0 1612 0 1 3185
box -3 -3 3 3
use M3_M2  M3_M2_8418
timestamp 1745462530
transform 1 0 2084 0 1 3665
box -3 -3 3 3
use M3_M2  M3_M2_8419
timestamp 1745462530
transform 1 0 1716 0 1 3665
box -3 -3 3 3
use M3_M2  M3_M2_8420
timestamp 1745462530
transform 1 0 2116 0 1 3705
box -3 -3 3 3
use M3_M2  M3_M2_8421
timestamp 1745462530
transform 1 0 2068 0 1 3705
box -3 -3 3 3
use M3_M2  M3_M2_8422
timestamp 1745462530
transform 1 0 2356 0 1 4045
box -3 -3 3 3
use M3_M2  M3_M2_8423
timestamp 1745462530
transform 1 0 2332 0 1 4045
box -3 -3 3 3
use M3_M2  M3_M2_8424
timestamp 1745462530
transform 1 0 2164 0 1 3545
box -3 -3 3 3
use M3_M2  M3_M2_8425
timestamp 1745462530
transform 1 0 1532 0 1 3525
box -3 -3 3 3
use M3_M2  M3_M2_8426
timestamp 1745462530
transform 1 0 1492 0 1 3525
box -3 -3 3 3
use M3_M2  M3_M2_8427
timestamp 1745462530
transform 1 0 2052 0 1 3825
box -3 -3 3 3
use M3_M2  M3_M2_8428
timestamp 1745462530
transform 1 0 1740 0 1 3825
box -3 -3 3 3
use M3_M2  M3_M2_8429
timestamp 1745462530
transform 1 0 2084 0 1 3835
box -3 -3 3 3
use M3_M2  M3_M2_8430
timestamp 1745462530
transform 1 0 2036 0 1 3835
box -3 -3 3 3
use M3_M2  M3_M2_8431
timestamp 1745462530
transform 1 0 2236 0 1 4065
box -3 -3 3 3
use M3_M2  M3_M2_8432
timestamp 1745462530
transform 1 0 2116 0 1 4065
box -3 -3 3 3
use M3_M2  M3_M2_8433
timestamp 1745462530
transform 1 0 2172 0 1 4045
box -3 -3 3 3
use M3_M2  M3_M2_8434
timestamp 1745462530
transform 1 0 2124 0 1 4045
box -3 -3 3 3
use M3_M2  M3_M2_8435
timestamp 1745462530
transform 1 0 2764 0 1 3815
box -3 -3 3 3
use M3_M2  M3_M2_8436
timestamp 1745462530
transform 1 0 2716 0 1 3815
box -3 -3 3 3
use M3_M2  M3_M2_8437
timestamp 1745462530
transform 1 0 3524 0 1 3675
box -3 -3 3 3
use M3_M2  M3_M2_8438
timestamp 1745462530
transform 1 0 2732 0 1 3675
box -3 -3 3 3
use M3_M2  M3_M2_8439
timestamp 1745462530
transform 1 0 3596 0 1 3775
box -3 -3 3 3
use M3_M2  M3_M2_8440
timestamp 1745462530
transform 1 0 3516 0 1 3775
box -3 -3 3 3
use M3_M2  M3_M2_8441
timestamp 1745462530
transform 1 0 3540 0 1 3955
box -3 -3 3 3
use M3_M2  M3_M2_8442
timestamp 1745462530
transform 1 0 3508 0 1 3955
box -3 -3 3 3
use M3_M2  M3_M2_8443
timestamp 1745462530
transform 1 0 3516 0 1 3915
box -3 -3 3 3
use M3_M2  M3_M2_8444
timestamp 1745462530
transform 1 0 3484 0 1 3915
box -3 -3 3 3
use M3_M2  M3_M2_8445
timestamp 1745462530
transform 1 0 4116 0 1 3875
box -3 -3 3 3
use M3_M2  M3_M2_8446
timestamp 1745462530
transform 1 0 3524 0 1 3875
box -3 -3 3 3
use M3_M2  M3_M2_8447
timestamp 1745462530
transform 1 0 1620 0 1 3325
box -3 -3 3 3
use M3_M2  M3_M2_8448
timestamp 1745462530
transform 1 0 1564 0 1 3405
box -3 -3 3 3
use M3_M2  M3_M2_8449
timestamp 1745462530
transform 1 0 1564 0 1 3325
box -3 -3 3 3
use M3_M2  M3_M2_8450
timestamp 1745462530
transform 1 0 1500 0 1 3405
box -3 -3 3 3
use M3_M2  M3_M2_8451
timestamp 1745462530
transform 1 0 3580 0 1 3795
box -3 -3 3 3
use M3_M2  M3_M2_8452
timestamp 1745462530
transform 1 0 3492 0 1 3795
box -3 -3 3 3
use M3_M2  M3_M2_8453
timestamp 1745462530
transform 1 0 4212 0 1 3755
box -3 -3 3 3
use M3_M2  M3_M2_8454
timestamp 1745462530
transform 1 0 3588 0 1 3755
box -3 -3 3 3
use M3_M2  M3_M2_8455
timestamp 1745462530
transform 1 0 4204 0 1 3745
box -3 -3 3 3
use M3_M2  M3_M2_8456
timestamp 1745462530
transform 1 0 4116 0 1 3745
box -3 -3 3 3
use M3_M2  M3_M2_8457
timestamp 1745462530
transform 1 0 4244 0 1 3695
box -3 -3 3 3
use M3_M2  M3_M2_8458
timestamp 1745462530
transform 1 0 4228 0 1 3695
box -3 -3 3 3
use M3_M2  M3_M2_8459
timestamp 1745462530
transform 1 0 2732 0 1 3845
box -3 -3 3 3
use M3_M2  M3_M2_8460
timestamp 1745462530
transform 1 0 2668 0 1 3845
box -3 -3 3 3
use M3_M2  M3_M2_8461
timestamp 1745462530
transform 1 0 2660 0 1 3865
box -3 -3 3 3
use M3_M2  M3_M2_8462
timestamp 1745462530
transform 1 0 2524 0 1 3865
box -3 -3 3 3
use M3_M2  M3_M2_8463
timestamp 1745462530
transform 1 0 2492 0 1 3815
box -3 -3 3 3
use M3_M2  M3_M2_8464
timestamp 1745462530
transform 1 0 1844 0 1 3845
box -3 -3 3 3
use M3_M2  M3_M2_8465
timestamp 1745462530
transform 1 0 2556 0 1 3845
box -3 -3 3 3
use M3_M2  M3_M2_8466
timestamp 1745462530
transform 1 0 2532 0 1 3845
box -3 -3 3 3
use M3_M2  M3_M2_8467
timestamp 1745462530
transform 1 0 2724 0 1 3995
box -3 -3 3 3
use M3_M2  M3_M2_8468
timestamp 1745462530
transform 1 0 2684 0 1 3995
box -3 -3 3 3
use M3_M2  M3_M2_8469
timestamp 1745462530
transform 1 0 2780 0 1 3935
box -3 -3 3 3
use M3_M2  M3_M2_8470
timestamp 1745462530
transform 1 0 2756 0 1 3935
box -3 -3 3 3
use M3_M2  M3_M2_8471
timestamp 1745462530
transform 1 0 3004 0 1 3865
box -3 -3 3 3
use M3_M2  M3_M2_8472
timestamp 1745462530
transform 1 0 2740 0 1 3865
box -3 -3 3 3
use M3_M2  M3_M2_8473
timestamp 1745462530
transform 1 0 2748 0 1 3795
box -3 -3 3 3
use M3_M2  M3_M2_8474
timestamp 1745462530
transform 1 0 2612 0 1 3795
box -3 -3 3 3
use M3_M2  M3_M2_8475
timestamp 1745462530
transform 1 0 2572 0 1 3785
box -3 -3 3 3
use M3_M2  M3_M2_8476
timestamp 1745462530
transform 1 0 1796 0 1 3785
box -3 -3 3 3
use M3_M2  M3_M2_8477
timestamp 1745462530
transform 1 0 1908 0 1 3705
box -3 -3 3 3
use M3_M2  M3_M2_8478
timestamp 1745462530
transform 1 0 1860 0 1 3705
box -3 -3 3 3
use M3_M2  M3_M2_8479
timestamp 1745462530
transform 1 0 1652 0 1 3705
box -3 -3 3 3
use M3_M2  M3_M2_8480
timestamp 1745462530
transform 1 0 1756 0 1 3725
box -3 -3 3 3
use M3_M2  M3_M2_8481
timestamp 1745462530
transform 1 0 1628 0 1 3725
box -3 -3 3 3
use M3_M2  M3_M2_8482
timestamp 1745462530
transform 1 0 3052 0 1 3955
box -3 -3 3 3
use M3_M2  M3_M2_8483
timestamp 1745462530
transform 1 0 2996 0 1 3955
box -3 -3 3 3
use M3_M2  M3_M2_8484
timestamp 1745462530
transform 1 0 3052 0 1 3935
box -3 -3 3 3
use M3_M2  M3_M2_8485
timestamp 1745462530
transform 1 0 3012 0 1 3935
box -3 -3 3 3
use M3_M2  M3_M2_8486
timestamp 1745462530
transform 1 0 1820 0 1 3685
box -3 -3 3 3
use M3_M2  M3_M2_8487
timestamp 1745462530
transform 1 0 1612 0 1 3675
box -3 -3 3 3
use M3_M2  M3_M2_8488
timestamp 1745462530
transform 1 0 1444 0 1 3675
box -3 -3 3 3
use M3_M2  M3_M2_8489
timestamp 1745462530
transform 1 0 2068 0 1 3555
box -3 -3 3 3
use M3_M2  M3_M2_8490
timestamp 1745462530
transform 1 0 1572 0 1 3555
box -3 -3 3 3
use M3_M2  M3_M2_8491
timestamp 1745462530
transform 1 0 1108 0 1 3365
box -3 -3 3 3
use M3_M2  M3_M2_8492
timestamp 1745462530
transform 1 0 1068 0 1 3555
box -3 -3 3 3
use M3_M2  M3_M2_8493
timestamp 1745462530
transform 1 0 988 0 1 3555
box -3 -3 3 3
use M3_M2  M3_M2_8494
timestamp 1745462530
transform 1 0 844 0 1 3555
box -3 -3 3 3
use M3_M2  M3_M2_8495
timestamp 1745462530
transform 1 0 836 0 1 3365
box -3 -3 3 3
use M3_M2  M3_M2_8496
timestamp 1745462530
transform 1 0 948 0 1 3505
box -3 -3 3 3
use M3_M2  M3_M2_8497
timestamp 1745462530
transform 1 0 844 0 1 3505
box -3 -3 3 3
use M3_M2  M3_M2_8498
timestamp 1745462530
transform 1 0 1020 0 1 3635
box -3 -3 3 3
use M3_M2  M3_M2_8499
timestamp 1745462530
transform 1 0 964 0 1 3635
box -3 -3 3 3
use M3_M2  M3_M2_8500
timestamp 1745462530
transform 1 0 1140 0 1 3535
box -3 -3 3 3
use M3_M2  M3_M2_8501
timestamp 1745462530
transform 1 0 1116 0 1 3535
box -3 -3 3 3
use M3_M2  M3_M2_8502
timestamp 1745462530
transform 1 0 1604 0 1 3105
box -3 -3 3 3
use M3_M2  M3_M2_8503
timestamp 1745462530
transform 1 0 1564 0 1 3175
box -3 -3 3 3
use M3_M2  M3_M2_8504
timestamp 1745462530
transform 1 0 1564 0 1 3105
box -3 -3 3 3
use M3_M2  M3_M2_8505
timestamp 1745462530
transform 1 0 1428 0 1 3175
box -3 -3 3 3
use M3_M2  M3_M2_8506
timestamp 1745462530
transform 1 0 1372 0 1 3175
box -3 -3 3 3
use M3_M2  M3_M2_8507
timestamp 1745462530
transform 1 0 1364 0 1 3195
box -3 -3 3 3
use M3_M2  M3_M2_8508
timestamp 1745462530
transform 1 0 1316 0 1 3195
box -3 -3 3 3
use M3_M2  M3_M2_8509
timestamp 1745462530
transform 1 0 1636 0 1 3155
box -3 -3 3 3
use M3_M2  M3_M2_8510
timestamp 1745462530
transform 1 0 1636 0 1 3115
box -3 -3 3 3
use M3_M2  M3_M2_8511
timestamp 1745462530
transform 1 0 1596 0 1 3115
box -3 -3 3 3
use M3_M2  M3_M2_8512
timestamp 1745462530
transform 1 0 1356 0 1 3155
box -3 -3 3 3
use M3_M2  M3_M2_8513
timestamp 1745462530
transform 1 0 1340 0 1 3155
box -3 -3 3 3
use M3_M2  M3_M2_8514
timestamp 1745462530
transform 1 0 1860 0 1 2865
box -3 -3 3 3
use M3_M2  M3_M2_8515
timestamp 1745462530
transform 1 0 1796 0 1 2865
box -3 -3 3 3
use M3_M2  M3_M2_8516
timestamp 1745462530
transform 1 0 1732 0 1 2865
box -3 -3 3 3
use M3_M2  M3_M2_8517
timestamp 1745462530
transform 1 0 1636 0 1 2785
box -3 -3 3 3
use M3_M2  M3_M2_8518
timestamp 1745462530
transform 1 0 1580 0 1 2785
box -3 -3 3 3
use M3_M2  M3_M2_8519
timestamp 1745462530
transform 1 0 1572 0 1 2865
box -3 -3 3 3
use M3_M2  M3_M2_8520
timestamp 1745462530
transform 1 0 1492 0 1 2865
box -3 -3 3 3
use M3_M2  M3_M2_8521
timestamp 1745462530
transform 1 0 1492 0 1 2845
box -3 -3 3 3
use M3_M2  M3_M2_8522
timestamp 1745462530
transform 1 0 1292 0 1 2845
box -3 -3 3 3
use M3_M2  M3_M2_8523
timestamp 1745462530
transform 1 0 1292 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_8524
timestamp 1745462530
transform 1 0 1236 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_8525
timestamp 1745462530
transform 1 0 2452 0 1 2165
box -3 -3 3 3
use M3_M2  M3_M2_8526
timestamp 1745462530
transform 1 0 1836 0 1 2165
box -3 -3 3 3
use M3_M2  M3_M2_8527
timestamp 1745462530
transform 1 0 1972 0 1 2215
box -3 -3 3 3
use M3_M2  M3_M2_8528
timestamp 1745462530
transform 1 0 1892 0 1 2215
box -3 -3 3 3
use M3_M2  M3_M2_8529
timestamp 1745462530
transform 1 0 1692 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_8530
timestamp 1745462530
transform 1 0 1636 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_8531
timestamp 1745462530
transform 1 0 1548 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_8532
timestamp 1745462530
transform 1 0 1476 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_8533
timestamp 1745462530
transform 1 0 1468 0 1 2165
box -3 -3 3 3
use M3_M2  M3_M2_8534
timestamp 1745462530
transform 1 0 1276 0 1 2165
box -3 -3 3 3
use M3_M2  M3_M2_8535
timestamp 1745462530
transform 1 0 1244 0 1 2165
box -3 -3 3 3
use M3_M2  M3_M2_8536
timestamp 1745462530
transform 1 0 1884 0 1 2585
box -3 -3 3 3
use M3_M2  M3_M2_8537
timestamp 1745462530
transform 1 0 1820 0 1 2635
box -3 -3 3 3
use M3_M2  M3_M2_8538
timestamp 1745462530
transform 1 0 1812 0 1 2585
box -3 -3 3 3
use M3_M2  M3_M2_8539
timestamp 1745462530
transform 1 0 1668 0 1 2755
box -3 -3 3 3
use M3_M2  M3_M2_8540
timestamp 1745462530
transform 1 0 1660 0 1 2635
box -3 -3 3 3
use M3_M2  M3_M2_8541
timestamp 1745462530
transform 1 0 1540 0 1 2565
box -3 -3 3 3
use M3_M2  M3_M2_8542
timestamp 1745462530
transform 1 0 1484 0 1 2565
box -3 -3 3 3
use M3_M2  M3_M2_8543
timestamp 1745462530
transform 1 0 1452 0 1 2755
box -3 -3 3 3
use M3_M2  M3_M2_8544
timestamp 1745462530
transform 1 0 1452 0 1 2565
box -3 -3 3 3
use M3_M2  M3_M2_8545
timestamp 1745462530
transform 1 0 1268 0 1 2755
box -3 -3 3 3
use M3_M2  M3_M2_8546
timestamp 1745462530
transform 1 0 1220 0 1 2755
box -3 -3 3 3
use M3_M2  M3_M2_8547
timestamp 1745462530
transform 1 0 1852 0 1 2055
box -3 -3 3 3
use M3_M2  M3_M2_8548
timestamp 1745462530
transform 1 0 1812 0 1 2055
box -3 -3 3 3
use M3_M2  M3_M2_8549
timestamp 1745462530
transform 1 0 1604 0 1 2055
box -3 -3 3 3
use M3_M2  M3_M2_8550
timestamp 1745462530
transform 1 0 1604 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_8551
timestamp 1745462530
transform 1 0 1444 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_8552
timestamp 1745462530
transform 1 0 1420 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_8553
timestamp 1745462530
transform 1 0 1244 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_8554
timestamp 1745462530
transform 1 0 1796 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_8555
timestamp 1745462530
transform 1 0 1732 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_8556
timestamp 1745462530
transform 1 0 1540 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_8557
timestamp 1745462530
transform 1 0 1404 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_8558
timestamp 1745462530
transform 1 0 1340 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_8559
timestamp 1745462530
transform 1 0 1260 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_8560
timestamp 1745462530
transform 1 0 1228 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_8561
timestamp 1745462530
transform 1 0 1796 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_8562
timestamp 1745462530
transform 1 0 1740 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_8563
timestamp 1745462530
transform 1 0 1580 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_8564
timestamp 1745462530
transform 1 0 1492 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_8565
timestamp 1745462530
transform 1 0 1348 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_8566
timestamp 1745462530
transform 1 0 1252 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_8567
timestamp 1745462530
transform 1 0 1180 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_8568
timestamp 1745462530
transform 1 0 1012 0 1 2865
box -3 -3 3 3
use M3_M2  M3_M2_8569
timestamp 1745462530
transform 1 0 852 0 1 2945
box -3 -3 3 3
use M3_M2  M3_M2_8570
timestamp 1745462530
transform 1 0 852 0 1 2865
box -3 -3 3 3
use M3_M2  M3_M2_8571
timestamp 1745462530
transform 1 0 772 0 1 2945
box -3 -3 3 3
use M3_M2  M3_M2_8572
timestamp 1745462530
transform 1 0 444 0 1 2775
box -3 -3 3 3
use M3_M2  M3_M2_8573
timestamp 1745462530
transform 1 0 404 0 1 2945
box -3 -3 3 3
use M3_M2  M3_M2_8574
timestamp 1745462530
transform 1 0 404 0 1 2775
box -3 -3 3 3
use M3_M2  M3_M2_8575
timestamp 1745462530
transform 1 0 332 0 1 2775
box -3 -3 3 3
use M3_M2  M3_M2_8576
timestamp 1745462530
transform 1 0 284 0 1 2775
box -3 -3 3 3
use M3_M2  M3_M2_8577
timestamp 1745462530
transform 1 0 796 0 1 2655
box -3 -3 3 3
use M3_M2  M3_M2_8578
timestamp 1745462530
transform 1 0 764 0 1 2475
box -3 -3 3 3
use M3_M2  M3_M2_8579
timestamp 1745462530
transform 1 0 716 0 1 2655
box -3 -3 3 3
use M3_M2  M3_M2_8580
timestamp 1745462530
transform 1 0 700 0 1 2865
box -3 -3 3 3
use M3_M2  M3_M2_8581
timestamp 1745462530
transform 1 0 604 0 1 2475
box -3 -3 3 3
use M3_M2  M3_M2_8582
timestamp 1745462530
transform 1 0 596 0 1 2705
box -3 -3 3 3
use M3_M2  M3_M2_8583
timestamp 1745462530
transform 1 0 556 0 1 2705
box -3 -3 3 3
use M3_M2  M3_M2_8584
timestamp 1745462530
transform 1 0 548 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_8585
timestamp 1745462530
transform 1 0 524 0 1 2475
box -3 -3 3 3
use M3_M2  M3_M2_8586
timestamp 1745462530
transform 1 0 508 0 1 2865
box -3 -3 3 3
use M3_M2  M3_M2_8587
timestamp 1745462530
transform 1 0 508 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_8588
timestamp 1745462530
transform 1 0 540 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_8589
timestamp 1745462530
transform 1 0 460 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_8590
timestamp 1745462530
transform 1 0 444 0 1 2615
box -3 -3 3 3
use M3_M2  M3_M2_8591
timestamp 1745462530
transform 1 0 444 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_8592
timestamp 1745462530
transform 1 0 348 0 1 2615
box -3 -3 3 3
use M3_M2  M3_M2_8593
timestamp 1745462530
transform 1 0 308 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_8594
timestamp 1745462530
transform 1 0 260 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_8595
timestamp 1745462530
transform 1 0 236 0 1 2615
box -3 -3 3 3
use M3_M2  M3_M2_8596
timestamp 1745462530
transform 1 0 972 0 1 2935
box -3 -3 3 3
use M3_M2  M3_M2_8597
timestamp 1745462530
transform 1 0 924 0 1 2935
box -3 -3 3 3
use M3_M2  M3_M2_8598
timestamp 1745462530
transform 1 0 476 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_8599
timestamp 1745462530
transform 1 0 412 0 1 2435
box -3 -3 3 3
use M3_M2  M3_M2_8600
timestamp 1745462530
transform 1 0 372 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_8601
timestamp 1745462530
transform 1 0 340 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_8602
timestamp 1745462530
transform 1 0 292 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_8603
timestamp 1745462530
transform 1 0 236 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_8604
timestamp 1745462530
transform 1 0 228 0 1 2435
box -3 -3 3 3
use M3_M2  M3_M2_8605
timestamp 1745462530
transform 1 0 180 0 1 2435
box -3 -3 3 3
use M3_M2  M3_M2_8606
timestamp 1745462530
transform 1 0 556 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_8607
timestamp 1745462530
transform 1 0 444 0 1 2185
box -3 -3 3 3
use M3_M2  M3_M2_8608
timestamp 1745462530
transform 1 0 444 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_8609
timestamp 1745462530
transform 1 0 404 0 1 1975
box -3 -3 3 3
use M3_M2  M3_M2_8610
timestamp 1745462530
transform 1 0 340 0 1 1975
box -3 -3 3 3
use M3_M2  M3_M2_8611
timestamp 1745462530
transform 1 0 268 0 1 2175
box -3 -3 3 3
use M3_M2  M3_M2_8612
timestamp 1745462530
transform 1 0 236 0 1 1975
box -3 -3 3 3
use M3_M2  M3_M2_8613
timestamp 1745462530
transform 1 0 204 0 1 2175
box -3 -3 3 3
use M3_M2  M3_M2_8614
timestamp 1745462530
transform 1 0 196 0 1 1975
box -3 -3 3 3
use M3_M2  M3_M2_8615
timestamp 1745462530
transform 1 0 676 0 1 2015
box -3 -3 3 3
use M3_M2  M3_M2_8616
timestamp 1745462530
transform 1 0 396 0 1 2015
box -3 -3 3 3
use M3_M2  M3_M2_8617
timestamp 1745462530
transform 1 0 396 0 1 1835
box -3 -3 3 3
use M3_M2  M3_M2_8618
timestamp 1745462530
transform 1 0 316 0 1 1835
box -3 -3 3 3
use M3_M2  M3_M2_8619
timestamp 1745462530
transform 1 0 244 0 1 1835
box -3 -3 3 3
use M3_M2  M3_M2_8620
timestamp 1745462530
transform 1 0 740 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_8621
timestamp 1745462530
transform 1 0 708 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_8622
timestamp 1745462530
transform 1 0 708 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_8623
timestamp 1745462530
transform 1 0 620 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_8624
timestamp 1745462530
transform 1 0 596 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_8625
timestamp 1745462530
transform 1 0 564 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_8626
timestamp 1745462530
transform 1 0 500 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_8627
timestamp 1745462530
transform 1 0 508 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_8628
timestamp 1745462530
transform 1 0 452 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_8629
timestamp 1745462530
transform 1 0 388 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_8630
timestamp 1745462530
transform 1 0 324 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_8631
timestamp 1745462530
transform 1 0 284 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_8632
timestamp 1745462530
transform 1 0 212 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_8633
timestamp 1745462530
transform 1 0 452 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_8634
timestamp 1745462530
transform 1 0 396 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_8635
timestamp 1745462530
transform 1 0 388 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_8636
timestamp 1745462530
transform 1 0 260 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_8637
timestamp 1745462530
transform 1 0 444 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_8638
timestamp 1745462530
transform 1 0 420 0 1 215
box -3 -3 3 3
use M3_M2  M3_M2_8639
timestamp 1745462530
transform 1 0 332 0 1 215
box -3 -3 3 3
use M3_M2  M3_M2_8640
timestamp 1745462530
transform 1 0 268 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_8641
timestamp 1745462530
transform 1 0 268 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_8642
timestamp 1745462530
transform 1 0 268 0 1 205
box -3 -3 3 3
use M3_M2  M3_M2_8643
timestamp 1745462530
transform 1 0 252 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_8644
timestamp 1745462530
transform 1 0 220 0 1 205
box -3 -3 3 3
use M3_M2  M3_M2_8645
timestamp 1745462530
transform 1 0 500 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_8646
timestamp 1745462530
transform 1 0 484 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_8647
timestamp 1745462530
transform 1 0 444 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_8648
timestamp 1745462530
transform 1 0 420 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_8649
timestamp 1745462530
transform 1 0 340 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_8650
timestamp 1745462530
transform 1 0 260 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_8651
timestamp 1745462530
transform 1 0 228 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_8652
timestamp 1745462530
transform 1 0 724 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_8653
timestamp 1745462530
transform 1 0 700 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_8654
timestamp 1745462530
transform 1 0 692 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_8655
timestamp 1745462530
transform 1 0 660 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_8656
timestamp 1745462530
transform 1 0 644 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_8657
timestamp 1745462530
transform 1 0 556 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_8658
timestamp 1745462530
transform 1 0 556 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_8659
timestamp 1745462530
transform 1 0 948 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_8660
timestamp 1745462530
transform 1 0 924 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_8661
timestamp 1745462530
transform 1 0 924 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_8662
timestamp 1745462530
transform 1 0 908 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_8663
timestamp 1745462530
transform 1 0 892 0 1 215
box -3 -3 3 3
use M3_M2  M3_M2_8664
timestamp 1745462530
transform 1 0 884 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_8665
timestamp 1745462530
transform 1 0 884 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_8666
timestamp 1745462530
transform 1 0 860 0 1 325
box -3 -3 3 3
use M3_M2  M3_M2_8667
timestamp 1745462530
transform 1 0 836 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_8668
timestamp 1745462530
transform 1 0 820 0 1 215
box -3 -3 3 3
use M3_M2  M3_M2_8669
timestamp 1745462530
transform 1 0 812 0 1 325
box -3 -3 3 3
use M3_M2  M3_M2_8670
timestamp 1745462530
transform 1 0 1004 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_8671
timestamp 1745462530
transform 1 0 452 0 1 1285
box -3 -3 3 3
use M3_M2  M3_M2_8672
timestamp 1745462530
transform 1 0 452 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_8673
timestamp 1745462530
transform 1 0 380 0 1 1285
box -3 -3 3 3
use M3_M2  M3_M2_8674
timestamp 1745462530
transform 1 0 372 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_8675
timestamp 1745462530
transform 1 0 220 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_8676
timestamp 1745462530
transform 1 0 172 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_8677
timestamp 1745462530
transform 1 0 1076 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_8678
timestamp 1745462530
transform 1 0 940 0 1 1415
box -3 -3 3 3
use M3_M2  M3_M2_8679
timestamp 1745462530
transform 1 0 940 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_8680
timestamp 1745462530
transform 1 0 836 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_8681
timestamp 1745462530
transform 1 0 820 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_8682
timestamp 1745462530
transform 1 0 804 0 1 1415
box -3 -3 3 3
use M3_M2  M3_M2_8683
timestamp 1745462530
transform 1 0 740 0 1 1415
box -3 -3 3 3
use M3_M2  M3_M2_8684
timestamp 1745462530
transform 1 0 676 0 1 1415
box -3 -3 3 3
use M3_M2  M3_M2_8685
timestamp 1745462530
transform 1 0 1668 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_8686
timestamp 1745462530
transform 1 0 1588 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_8687
timestamp 1745462530
transform 1 0 1460 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_8688
timestamp 1745462530
transform 1 0 1148 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_8689
timestamp 1745462530
transform 1 0 1940 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_8690
timestamp 1745462530
transform 1 0 1852 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_8691
timestamp 1745462530
transform 1 0 1692 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_8692
timestamp 1745462530
transform 1 0 1452 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_8693
timestamp 1745462530
transform 1 0 1244 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_8694
timestamp 1745462530
transform 1 0 1172 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_8695
timestamp 1745462530
transform 1 0 1036 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_8696
timestamp 1745462530
transform 1 0 1908 0 1 205
box -3 -3 3 3
use M3_M2  M3_M2_8697
timestamp 1745462530
transform 1 0 1812 0 1 205
box -3 -3 3 3
use M3_M2  M3_M2_8698
timestamp 1745462530
transform 1 0 1676 0 1 205
box -3 -3 3 3
use M3_M2  M3_M2_8699
timestamp 1745462530
transform 1 0 1524 0 1 205
box -3 -3 3 3
use M3_M2  M3_M2_8700
timestamp 1745462530
transform 1 0 1468 0 1 205
box -3 -3 3 3
use M3_M2  M3_M2_8701
timestamp 1745462530
transform 1 0 1380 0 1 205
box -3 -3 3 3
use M3_M2  M3_M2_8702
timestamp 1745462530
transform 1 0 1908 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_8703
timestamp 1745462530
transform 1 0 1844 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_8704
timestamp 1745462530
transform 1 0 1764 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_8705
timestamp 1745462530
transform 1 0 1748 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_8706
timestamp 1745462530
transform 1 0 1588 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_8707
timestamp 1745462530
transform 1 0 1580 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_8708
timestamp 1745462530
transform 1 0 1436 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_8709
timestamp 1745462530
transform 1 0 1364 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_8710
timestamp 1745462530
transform 1 0 1276 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_8711
timestamp 1745462530
transform 1 0 2036 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_8712
timestamp 1745462530
transform 1 0 1916 0 1 335
box -3 -3 3 3
use M3_M2  M3_M2_8713
timestamp 1745462530
transform 1 0 1740 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_8714
timestamp 1745462530
transform 1 0 1524 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_8715
timestamp 1745462530
transform 1 0 1508 0 1 135
box -3 -3 3 3
use M3_M2  M3_M2_8716
timestamp 1745462530
transform 1 0 1428 0 1 135
box -3 -3 3 3
use M3_M2  M3_M2_8717
timestamp 1745462530
transform 1 0 1332 0 1 135
box -3 -3 3 3
use M3_M2  M3_M2_8718
timestamp 1745462530
transform 1 0 2020 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_8719
timestamp 1745462530
transform 1 0 1988 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_8720
timestamp 1745462530
transform 1 0 1940 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_8721
timestamp 1745462530
transform 1 0 1788 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_8722
timestamp 1745462530
transform 1 0 1588 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_8723
timestamp 1745462530
transform 1 0 1500 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_8724
timestamp 1745462530
transform 1 0 1396 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_8725
timestamp 1745462530
transform 1 0 1980 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_8726
timestamp 1745462530
transform 1 0 1972 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_8727
timestamp 1745462530
transform 1 0 1916 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_8728
timestamp 1745462530
transform 1 0 1916 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_8729
timestamp 1745462530
transform 1 0 1820 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_8730
timestamp 1745462530
transform 1 0 1620 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_8731
timestamp 1745462530
transform 1 0 1580 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_8732
timestamp 1745462530
transform 1 0 1556 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_8733
timestamp 1745462530
transform 1 0 1500 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_8734
timestamp 1745462530
transform 1 0 1500 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_8735
timestamp 1745462530
transform 1 0 1404 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_8736
timestamp 1745462530
transform 1 0 2020 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_8737
timestamp 1745462530
transform 1 0 1956 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_8738
timestamp 1745462530
transform 1 0 1908 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_8739
timestamp 1745462530
transform 1 0 1828 0 1 1375
box -3 -3 3 3
use M3_M2  M3_M2_8740
timestamp 1745462530
transform 1 0 1612 0 1 1375
box -3 -3 3 3
use M3_M2  M3_M2_8741
timestamp 1745462530
transform 1 0 1604 0 1 1335
box -3 -3 3 3
use M3_M2  M3_M2_8742
timestamp 1745462530
transform 1 0 1556 0 1 1335
box -3 -3 3 3
use M3_M2  M3_M2_8743
timestamp 1745462530
transform 1 0 1508 0 1 1335
box -3 -3 3 3
use M3_M2  M3_M2_8744
timestamp 1745462530
transform 1 0 2884 0 1 375
box -3 -3 3 3
use M3_M2  M3_M2_8745
timestamp 1745462530
transform 1 0 2812 0 1 375
box -3 -3 3 3
use M3_M2  M3_M2_8746
timestamp 1745462530
transform 1 0 2692 0 1 375
box -3 -3 3 3
use M3_M2  M3_M2_8747
timestamp 1745462530
transform 1 0 2564 0 1 375
box -3 -3 3 3
use M3_M2  M3_M2_8748
timestamp 1745462530
transform 1 0 2340 0 1 365
box -3 -3 3 3
use M3_M2  M3_M2_8749
timestamp 1745462530
transform 1 0 2324 0 1 375
box -3 -3 3 3
use M3_M2  M3_M2_8750
timestamp 1745462530
transform 1 0 2268 0 1 365
box -3 -3 3 3
use M3_M2  M3_M2_8751
timestamp 1745462530
transform 1 0 2228 0 1 365
box -3 -3 3 3
use M3_M2  M3_M2_8752
timestamp 1745462530
transform 1 0 3084 0 1 675
box -3 -3 3 3
use M3_M2  M3_M2_8753
timestamp 1745462530
transform 1 0 3060 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_8754
timestamp 1745462530
transform 1 0 3044 0 1 675
box -3 -3 3 3
use M3_M2  M3_M2_8755
timestamp 1745462530
transform 1 0 2764 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_8756
timestamp 1745462530
transform 1 0 2764 0 1 685
box -3 -3 3 3
use M3_M2  M3_M2_8757
timestamp 1745462530
transform 1 0 2700 0 1 685
box -3 -3 3 3
use M3_M2  M3_M2_8758
timestamp 1745462530
transform 1 0 2628 0 1 685
box -3 -3 3 3
use M3_M2  M3_M2_8759
timestamp 1745462530
transform 1 0 2300 0 1 685
box -3 -3 3 3
use M3_M2  M3_M2_8760
timestamp 1745462530
transform 1 0 2212 0 1 685
box -3 -3 3 3
use M3_M2  M3_M2_8761
timestamp 1745462530
transform 1 0 2828 0 1 235
box -3 -3 3 3
use M3_M2  M3_M2_8762
timestamp 1745462530
transform 1 0 2668 0 1 245
box -3 -3 3 3
use M3_M2  M3_M2_8763
timestamp 1745462530
transform 1 0 2628 0 1 245
box -3 -3 3 3
use M3_M2  M3_M2_8764
timestamp 1745462530
transform 1 0 2604 0 1 485
box -3 -3 3 3
use M3_M2  M3_M2_8765
timestamp 1745462530
transform 1 0 2572 0 1 485
box -3 -3 3 3
use M3_M2  M3_M2_8766
timestamp 1745462530
transform 1 0 2572 0 1 245
box -3 -3 3 3
use M3_M2  M3_M2_8767
timestamp 1745462530
transform 1 0 2532 0 1 245
box -3 -3 3 3
use M3_M2  M3_M2_8768
timestamp 1745462530
transform 1 0 2316 0 1 245
box -3 -3 3 3
use M3_M2  M3_M2_8769
timestamp 1745462530
transform 1 0 2316 0 1 205
box -3 -3 3 3
use M3_M2  M3_M2_8770
timestamp 1745462530
transform 1 0 2252 0 1 205
box -3 -3 3 3
use M3_M2  M3_M2_8771
timestamp 1745462530
transform 1 0 3020 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_8772
timestamp 1745462530
transform 1 0 2964 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_8773
timestamp 1745462530
transform 1 0 2788 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_8774
timestamp 1745462530
transform 1 0 2788 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_8775
timestamp 1745462530
transform 1 0 2692 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_8776
timestamp 1745462530
transform 1 0 2644 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_8777
timestamp 1745462530
transform 1 0 2316 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_8778
timestamp 1745462530
transform 1 0 2252 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_8779
timestamp 1745462530
transform 1 0 3124 0 1 325
box -3 -3 3 3
use M3_M2  M3_M2_8780
timestamp 1745462530
transform 1 0 3108 0 1 205
box -3 -3 3 3
use M3_M2  M3_M2_8781
timestamp 1745462530
transform 1 0 3052 0 1 205
box -3 -3 3 3
use M3_M2  M3_M2_8782
timestamp 1745462530
transform 1 0 2972 0 1 325
box -3 -3 3 3
use M3_M2  M3_M2_8783
timestamp 1745462530
transform 1 0 2652 0 1 335
box -3 -3 3 3
use M3_M2  M3_M2_8784
timestamp 1745462530
transform 1 0 2652 0 1 325
box -3 -3 3 3
use M3_M2  M3_M2_8785
timestamp 1745462530
transform 1 0 2620 0 1 335
box -3 -3 3 3
use M3_M2  M3_M2_8786
timestamp 1745462530
transform 1 0 2500 0 1 325
box -3 -3 3 3
use M3_M2  M3_M2_8787
timestamp 1745462530
transform 1 0 2468 0 1 335
box -3 -3 3 3
use M3_M2  M3_M2_8788
timestamp 1745462530
transform 1 0 2876 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_8789
timestamp 1745462530
transform 1 0 2764 0 1 1055
box -3 -3 3 3
use M3_M2  M3_M2_8790
timestamp 1745462530
transform 1 0 2764 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_8791
timestamp 1745462530
transform 1 0 2716 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_8792
timestamp 1745462530
transform 1 0 2716 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_8793
timestamp 1745462530
transform 1 0 2548 0 1 1055
box -3 -3 3 3
use M3_M2  M3_M2_8794
timestamp 1745462530
transform 1 0 2316 0 1 1055
box -3 -3 3 3
use M3_M2  M3_M2_8795
timestamp 1745462530
transform 1 0 2836 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_8796
timestamp 1745462530
transform 1 0 2668 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_8797
timestamp 1745462530
transform 1 0 2636 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_8798
timestamp 1745462530
transform 1 0 2596 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_8799
timestamp 1745462530
transform 1 0 2348 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_8800
timestamp 1745462530
transform 1 0 2292 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_8801
timestamp 1745462530
transform 1 0 2796 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_8802
timestamp 1745462530
transform 1 0 2772 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_8803
timestamp 1745462530
transform 1 0 2684 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_8804
timestamp 1745462530
transform 1 0 2604 0 1 1375
box -3 -3 3 3
use M3_M2  M3_M2_8805
timestamp 1745462530
transform 1 0 2580 0 1 1375
box -3 -3 3 3
use M3_M2  M3_M2_8806
timestamp 1745462530
transform 1 0 2372 0 1 1375
box -3 -3 3 3
use M3_M2  M3_M2_8807
timestamp 1745462530
transform 1 0 3396 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_8808
timestamp 1745462530
transform 1 0 3364 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_8809
timestamp 1745462530
transform 1 0 3356 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_8810
timestamp 1745462530
transform 1 0 3300 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_8811
timestamp 1745462530
transform 1 0 3300 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_8812
timestamp 1745462530
transform 1 0 3244 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_8813
timestamp 1745462530
transform 1 0 3180 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_8814
timestamp 1745462530
transform 1 0 3900 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_8815
timestamp 1745462530
transform 1 0 3828 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_8816
timestamp 1745462530
transform 1 0 3804 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_8817
timestamp 1745462530
transform 1 0 3756 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_8818
timestamp 1745462530
transform 1 0 3540 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_8819
timestamp 1745462530
transform 1 0 3372 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_8820
timestamp 1745462530
transform 1 0 4236 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_8821
timestamp 1745462530
transform 1 0 4236 0 1 235
box -3 -3 3 3
use M3_M2  M3_M2_8822
timestamp 1745462530
transform 1 0 4164 0 1 235
box -3 -3 3 3
use M3_M2  M3_M2_8823
timestamp 1745462530
transform 1 0 4092 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_8824
timestamp 1745462530
transform 1 0 4076 0 1 235
box -3 -3 3 3
use M3_M2  M3_M2_8825
timestamp 1745462530
transform 1 0 4028 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_8826
timestamp 1745462530
transform 1 0 3764 0 1 255
box -3 -3 3 3
use M3_M2  M3_M2_8827
timestamp 1745462530
transform 1 0 3620 0 1 255
box -3 -3 3 3
use M3_M2  M3_M2_8828
timestamp 1745462530
transform 1 0 4004 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_8829
timestamp 1745462530
transform 1 0 3796 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_8830
timestamp 1745462530
transform 1 0 3700 0 1 335
box -3 -3 3 3
use M3_M2  M3_M2_8831
timestamp 1745462530
transform 1 0 3660 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_8832
timestamp 1745462530
transform 1 0 3660 0 1 335
box -3 -3 3 3
use M3_M2  M3_M2_8833
timestamp 1745462530
transform 1 0 3572 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_8834
timestamp 1745462530
transform 1 0 3532 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_8835
timestamp 1745462530
transform 1 0 3532 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_8836
timestamp 1745462530
transform 1 0 3388 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_8837
timestamp 1745462530
transform 1 0 4340 0 1 605
box -3 -3 3 3
use M3_M2  M3_M2_8838
timestamp 1745462530
transform 1 0 4324 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_8839
timestamp 1745462530
transform 1 0 4268 0 1 405
box -3 -3 3 3
use M3_M2  M3_M2_8840
timestamp 1745462530
transform 1 0 4268 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_8841
timestamp 1745462530
transform 1 0 4236 0 1 605
box -3 -3 3 3
use M3_M2  M3_M2_8842
timestamp 1745462530
transform 1 0 4172 0 1 405
box -3 -3 3 3
use M3_M2  M3_M2_8843
timestamp 1745462530
transform 1 0 4164 0 1 605
box -3 -3 3 3
use M3_M2  M3_M2_8844
timestamp 1745462530
transform 1 0 4108 0 1 605
box -3 -3 3 3
use M3_M2  M3_M2_8845
timestamp 1745462530
transform 1 0 3820 0 1 605
box -3 -3 3 3
use M3_M2  M3_M2_8846
timestamp 1745462530
transform 1 0 4276 0 1 885
box -3 -3 3 3
use M3_M2  M3_M2_8847
timestamp 1745462530
transform 1 0 4212 0 1 885
box -3 -3 3 3
use M3_M2  M3_M2_8848
timestamp 1745462530
transform 1 0 4124 0 1 885
box -3 -3 3 3
use M3_M2  M3_M2_8849
timestamp 1745462530
transform 1 0 4044 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_8850
timestamp 1745462530
transform 1 0 3932 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_8851
timestamp 1745462530
transform 1 0 3292 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_8852
timestamp 1745462530
transform 1 0 4188 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_8853
timestamp 1745462530
transform 1 0 4148 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_8854
timestamp 1745462530
transform 1 0 4116 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_8855
timestamp 1745462530
transform 1 0 4084 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_8856
timestamp 1745462530
transform 1 0 3780 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_8857
timestamp 1745462530
transform 1 0 3780 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_8858
timestamp 1745462530
transform 1 0 3428 0 1 1015
box -3 -3 3 3
use M3_M2  M3_M2_8859
timestamp 1745462530
transform 1 0 3396 0 1 1015
box -3 -3 3 3
use M3_M2  M3_M2_8860
timestamp 1745462530
transform 1 0 3380 0 1 1015
box -3 -3 3 3
use M3_M2  M3_M2_8861
timestamp 1745462530
transform 1 0 3916 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_8862
timestamp 1745462530
transform 1 0 3860 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_8863
timestamp 1745462530
transform 1 0 3812 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_8864
timestamp 1745462530
transform 1 0 3772 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_8865
timestamp 1745462530
transform 1 0 3604 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_8866
timestamp 1745462530
transform 1 0 3460 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_8867
timestamp 1745462530
transform 1 0 3444 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_8868
timestamp 1745462530
transform 1 0 3364 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_8869
timestamp 1745462530
transform 1 0 4204 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_8870
timestamp 1745462530
transform 1 0 4204 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_8871
timestamp 1745462530
transform 1 0 4140 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_8872
timestamp 1745462530
transform 1 0 4116 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_8873
timestamp 1745462530
transform 1 0 4100 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_8874
timestamp 1745462530
transform 1 0 4076 0 1 1485
box -3 -3 3 3
use M3_M2  M3_M2_8875
timestamp 1745462530
transform 1 0 4076 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_8876
timestamp 1745462530
transform 1 0 4068 0 1 1535
box -3 -3 3 3
use M3_M2  M3_M2_8877
timestamp 1745462530
transform 1 0 3964 0 1 1535
box -3 -3 3 3
use M3_M2  M3_M2_8878
timestamp 1745462530
transform 1 0 3964 0 1 1485
box -3 -3 3 3
use M3_M2  M3_M2_8879
timestamp 1745462530
transform 1 0 3492 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_8880
timestamp 1745462530
transform 1 0 3836 0 1 1815
box -3 -3 3 3
use M3_M2  M3_M2_8881
timestamp 1745462530
transform 1 0 3820 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_8882
timestamp 1745462530
transform 1 0 3692 0 1 1815
box -3 -3 3 3
use M3_M2  M3_M2_8883
timestamp 1745462530
transform 1 0 3692 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_8884
timestamp 1745462530
transform 1 0 3692 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_8885
timestamp 1745462530
transform 1 0 3524 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_8886
timestamp 1745462530
transform 1 0 3492 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_8887
timestamp 1745462530
transform 1 0 4252 0 1 1775
box -3 -3 3 3
use M3_M2  M3_M2_8888
timestamp 1745462530
transform 1 0 4244 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_8889
timestamp 1745462530
transform 1 0 4236 0 1 1935
box -3 -3 3 3
use M3_M2  M3_M2_8890
timestamp 1745462530
transform 1 0 4228 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_8891
timestamp 1745462530
transform 1 0 4196 0 1 1935
box -3 -3 3 3
use M3_M2  M3_M2_8892
timestamp 1745462530
transform 1 0 4188 0 1 1775
box -3 -3 3 3
use M3_M2  M3_M2_8893
timestamp 1745462530
transform 1 0 4164 0 1 1935
box -3 -3 3 3
use M3_M2  M3_M2_8894
timestamp 1745462530
transform 1 0 4132 0 1 1935
box -3 -3 3 3
use M3_M2  M3_M2_8895
timestamp 1745462530
transform 1 0 4084 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_8896
timestamp 1745462530
transform 1 0 4028 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_8897
timestamp 1745462530
transform 1 0 3868 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_8898
timestamp 1745462530
transform 1 0 3852 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_8899
timestamp 1745462530
transform 1 0 3828 0 1 1655
box -3 -3 3 3
use M3_M2  M3_M2_8900
timestamp 1745462530
transform 1 0 3796 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_8901
timestamp 1745462530
transform 1 0 3708 0 1 2015
box -3 -3 3 3
use M3_M2  M3_M2_8902
timestamp 1745462530
transform 1 0 3668 0 1 1655
box -3 -3 3 3
use M3_M2  M3_M2_8903
timestamp 1745462530
transform 1 0 3668 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_8904
timestamp 1745462530
transform 1 0 3588 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_8905
timestamp 1745462530
transform 1 0 4332 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_8906
timestamp 1745462530
transform 1 0 4308 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_8907
timestamp 1745462530
transform 1 0 4252 0 1 1835
box -3 -3 3 3
use M3_M2  M3_M2_8908
timestamp 1745462530
transform 1 0 4236 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_8909
timestamp 1745462530
transform 1 0 4172 0 1 1615
box -3 -3 3 3
use M3_M2  M3_M2_8910
timestamp 1745462530
transform 1 0 4156 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_8911
timestamp 1745462530
transform 1 0 4148 0 1 1835
box -3 -3 3 3
use M3_M2  M3_M2_8912
timestamp 1745462530
transform 1 0 4148 0 1 1615
box -3 -3 3 3
use M3_M2  M3_M2_8913
timestamp 1745462530
transform 1 0 4148 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_8914
timestamp 1745462530
transform 1 0 4004 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_8915
timestamp 1745462530
transform 1 0 3980 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_8916
timestamp 1745462530
transform 1 0 3860 0 1 2015
box -3 -3 3 3
use M3_M2  M3_M2_8917
timestamp 1745462530
transform 1 0 3860 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_8918
timestamp 1745462530
transform 1 0 3852 0 1 2205
box -3 -3 3 3
use M3_M2  M3_M2_8919
timestamp 1745462530
transform 1 0 3732 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_8920
timestamp 1745462530
transform 1 0 3564 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_8921
timestamp 1745462530
transform 1 0 3564 0 1 2175
box -3 -3 3 3
use M3_M2  M3_M2_8922
timestamp 1745462530
transform 1 0 3340 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_8923
timestamp 1745462530
transform 1 0 3340 0 1 2175
box -3 -3 3 3
use M3_M2  M3_M2_8924
timestamp 1745462530
transform 1 0 3268 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_8925
timestamp 1745462530
transform 1 0 3212 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_8926
timestamp 1745462530
transform 1 0 3212 0 1 2135
box -3 -3 3 3
use M3_M2  M3_M2_8927
timestamp 1745462530
transform 1 0 3196 0 1 2135
box -3 -3 3 3
use M3_M2  M3_M2_8928
timestamp 1745462530
transform 1 0 3196 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_8929
timestamp 1745462530
transform 1 0 3100 0 1 2175
box -3 -3 3 3
use M3_M2  M3_M2_8930
timestamp 1745462530
transform 1 0 2980 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_8931
timestamp 1745462530
transform 1 0 2956 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_8932
timestamp 1745462530
transform 1 0 2844 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_8933
timestamp 1745462530
transform 1 0 2836 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_8934
timestamp 1745462530
transform 1 0 2828 0 1 2165
box -3 -3 3 3
use M3_M2  M3_M2_8935
timestamp 1745462530
transform 1 0 2804 0 1 2165
box -3 -3 3 3
use M3_M2  M3_M2_8936
timestamp 1745462530
transform 1 0 2780 0 1 2165
box -3 -3 3 3
use M3_M2  M3_M2_8937
timestamp 1745462530
transform 1 0 2764 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_8938
timestamp 1745462530
transform 1 0 2956 0 1 2135
box -3 -3 3 3
use M3_M2  M3_M2_8939
timestamp 1745462530
transform 1 0 2924 0 1 2135
box -3 -3 3 3
use M3_M2  M3_M2_8940
timestamp 1745462530
transform 1 0 2732 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_8941
timestamp 1745462530
transform 1 0 2692 0 1 2135
box -3 -3 3 3
use M3_M2  M3_M2_8942
timestamp 1745462530
transform 1 0 2668 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_8943
timestamp 1745462530
transform 1 0 2660 0 1 2135
box -3 -3 3 3
use M3_M2  M3_M2_8944
timestamp 1745462530
transform 1 0 2612 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_8945
timestamp 1745462530
transform 1 0 4180 0 1 2715
box -3 -3 3 3
use M3_M2  M3_M2_8946
timestamp 1745462530
transform 1 0 3836 0 1 2735
box -3 -3 3 3
use M3_M2  M3_M2_8947
timestamp 1745462530
transform 1 0 3748 0 1 2735
box -3 -3 3 3
use M3_M2  M3_M2_8948
timestamp 1745462530
transform 1 0 3644 0 1 2735
box -3 -3 3 3
use M3_M2  M3_M2_8949
timestamp 1745462530
transform 1 0 3420 0 1 2725
box -3 -3 3 3
use M3_M2  M3_M2_8950
timestamp 1745462530
transform 1 0 3268 0 1 2725
box -3 -3 3 3
use M3_M2  M3_M2_8951
timestamp 1745462530
transform 1 0 3076 0 1 2725
box -3 -3 3 3
use M3_M2  M3_M2_8952
timestamp 1745462530
transform 1 0 3916 0 1 3005
box -3 -3 3 3
use M3_M2  M3_M2_8953
timestamp 1745462530
transform 1 0 3884 0 1 3005
box -3 -3 3 3
use M3_M2  M3_M2_8954
timestamp 1745462530
transform 1 0 3748 0 1 3005
box -3 -3 3 3
use M3_M2  M3_M2_8955
timestamp 1745462530
transform 1 0 3684 0 1 3005
box -3 -3 3 3
use M3_M2  M3_M2_8956
timestamp 1745462530
transform 1 0 3236 0 1 3005
box -3 -3 3 3
use M3_M2  M3_M2_8957
timestamp 1745462530
transform 1 0 3212 0 1 2945
box -3 -3 3 3
use M3_M2  M3_M2_8958
timestamp 1745462530
transform 1 0 3100 0 1 2945
box -3 -3 3 3
use M3_M2  M3_M2_8959
timestamp 1745462530
transform 1 0 2996 0 1 2945
box -3 -3 3 3
use M3_M2  M3_M2_8960
timestamp 1745462530
transform 1 0 4148 0 1 2805
box -3 -3 3 3
use M3_M2  M3_M2_8961
timestamp 1745462530
transform 1 0 4060 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_8962
timestamp 1745462530
transform 1 0 3988 0 1 2785
box -3 -3 3 3
use M3_M2  M3_M2_8963
timestamp 1745462530
transform 1 0 3852 0 1 2785
box -3 -3 3 3
use M3_M2  M3_M2_8964
timestamp 1745462530
transform 1 0 3620 0 1 2785
box -3 -3 3 3
use M3_M2  M3_M2_8965
timestamp 1745462530
transform 1 0 3396 0 1 2805
box -3 -3 3 3
use M3_M2  M3_M2_8966
timestamp 1745462530
transform 1 0 3244 0 1 2785
box -3 -3 3 3
use M3_M2  M3_M2_8967
timestamp 1745462530
transform 1 0 3148 0 1 2785
box -3 -3 3 3
use M3_M2  M3_M2_8968
timestamp 1745462530
transform 1 0 4196 0 1 2965
box -3 -3 3 3
use M3_M2  M3_M2_8969
timestamp 1745462530
transform 1 0 4140 0 1 2965
box -3 -3 3 3
use M3_M2  M3_M2_8970
timestamp 1745462530
transform 1 0 3724 0 1 2965
box -3 -3 3 3
use M3_M2  M3_M2_8971
timestamp 1745462530
transform 1 0 3524 0 1 2965
box -3 -3 3 3
use M3_M2  M3_M2_8972
timestamp 1745462530
transform 1 0 3284 0 1 2975
box -3 -3 3 3
use M3_M2  M3_M2_8973
timestamp 1745462530
transform 1 0 3196 0 1 2975
box -3 -3 3 3
use M3_M2  M3_M2_8974
timestamp 1745462530
transform 1 0 2980 0 1 2975
box -3 -3 3 3
use M3_M2  M3_M2_8975
timestamp 1745462530
transform 1 0 4204 0 1 2465
box -3 -3 3 3
use M3_M2  M3_M2_8976
timestamp 1745462530
transform 1 0 3932 0 1 2465
box -3 -3 3 3
use M3_M2  M3_M2_8977
timestamp 1745462530
transform 1 0 3828 0 1 2485
box -3 -3 3 3
use M3_M2  M3_M2_8978
timestamp 1745462530
transform 1 0 3628 0 1 2485
box -3 -3 3 3
use M3_M2  M3_M2_8979
timestamp 1745462530
transform 1 0 3572 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_8980
timestamp 1745462530
transform 1 0 3572 0 1 2485
box -3 -3 3 3
use M3_M2  M3_M2_8981
timestamp 1745462530
transform 1 0 3500 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_8982
timestamp 1745462530
transform 1 0 3284 0 1 2495
box -3 -3 3 3
use M3_M2  M3_M2_8983
timestamp 1745462530
transform 1 0 3052 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_8984
timestamp 1745462530
transform 1 0 4236 0 1 2285
box -3 -3 3 3
use M3_M2  M3_M2_8985
timestamp 1745462530
transform 1 0 4196 0 1 2285
box -3 -3 3 3
use M3_M2  M3_M2_8986
timestamp 1745462530
transform 1 0 4156 0 1 2285
box -3 -3 3 3
use M3_M2  M3_M2_8987
timestamp 1745462530
transform 1 0 3948 0 1 2285
box -3 -3 3 3
use M3_M2  M3_M2_8988
timestamp 1745462530
transform 1 0 3892 0 1 2275
box -3 -3 3 3
use M3_M2  M3_M2_8989
timestamp 1745462530
transform 1 0 3636 0 1 2275
box -3 -3 3 3
use M3_M2  M3_M2_8990
timestamp 1745462530
transform 1 0 3388 0 1 2335
box -3 -3 3 3
use M3_M2  M3_M2_8991
timestamp 1745462530
transform 1 0 3388 0 1 2275
box -3 -3 3 3
use M3_M2  M3_M2_8992
timestamp 1745462530
transform 1 0 3260 0 1 2335
box -3 -3 3 3
use M3_M2  M3_M2_8993
timestamp 1745462530
transform 1 0 4116 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_8994
timestamp 1745462530
transform 1 0 4076 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_8995
timestamp 1745462530
transform 1 0 3860 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_8996
timestamp 1745462530
transform 1 0 3860 0 1 2885
box -3 -3 3 3
use M3_M2  M3_M2_8997
timestamp 1745462530
transform 1 0 3836 0 1 2885
box -3 -3 3 3
use M3_M2  M3_M2_8998
timestamp 1745462530
transform 1 0 3700 0 1 2885
box -3 -3 3 3
use M3_M2  M3_M2_8999
timestamp 1745462530
transform 1 0 3484 0 1 2885
box -3 -3 3 3
use M3_M2  M3_M2_9000
timestamp 1745462530
transform 1 0 3220 0 1 2935
box -3 -3 3 3
use M3_M2  M3_M2_9001
timestamp 1745462530
transform 1 0 3220 0 1 2885
box -3 -3 3 3
use M3_M2  M3_M2_9002
timestamp 1745462530
transform 1 0 3196 0 1 2935
box -3 -3 3 3
use M3_M2  M3_M2_9003
timestamp 1745462530
transform 1 0 3020 0 1 2645
box -3 -3 3 3
use M3_M2  M3_M2_9004
timestamp 1745462530
transform 1 0 2932 0 1 2415
box -3 -3 3 3
use M3_M2  M3_M2_9005
timestamp 1745462530
transform 1 0 2852 0 1 2645
box -3 -3 3 3
use M3_M2  M3_M2_9006
timestamp 1745462530
transform 1 0 2836 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_9007
timestamp 1745462530
transform 1 0 2804 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_9008
timestamp 1745462530
transform 1 0 2804 0 1 2405
box -3 -3 3 3
use M3_M2  M3_M2_9009
timestamp 1745462530
transform 1 0 2748 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_9010
timestamp 1745462530
transform 1 0 2828 0 1 2775
box -3 -3 3 3
use M3_M2  M3_M2_9011
timestamp 1745462530
transform 1 0 2788 0 1 2775
box -3 -3 3 3
use M3_M2  M3_M2_9012
timestamp 1745462530
transform 1 0 2764 0 1 2775
box -3 -3 3 3
use M3_M2  M3_M2_9013
timestamp 1745462530
transform 1 0 2676 0 1 2775
box -3 -3 3 3
use M3_M2  M3_M2_9014
timestamp 1745462530
transform 1 0 2604 0 1 2775
box -3 -3 3 3
use M3_M2  M3_M2_9015
timestamp 1745462530
transform 1 0 2484 0 1 2775
box -3 -3 3 3
use M3_M2  M3_M2_9016
timestamp 1745462530
transform 1 0 2484 0 1 2755
box -3 -3 3 3
use M3_M2  M3_M2_9017
timestamp 1745462530
transform 1 0 2420 0 1 2755
box -3 -3 3 3
use M3_M2  M3_M2_9018
timestamp 1745462530
transform 1 0 1764 0 1 1075
box -3 -3 3 3
use M3_M2  M3_M2_9019
timestamp 1745462530
transform 1 0 1628 0 1 1075
box -3 -3 3 3
use M3_M2  M3_M2_9020
timestamp 1745462530
transform 1 0 1788 0 1 2185
box -3 -3 3 3
use M3_M2  M3_M2_9021
timestamp 1745462530
transform 1 0 1764 0 1 2185
box -3 -3 3 3
use M3_M2  M3_M2_9022
timestamp 1745462530
transform 1 0 3788 0 1 2315
box -3 -3 3 3
use M3_M2  M3_M2_9023
timestamp 1745462530
transform 1 0 1796 0 1 2315
box -3 -3 3 3
use M3_M2  M3_M2_9024
timestamp 1745462530
transform 1 0 3900 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_9025
timestamp 1745462530
transform 1 0 3764 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_9026
timestamp 1745462530
transform 1 0 3868 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_9027
timestamp 1745462530
transform 1 0 3852 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_9028
timestamp 1745462530
transform 1 0 3772 0 1 2265
box -3 -3 3 3
use M3_M2  M3_M2_9029
timestamp 1745462530
transform 1 0 3740 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_9030
timestamp 1745462530
transform 1 0 3620 0 1 1855
box -3 -3 3 3
use M3_M2  M3_M2_9031
timestamp 1745462530
transform 1 0 3620 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_9032
timestamp 1745462530
transform 1 0 3532 0 1 1885
box -3 -3 3 3
use M3_M2  M3_M2_9033
timestamp 1745462530
transform 1 0 3532 0 1 1855
box -3 -3 3 3
use M3_M2  M3_M2_9034
timestamp 1745462530
transform 1 0 3508 0 1 2265
box -3 -3 3 3
use M3_M2  M3_M2_9035
timestamp 1745462530
transform 1 0 3508 0 1 2125
box -3 -3 3 3
use M3_M2  M3_M2_9036
timestamp 1745462530
transform 1 0 3500 0 1 1885
box -3 -3 3 3
use M3_M2  M3_M2_9037
timestamp 1745462530
transform 1 0 3476 0 1 2125
box -3 -3 3 3
use M3_M2  M3_M2_9038
timestamp 1745462530
transform 1 0 3716 0 1 1005
box -3 -3 3 3
use M3_M2  M3_M2_9039
timestamp 1745462530
transform 1 0 3004 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_9040
timestamp 1745462530
transform 1 0 3892 0 1 1005
box -3 -3 3 3
use M3_M2  M3_M2_9041
timestamp 1745462530
transform 1 0 3748 0 1 1005
box -3 -3 3 3
use M3_M2  M3_M2_9042
timestamp 1745462530
transform 1 0 3932 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_9043
timestamp 1745462530
transform 1 0 3868 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_9044
timestamp 1745462530
transform 1 0 3852 0 1 335
box -3 -3 3 3
use M3_M2  M3_M2_9045
timestamp 1745462530
transform 1 0 3772 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_9046
timestamp 1745462530
transform 1 0 3892 0 1 365
box -3 -3 3 3
use M3_M2  M3_M2_9047
timestamp 1745462530
transform 1 0 3788 0 1 365
box -3 -3 3 3
use M3_M2  M3_M2_9048
timestamp 1745462530
transform 1 0 3772 0 1 575
box -3 -3 3 3
use M3_M2  M3_M2_9049
timestamp 1745462530
transform 1 0 3692 0 1 575
box -3 -3 3 3
use M3_M2  M3_M2_9050
timestamp 1745462530
transform 1 0 3636 0 1 465
box -3 -3 3 3
use M3_M2  M3_M2_9051
timestamp 1745462530
transform 1 0 3564 0 1 575
box -3 -3 3 3
use M3_M2  M3_M2_9052
timestamp 1745462530
transform 1 0 3524 0 1 575
box -3 -3 3 3
use M3_M2  M3_M2_9053
timestamp 1745462530
transform 1 0 3524 0 1 465
box -3 -3 3 3
use M3_M2  M3_M2_9054
timestamp 1745462530
transform 1 0 3340 0 1 575
box -3 -3 3 3
use M3_M2  M3_M2_9055
timestamp 1745462530
transform 1 0 3964 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_9056
timestamp 1745462530
transform 1 0 3740 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_9057
timestamp 1745462530
transform 1 0 3700 0 1 455
box -3 -3 3 3
use M3_M2  M3_M2_9058
timestamp 1745462530
transform 1 0 3668 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_9059
timestamp 1745462530
transform 1 0 3668 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_9060
timestamp 1745462530
transform 1 0 3668 0 1 455
box -3 -3 3 3
use M3_M2  M3_M2_9061
timestamp 1745462530
transform 1 0 3596 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_9062
timestamp 1745462530
transform 1 0 3548 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_9063
timestamp 1745462530
transform 1 0 3396 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_9064
timestamp 1745462530
transform 1 0 3300 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_9065
timestamp 1745462530
transform 1 0 3772 0 1 365
box -3 -3 3 3
use M3_M2  M3_M2_9066
timestamp 1745462530
transform 1 0 3724 0 1 365
box -3 -3 3 3
use M3_M2  M3_M2_9067
timestamp 1745462530
transform 1 0 3580 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_9068
timestamp 1745462530
transform 1 0 3556 0 1 365
box -3 -3 3 3
use M3_M2  M3_M2_9069
timestamp 1745462530
transform 1 0 3436 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_9070
timestamp 1745462530
transform 1 0 3236 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_9071
timestamp 1745462530
transform 1 0 3852 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_9072
timestamp 1745462530
transform 1 0 3788 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_9073
timestamp 1745462530
transform 1 0 3636 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_9074
timestamp 1745462530
transform 1 0 3596 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_9075
timestamp 1745462530
transform 1 0 3596 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_9076
timestamp 1745462530
transform 1 0 3476 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_9077
timestamp 1745462530
transform 1 0 3300 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_9078
timestamp 1745462530
transform 1 0 3908 0 1 865
box -3 -3 3 3
use M3_M2  M3_M2_9079
timestamp 1745462530
transform 1 0 3860 0 1 865
box -3 -3 3 3
use M3_M2  M3_M2_9080
timestamp 1745462530
transform 1 0 3620 0 1 865
box -3 -3 3 3
use M3_M2  M3_M2_9081
timestamp 1745462530
transform 1 0 3484 0 1 1005
box -3 -3 3 3
use M3_M2  M3_M2_9082
timestamp 1745462530
transform 1 0 3484 0 1 865
box -3 -3 3 3
use M3_M2  M3_M2_9083
timestamp 1745462530
transform 1 0 3388 0 1 865
box -3 -3 3 3
use M3_M2  M3_M2_9084
timestamp 1745462530
transform 1 0 3388 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_9085
timestamp 1745462530
transform 1 0 3340 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_9086
timestamp 1745462530
transform 1 0 3244 0 1 1005
box -3 -3 3 3
use M3_M2  M3_M2_9087
timestamp 1745462530
transform 1 0 3940 0 1 845
box -3 -3 3 3
use M3_M2  M3_M2_9088
timestamp 1745462530
transform 1 0 3884 0 1 845
box -3 -3 3 3
use M3_M2  M3_M2_9089
timestamp 1745462530
transform 1 0 3652 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_9090
timestamp 1745462530
transform 1 0 3508 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_9091
timestamp 1745462530
transform 1 0 3508 0 1 845
box -3 -3 3 3
use M3_M2  M3_M2_9092
timestamp 1745462530
transform 1 0 3508 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_9093
timestamp 1745462530
transform 1 0 3380 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_9094
timestamp 1745462530
transform 1 0 3380 0 1 1085
box -3 -3 3 3
use M3_M2  M3_M2_9095
timestamp 1745462530
transform 1 0 3364 0 1 845
box -3 -3 3 3
use M3_M2  M3_M2_9096
timestamp 1745462530
transform 1 0 3236 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_9097
timestamp 1745462530
transform 1 0 3876 0 1 1075
box -3 -3 3 3
use M3_M2  M3_M2_9098
timestamp 1745462530
transform 1 0 3820 0 1 1075
box -3 -3 3 3
use M3_M2  M3_M2_9099
timestamp 1745462530
transform 1 0 3636 0 1 1075
box -3 -3 3 3
use M3_M2  M3_M2_9100
timestamp 1745462530
transform 1 0 3612 0 1 1075
box -3 -3 3 3
use M3_M2  M3_M2_9101
timestamp 1745462530
transform 1 0 3540 0 1 1075
box -3 -3 3 3
use M3_M2  M3_M2_9102
timestamp 1745462530
transform 1 0 3428 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_9103
timestamp 1745462530
transform 1 0 3428 0 1 1075
box -3 -3 3 3
use M3_M2  M3_M2_9104
timestamp 1745462530
transform 1 0 3308 0 1 1075
box -3 -3 3 3
use M3_M2  M3_M2_9105
timestamp 1745462530
transform 1 0 3268 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_9106
timestamp 1745462530
transform 1 0 3268 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_9107
timestamp 1745462530
transform 1 0 3196 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_9108
timestamp 1745462530
transform 1 0 3892 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_9109
timestamp 1745462530
transform 1 0 3852 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_9110
timestamp 1745462530
transform 1 0 3836 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_9111
timestamp 1745462530
transform 1 0 3692 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_9112
timestamp 1745462530
transform 1 0 3628 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_9113
timestamp 1745462530
transform 1 0 3572 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_9114
timestamp 1745462530
transform 1 0 3412 0 1 1335
box -3 -3 3 3
use M3_M2  M3_M2_9115
timestamp 1745462530
transform 1 0 3356 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_9116
timestamp 1745462530
transform 1 0 3332 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_9117
timestamp 1745462530
transform 1 0 3332 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_9118
timestamp 1745462530
transform 1 0 3212 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_9119
timestamp 1745462530
transform 1 0 2972 0 1 1005
box -3 -3 3 3
use M3_M2  M3_M2_9120
timestamp 1745462530
transform 1 0 2948 0 1 1005
box -3 -3 3 3
use M3_M2  M3_M2_9121
timestamp 1745462530
transform 1 0 3068 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_9122
timestamp 1745462530
transform 1 0 3044 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_9123
timestamp 1745462530
transform 1 0 3044 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_9124
timestamp 1745462530
transform 1 0 2988 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_9125
timestamp 1745462530
transform 1 0 2996 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_9126
timestamp 1745462530
transform 1 0 2964 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_9127
timestamp 1745462530
transform 1 0 2908 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_9128
timestamp 1745462530
transform 1 0 2812 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_9129
timestamp 1745462530
transform 1 0 2804 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_9130
timestamp 1745462530
transform 1 0 2684 0 1 495
box -3 -3 3 3
use M3_M2  M3_M2_9131
timestamp 1745462530
transform 1 0 2644 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_9132
timestamp 1745462530
transform 1 0 2572 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_9133
timestamp 1745462530
transform 1 0 2508 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_9134
timestamp 1745462530
transform 1 0 2508 0 1 495
box -3 -3 3 3
use M3_M2  M3_M2_9135
timestamp 1745462530
transform 1 0 2508 0 1 465
box -3 -3 3 3
use M3_M2  M3_M2_9136
timestamp 1745462530
transform 1 0 2452 0 1 495
box -3 -3 3 3
use M3_M2  M3_M2_9137
timestamp 1745462530
transform 1 0 2452 0 1 465
box -3 -3 3 3
use M3_M2  M3_M2_9138
timestamp 1745462530
transform 1 0 2372 0 1 495
box -3 -3 3 3
use M3_M2  M3_M2_9139
timestamp 1745462530
transform 1 0 2964 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_9140
timestamp 1745462530
transform 1 0 2860 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_9141
timestamp 1745462530
transform 1 0 2724 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_9142
timestamp 1745462530
transform 1 0 2604 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_9143
timestamp 1745462530
transform 1 0 2532 0 1 535
box -3 -3 3 3
use M3_M2  M3_M2_9144
timestamp 1745462530
transform 1 0 2484 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_9145
timestamp 1745462530
transform 1 0 2420 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_9146
timestamp 1745462530
transform 1 0 2908 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_9147
timestamp 1745462530
transform 1 0 2868 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_9148
timestamp 1745462530
transform 1 0 2836 0 1 675
box -3 -3 3 3
use M3_M2  M3_M2_9149
timestamp 1745462530
transform 1 0 2764 0 1 675
box -3 -3 3 3
use M3_M2  M3_M2_9150
timestamp 1745462530
transform 1 0 2644 0 1 675
box -3 -3 3 3
use M3_M2  M3_M2_9151
timestamp 1745462530
transform 1 0 2612 0 1 675
box -3 -3 3 3
use M3_M2  M3_M2_9152
timestamp 1745462530
transform 1 0 2460 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_9153
timestamp 1745462530
transform 1 0 2460 0 1 675
box -3 -3 3 3
use M3_M2  M3_M2_9154
timestamp 1745462530
transform 1 0 2316 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_9155
timestamp 1745462530
transform 1 0 2316 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_9156
timestamp 1745462530
transform 1 0 2252 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_9157
timestamp 1745462530
transform 1 0 2964 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_9158
timestamp 1745462530
transform 1 0 2908 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_9159
timestamp 1745462530
transform 1 0 2900 0 1 645
box -3 -3 3 3
use M3_M2  M3_M2_9160
timestamp 1745462530
transform 1 0 2796 0 1 645
box -3 -3 3 3
use M3_M2  M3_M2_9161
timestamp 1745462530
transform 1 0 2636 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_9162
timestamp 1745462530
transform 1 0 2604 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_9163
timestamp 1745462530
transform 1 0 2492 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_9164
timestamp 1745462530
transform 1 0 2348 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_9165
timestamp 1745462530
transform 1 0 2308 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_9166
timestamp 1745462530
transform 1 0 3036 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_9167
timestamp 1745462530
transform 1 0 2844 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_9168
timestamp 1745462530
transform 1 0 2828 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_9169
timestamp 1745462530
transform 1 0 2748 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_9170
timestamp 1745462530
transform 1 0 2748 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_9171
timestamp 1745462530
transform 1 0 2676 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_9172
timestamp 1745462530
transform 1 0 2636 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_9173
timestamp 1745462530
transform 1 0 2508 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_9174
timestamp 1745462530
transform 1 0 3100 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_9175
timestamp 1745462530
transform 1 0 3068 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_9176
timestamp 1745462530
transform 1 0 2980 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_9177
timestamp 1745462530
transform 1 0 2980 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_9178
timestamp 1745462530
transform 1 0 2852 0 1 1005
box -3 -3 3 3
use M3_M2  M3_M2_9179
timestamp 1745462530
transform 1 0 2852 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_9180
timestamp 1745462530
transform 1 0 2788 0 1 1005
box -3 -3 3 3
use M3_M2  M3_M2_9181
timestamp 1745462530
transform 1 0 2708 0 1 1005
box -3 -3 3 3
use M3_M2  M3_M2_9182
timestamp 1745462530
transform 1 0 2700 0 1 875
box -3 -3 3 3
use M3_M2  M3_M2_9183
timestamp 1745462530
transform 1 0 2652 0 1 875
box -3 -3 3 3
use M3_M2  M3_M2_9184
timestamp 1745462530
transform 1 0 2524 0 1 875
box -3 -3 3 3
use M3_M2  M3_M2_9185
timestamp 1745462530
transform 1 0 2964 0 1 1215
box -3 -3 3 3
use M3_M2  M3_M2_9186
timestamp 1745462530
transform 1 0 2916 0 1 1215
box -3 -3 3 3
use M3_M2  M3_M2_9187
timestamp 1745462530
transform 1 0 2756 0 1 1215
box -3 -3 3 3
use M3_M2  M3_M2_9188
timestamp 1745462530
transform 1 0 2724 0 1 1285
box -3 -3 3 3
use M3_M2  M3_M2_9189
timestamp 1745462530
transform 1 0 2532 0 1 1285
box -3 -3 3 3
use M3_M2  M3_M2_9190
timestamp 1745462530
transform 1 0 2508 0 1 1215
box -3 -3 3 3
use M3_M2  M3_M2_9191
timestamp 1745462530
transform 1 0 2436 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_9192
timestamp 1745462530
transform 1 0 3140 0 1 1065
box -3 -3 3 3
use M3_M2  M3_M2_9193
timestamp 1745462530
transform 1 0 3012 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_9194
timestamp 1745462530
transform 1 0 3012 0 1 1065
box -3 -3 3 3
use M3_M2  M3_M2_9195
timestamp 1745462530
transform 1 0 2948 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_9196
timestamp 1745462530
transform 1 0 2948 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_9197
timestamp 1745462530
transform 1 0 2820 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_9198
timestamp 1745462530
transform 1 0 2652 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_9199
timestamp 1745462530
transform 1 0 2524 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_9200
timestamp 1745462530
transform 1 0 2524 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_9201
timestamp 1745462530
transform 1 0 2492 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_9202
timestamp 1745462530
transform 1 0 4012 0 1 2675
box -3 -3 3 3
use M3_M2  M3_M2_9203
timestamp 1745462530
transform 1 0 3972 0 1 2675
box -3 -3 3 3
use M3_M2  M3_M2_9204
timestamp 1745462530
transform 1 0 4060 0 1 2705
box -3 -3 3 3
use M3_M2  M3_M2_9205
timestamp 1745462530
transform 1 0 3988 0 1 2705
box -3 -3 3 3
use M3_M2  M3_M2_9206
timestamp 1745462530
transform 1 0 4100 0 1 2685
box -3 -3 3 3
use M3_M2  M3_M2_9207
timestamp 1745462530
transform 1 0 4004 0 1 2685
box -3 -3 3 3
use M3_M2  M3_M2_9208
timestamp 1745462530
transform 1 0 4092 0 1 2605
box -3 -3 3 3
use M3_M2  M3_M2_9209
timestamp 1745462530
transform 1 0 4060 0 1 2605
box -3 -3 3 3
use M3_M2  M3_M2_9210
timestamp 1745462530
transform 1 0 3844 0 1 2605
box -3 -3 3 3
use M3_M2  M3_M2_9211
timestamp 1745462530
transform 1 0 3492 0 1 2605
box -3 -3 3 3
use M3_M2  M3_M2_9212
timestamp 1745462530
transform 1 0 3484 0 1 2545
box -3 -3 3 3
use M3_M2  M3_M2_9213
timestamp 1745462530
transform 1 0 3308 0 1 2535
box -3 -3 3 3
use M3_M2  M3_M2_9214
timestamp 1745462530
transform 1 0 3172 0 1 2565
box -3 -3 3 3
use M3_M2  M3_M2_9215
timestamp 1745462530
transform 1 0 3172 0 1 2545
box -3 -3 3 3
use M3_M2  M3_M2_9216
timestamp 1745462530
transform 1 0 3060 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_9217
timestamp 1745462530
transform 1 0 3060 0 1 2565
box -3 -3 3 3
use M3_M2  M3_M2_9218
timestamp 1745462530
transform 1 0 2980 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_9219
timestamp 1745462530
transform 1 0 2940 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_9220
timestamp 1745462530
transform 1 0 2940 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_9221
timestamp 1745462530
transform 1 0 2900 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_9222
timestamp 1745462530
transform 1 0 4172 0 1 2575
box -3 -3 3 3
use M3_M2  M3_M2_9223
timestamp 1745462530
transform 1 0 4108 0 1 2575
box -3 -3 3 3
use M3_M2  M3_M2_9224
timestamp 1745462530
transform 1 0 4148 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_9225
timestamp 1745462530
transform 1 0 4140 0 1 2415
box -3 -3 3 3
use M3_M2  M3_M2_9226
timestamp 1745462530
transform 1 0 4084 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_9227
timestamp 1745462530
transform 1 0 4084 0 1 2435
box -3 -3 3 3
use M3_M2  M3_M2_9228
timestamp 1745462530
transform 1 0 3868 0 1 2435
box -3 -3 3 3
use M3_M2  M3_M2_9229
timestamp 1745462530
transform 1 0 3804 0 1 2495
box -3 -3 3 3
use M3_M2  M3_M2_9230
timestamp 1745462530
transform 1 0 3804 0 1 2435
box -3 -3 3 3
use M3_M2  M3_M2_9231
timestamp 1745462530
transform 1 0 3524 0 1 2495
box -3 -3 3 3
use M3_M2  M3_M2_9232
timestamp 1745462530
transform 1 0 3356 0 1 2485
box -3 -3 3 3
use M3_M2  M3_M2_9233
timestamp 1745462530
transform 1 0 3188 0 1 2485
box -3 -3 3 3
use M3_M2  M3_M2_9234
timestamp 1745462530
transform 1 0 2604 0 1 2485
box -3 -3 3 3
use M3_M2  M3_M2_9235
timestamp 1745462530
transform 1 0 2604 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_9236
timestamp 1745462530
transform 1 0 2572 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_9237
timestamp 1745462530
transform 1 0 4188 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_9238
timestamp 1745462530
transform 1 0 4148 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_9239
timestamp 1745462530
transform 1 0 3916 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_9240
timestamp 1745462530
transform 1 0 3908 0 1 2405
box -3 -3 3 3
use M3_M2  M3_M2_9241
timestamp 1745462530
transform 1 0 3860 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_9242
timestamp 1745462530
transform 1 0 3548 0 1 2405
box -3 -3 3 3
use M3_M2  M3_M2_9243
timestamp 1745462530
transform 1 0 3396 0 1 2405
box -3 -3 3 3
use M3_M2  M3_M2_9244
timestamp 1745462530
transform 1 0 3220 0 1 2405
box -3 -3 3 3
use M3_M2  M3_M2_9245
timestamp 1745462530
transform 1 0 3220 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_9246
timestamp 1745462530
transform 1 0 2668 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_9247
timestamp 1745462530
transform 1 0 3988 0 1 2685
box -3 -3 3 3
use M3_M2  M3_M2_9248
timestamp 1745462530
transform 1 0 3900 0 1 2675
box -3 -3 3 3
use M3_M2  M3_M2_9249
timestamp 1745462530
transform 1 0 3724 0 1 2675
box -3 -3 3 3
use M3_M2  M3_M2_9250
timestamp 1745462530
transform 1 0 3556 0 1 2675
box -3 -3 3 3
use M3_M2  M3_M2_9251
timestamp 1745462530
transform 1 0 3412 0 1 2675
box -3 -3 3 3
use M3_M2  M3_M2_9252
timestamp 1745462530
transform 1 0 3412 0 1 2645
box -3 -3 3 3
use M3_M2  M3_M2_9253
timestamp 1745462530
transform 1 0 3100 0 1 2685
box -3 -3 3 3
use M3_M2  M3_M2_9254
timestamp 1745462530
transform 1 0 3100 0 1 2645
box -3 -3 3 3
use M3_M2  M3_M2_9255
timestamp 1745462530
transform 1 0 3068 0 1 2685
box -3 -3 3 3
use M3_M2  M3_M2_9256
timestamp 1745462530
transform 1 0 2708 0 1 2705
box -3 -3 3 3
use M3_M2  M3_M2_9257
timestamp 1745462530
transform 1 0 4004 0 1 2565
box -3 -3 3 3
use M3_M2  M3_M2_9258
timestamp 1745462530
transform 1 0 3940 0 1 2565
box -3 -3 3 3
use M3_M2  M3_M2_9259
timestamp 1745462530
transform 1 0 3764 0 1 2575
box -3 -3 3 3
use M3_M2  M3_M2_9260
timestamp 1745462530
transform 1 0 3612 0 1 2575
box -3 -3 3 3
use M3_M2  M3_M2_9261
timestamp 1745462530
transform 1 0 3404 0 1 2575
box -3 -3 3 3
use M3_M2  M3_M2_9262
timestamp 1745462530
transform 1 0 3396 0 1 2675
box -3 -3 3 3
use M3_M2  M3_M2_9263
timestamp 1745462530
transform 1 0 3108 0 1 2675
box -3 -3 3 3
use M3_M2  M3_M2_9264
timestamp 1745462530
transform 1 0 2764 0 1 2675
box -3 -3 3 3
use M3_M2  M3_M2_9265
timestamp 1745462530
transform 1 0 4036 0 1 2815
box -3 -3 3 3
use M3_M2  M3_M2_9266
timestamp 1745462530
transform 1 0 3780 0 1 2815
box -3 -3 3 3
use M3_M2  M3_M2_9267
timestamp 1745462530
transform 1 0 3532 0 1 2865
box -3 -3 3 3
use M3_M2  M3_M2_9268
timestamp 1745462530
transform 1 0 3532 0 1 2815
box -3 -3 3 3
use M3_M2  M3_M2_9269
timestamp 1745462530
transform 1 0 3300 0 1 2865
box -3 -3 3 3
use M3_M2  M3_M2_9270
timestamp 1745462530
transform 1 0 2988 0 1 2865
box -3 -3 3 3
use M3_M2  M3_M2_9271
timestamp 1745462530
transform 1 0 2956 0 1 2865
box -3 -3 3 3
use M3_M2  M3_M2_9272
timestamp 1745462530
transform 1 0 2644 0 1 2865
box -3 -3 3 3
use M3_M2  M3_M2_9273
timestamp 1745462530
transform 1 0 2644 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_9274
timestamp 1745462530
transform 1 0 2628 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_9275
timestamp 1745462530
transform 1 0 4052 0 1 2775
box -3 -3 3 3
use M3_M2  M3_M2_9276
timestamp 1745462530
transform 1 0 3812 0 1 2775
box -3 -3 3 3
use M3_M2  M3_M2_9277
timestamp 1745462530
transform 1 0 3572 0 1 2755
box -3 -3 3 3
use M3_M2  M3_M2_9278
timestamp 1745462530
transform 1 0 3340 0 1 2755
box -3 -3 3 3
use M3_M2  M3_M2_9279
timestamp 1745462530
transform 1 0 3020 0 1 2755
box -3 -3 3 3
use M3_M2  M3_M2_9280
timestamp 1745462530
transform 1 0 3004 0 1 2785
box -3 -3 3 3
use M3_M2  M3_M2_9281
timestamp 1745462530
transform 1 0 2708 0 1 2805
box -3 -3 3 3
use M3_M2  M3_M2_9282
timestamp 1745462530
transform 1 0 2708 0 1 2725
box -3 -3 3 3
use M3_M2  M3_M2_9283
timestamp 1745462530
transform 1 0 2676 0 1 2425
box -3 -3 3 3
use M3_M2  M3_M2_9284
timestamp 1745462530
transform 1 0 2612 0 1 2425
box -3 -3 3 3
use M3_M2  M3_M2_9285
timestamp 1745462530
transform 1 0 2596 0 1 2725
box -3 -3 3 3
use M3_M2  M3_M2_9286
timestamp 1745462530
transform 1 0 3868 0 1 2165
box -3 -3 3 3
use M3_M2  M3_M2_9287
timestamp 1745462530
transform 1 0 3820 0 1 2285
box -3 -3 3 3
use M3_M2  M3_M2_9288
timestamp 1745462530
transform 1 0 3820 0 1 2165
box -3 -3 3 3
use M3_M2  M3_M2_9289
timestamp 1745462530
transform 1 0 2988 0 1 2285
box -3 -3 3 3
use M3_M2  M3_M2_9290
timestamp 1745462530
transform 1 0 3924 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_9291
timestamp 1745462530
transform 1 0 3900 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_9292
timestamp 1745462530
transform 1 0 3964 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_9293
timestamp 1745462530
transform 1 0 3892 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_9294
timestamp 1745462530
transform 1 0 3844 0 1 1455
box -3 -3 3 3
use M3_M2  M3_M2_9295
timestamp 1745462530
transform 1 0 3732 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_9296
timestamp 1745462530
transform 1 0 3732 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_9297
timestamp 1745462530
transform 1 0 3676 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_9298
timestamp 1745462530
transform 1 0 3644 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_9299
timestamp 1745462530
transform 1 0 3588 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_9300
timestamp 1745462530
transform 1 0 3588 0 1 1455
box -3 -3 3 3
use M3_M2  M3_M2_9301
timestamp 1745462530
transform 1 0 3460 0 1 1455
box -3 -3 3 3
use M3_M2  M3_M2_9302
timestamp 1745462530
transform 1 0 3460 0 1 1435
box -3 -3 3 3
use M3_M2  M3_M2_9303
timestamp 1745462530
transform 1 0 3404 0 1 1435
box -3 -3 3 3
use M3_M2  M3_M2_9304
timestamp 1745462530
transform 1 0 3940 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_9305
timestamp 1745462530
transform 1 0 3924 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_9306
timestamp 1745462530
transform 1 0 3900 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_9307
timestamp 1745462530
transform 1 0 3828 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_9308
timestamp 1745462530
transform 1 0 3828 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_9309
timestamp 1745462530
transform 1 0 3772 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_9310
timestamp 1745462530
transform 1 0 3676 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_9311
timestamp 1745462530
transform 1 0 3668 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_9312
timestamp 1745462530
transform 1 0 3668 0 1 1465
box -3 -3 3 3
use M3_M2  M3_M2_9313
timestamp 1745462530
transform 1 0 3564 0 1 1465
box -3 -3 3 3
use M3_M2  M3_M2_9314
timestamp 1745462530
transform 1 0 3564 0 1 1375
box -3 -3 3 3
use M3_M2  M3_M2_9315
timestamp 1745462530
transform 1 0 3500 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_9316
timestamp 1745462530
transform 1 0 3492 0 1 1375
box -3 -3 3 3
use M3_M2  M3_M2_9317
timestamp 1745462530
transform 1 0 3340 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_9318
timestamp 1745462530
transform 1 0 3972 0 1 1885
box -3 -3 3 3
use M3_M2  M3_M2_9319
timestamp 1745462530
transform 1 0 3876 0 1 1885
box -3 -3 3 3
use M3_M2  M3_M2_9320
timestamp 1745462530
transform 1 0 3860 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_9321
timestamp 1745462530
transform 1 0 3748 0 1 1885
box -3 -3 3 3
use M3_M2  M3_M2_9322
timestamp 1745462530
transform 1 0 3748 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_9323
timestamp 1745462530
transform 1 0 3548 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_9324
timestamp 1745462530
transform 1 0 3516 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_9325
timestamp 1745462530
transform 1 0 3396 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_9326
timestamp 1745462530
transform 1 0 3364 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_9327
timestamp 1745462530
transform 1 0 3292 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_9328
timestamp 1745462530
transform 1 0 3932 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_9329
timestamp 1745462530
transform 1 0 3900 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_9330
timestamp 1745462530
transform 1 0 3788 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_9331
timestamp 1745462530
transform 1 0 3788 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_9332
timestamp 1745462530
transform 1 0 3780 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_9333
timestamp 1745462530
transform 1 0 3780 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_9334
timestamp 1745462530
transform 1 0 3780 0 1 1685
box -3 -3 3 3
use M3_M2  M3_M2_9335
timestamp 1745462530
transform 1 0 3772 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_9336
timestamp 1745462530
transform 1 0 3764 0 1 1685
box -3 -3 3 3
use M3_M2  M3_M2_9337
timestamp 1745462530
transform 1 0 3604 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_9338
timestamp 1745462530
transform 1 0 3572 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_9339
timestamp 1745462530
transform 1 0 3452 0 1 1375
box -3 -3 3 3
use M3_M2  M3_M2_9340
timestamp 1745462530
transform 1 0 3420 0 1 1375
box -3 -3 3 3
use M3_M2  M3_M2_9341
timestamp 1745462530
transform 1 0 3420 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_9342
timestamp 1745462530
transform 1 0 3268 0 1 1375
box -3 -3 3 3
use M3_M2  M3_M2_9343
timestamp 1745462530
transform 1 0 3820 0 1 1895
box -3 -3 3 3
use M3_M2  M3_M2_9344
timestamp 1745462530
transform 1 0 3804 0 1 2095
box -3 -3 3 3
use M3_M2  M3_M2_9345
timestamp 1745462530
transform 1 0 3748 0 1 2095
box -3 -3 3 3
use M3_M2  M3_M2_9346
timestamp 1745462530
transform 1 0 3748 0 1 1895
box -3 -3 3 3
use M3_M2  M3_M2_9347
timestamp 1745462530
transform 1 0 3548 0 1 2095
box -3 -3 3 3
use M3_M2  M3_M2_9348
timestamp 1745462530
transform 1 0 3444 0 1 2095
box -3 -3 3 3
use M3_M2  M3_M2_9349
timestamp 1745462530
transform 1 0 3316 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_9350
timestamp 1745462530
transform 1 0 3260 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_9351
timestamp 1745462530
transform 1 0 3204 0 1 2095
box -3 -3 3 3
use M3_M2  M3_M2_9352
timestamp 1745462530
transform 1 0 3172 0 1 2095
box -3 -3 3 3
use M3_M2  M3_M2_9353
timestamp 1745462530
transform 1 0 3844 0 1 2125
box -3 -3 3 3
use M3_M2  M3_M2_9354
timestamp 1745462530
transform 1 0 3812 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_9355
timestamp 1745462530
transform 1 0 3564 0 1 2125
box -3 -3 3 3
use M3_M2  M3_M2_9356
timestamp 1745462530
transform 1 0 3564 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_9357
timestamp 1745462530
transform 1 0 3460 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_9358
timestamp 1745462530
transform 1 0 3460 0 1 1935
box -3 -3 3 3
use M3_M2  M3_M2_9359
timestamp 1745462530
transform 1 0 3460 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_9360
timestamp 1745462530
transform 1 0 3460 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_9361
timestamp 1745462530
transform 1 0 3388 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_9362
timestamp 1745462530
transform 1 0 3252 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_9363
timestamp 1745462530
transform 1 0 3188 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_9364
timestamp 1745462530
transform 1 0 3060 0 1 2095
box -3 -3 3 3
use M3_M2  M3_M2_9365
timestamp 1745462530
transform 1 0 3020 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_9366
timestamp 1745462530
transform 1 0 3004 0 1 2455
box -3 -3 3 3
use M3_M2  M3_M2_9367
timestamp 1745462530
transform 1 0 3004 0 1 2385
box -3 -3 3 3
use M3_M2  M3_M2_9368
timestamp 1745462530
transform 1 0 3004 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_9369
timestamp 1745462530
transform 1 0 2948 0 1 2455
box -3 -3 3 3
use M3_M2  M3_M2_9370
timestamp 1745462530
transform 1 0 2948 0 1 2385
box -3 -3 3 3
use M3_M2  M3_M2_9371
timestamp 1745462530
transform 1 0 2948 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_9372
timestamp 1745462530
transform 1 0 2940 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_9373
timestamp 1745462530
transform 1 0 2876 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_9374
timestamp 1745462530
transform 1 0 1972 0 1 2285
box -3 -3 3 3
use M3_M2  M3_M2_9375
timestamp 1745462530
transform 1 0 1748 0 1 2285
box -3 -3 3 3
use M3_M2  M3_M2_9376
timestamp 1745462530
transform 1 0 1764 0 1 2215
box -3 -3 3 3
use M3_M2  M3_M2_9377
timestamp 1745462530
transform 1 0 684 0 1 2215
box -3 -3 3 3
use M3_M2  M3_M2_9378
timestamp 1745462530
transform 1 0 724 0 1 2085
box -3 -3 3 3
use M3_M2  M3_M2_9379
timestamp 1745462530
transform 1 0 684 0 1 2085
box -3 -3 3 3
use M3_M2  M3_M2_9380
timestamp 1745462530
transform 1 0 668 0 1 2235
box -3 -3 3 3
use M3_M2  M3_M2_9381
timestamp 1745462530
transform 1 0 620 0 1 2235
box -3 -3 3 3
use M3_M2  M3_M2_9382
timestamp 1745462530
transform 1 0 692 0 1 2465
box -3 -3 3 3
use M3_M2  M3_M2_9383
timestamp 1745462530
transform 1 0 652 0 1 2465
box -3 -3 3 3
use M3_M2  M3_M2_9384
timestamp 1745462530
transform 1 0 700 0 1 2405
box -3 -3 3 3
use M3_M2  M3_M2_9385
timestamp 1745462530
transform 1 0 668 0 1 2405
box -3 -3 3 3
use M3_M2  M3_M2_9386
timestamp 1745462530
transform 1 0 852 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_9387
timestamp 1745462530
transform 1 0 828 0 1 2445
box -3 -3 3 3
use M3_M2  M3_M2_9388
timestamp 1745462530
transform 1 0 724 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_9389
timestamp 1745462530
transform 1 0 724 0 1 2775
box -3 -3 3 3
use M3_M2  M3_M2_9390
timestamp 1745462530
transform 1 0 716 0 1 2445
box -3 -3 3 3
use M3_M2  M3_M2_9391
timestamp 1745462530
transform 1 0 692 0 1 2775
box -3 -3 3 3
use M3_M2  M3_M2_9392
timestamp 1745462530
transform 1 0 676 0 1 2435
box -3 -3 3 3
use M3_M2  M3_M2_9393
timestamp 1745462530
transform 1 0 452 0 1 2435
box -3 -3 3 3
use M3_M2  M3_M2_9394
timestamp 1745462530
transform 1 0 932 0 1 2725
box -3 -3 3 3
use M3_M2  M3_M2_9395
timestamp 1745462530
transform 1 0 908 0 1 2725
box -3 -3 3 3
use M3_M2  M3_M2_9396
timestamp 1745462530
transform 1 0 796 0 1 2725
box -3 -3 3 3
use M3_M2  M3_M2_9397
timestamp 1745462530
transform 1 0 788 0 1 2845
box -3 -3 3 3
use M3_M2  M3_M2_9398
timestamp 1745462530
transform 1 0 764 0 1 2845
box -3 -3 3 3
use M3_M2  M3_M2_9399
timestamp 1745462530
transform 1 0 756 0 1 2725
box -3 -3 3 3
use M3_M2  M3_M2_9400
timestamp 1745462530
transform 1 0 868 0 1 2465
box -3 -3 3 3
use M3_M2  M3_M2_9401
timestamp 1745462530
transform 1 0 804 0 1 2805
box -3 -3 3 3
use M3_M2  M3_M2_9402
timestamp 1745462530
transform 1 0 756 0 1 2805
box -3 -3 3 3
use M3_M2  M3_M2_9403
timestamp 1745462530
transform 1 0 676 0 1 2455
box -3 -3 3 3
use M3_M2  M3_M2_9404
timestamp 1745462530
transform 1 0 652 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_9405
timestamp 1745462530
transform 1 0 628 0 1 2665
box -3 -3 3 3
use M3_M2  M3_M2_9406
timestamp 1745462530
transform 1 0 516 0 1 2665
box -3 -3 3 3
use M3_M2  M3_M2_9407
timestamp 1745462530
transform 1 0 900 0 1 2565
box -3 -3 3 3
use M3_M2  M3_M2_9408
timestamp 1745462530
transform 1 0 868 0 1 2565
box -3 -3 3 3
use M3_M2  M3_M2_9409
timestamp 1745462530
transform 1 0 812 0 1 2765
box -3 -3 3 3
use M3_M2  M3_M2_9410
timestamp 1745462530
transform 1 0 716 0 1 2565
box -3 -3 3 3
use M3_M2  M3_M2_9411
timestamp 1745462530
transform 1 0 700 0 1 2765
box -3 -3 3 3
use M3_M2  M3_M2_9412
timestamp 1745462530
transform 1 0 692 0 1 2565
box -3 -3 3 3
use M3_M2  M3_M2_9413
timestamp 1745462530
transform 1 0 964 0 1 2245
box -3 -3 3 3
use M3_M2  M3_M2_9414
timestamp 1745462530
transform 1 0 788 0 1 2245
box -3 -3 3 3
use M3_M2  M3_M2_9415
timestamp 1745462530
transform 1 0 788 0 1 2165
box -3 -3 3 3
use M3_M2  M3_M2_9416
timestamp 1745462530
transform 1 0 692 0 1 2155
box -3 -3 3 3
use M3_M2  M3_M2_9417
timestamp 1745462530
transform 1 0 644 0 1 2155
box -3 -3 3 3
use M3_M2  M3_M2_9418
timestamp 1745462530
transform 1 0 588 0 1 2155
box -3 -3 3 3
use M3_M2  M3_M2_9419
timestamp 1745462530
transform 1 0 588 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_9420
timestamp 1745462530
transform 1 0 532 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_9421
timestamp 1745462530
transform 1 0 1012 0 1 2265
box -3 -3 3 3
use M3_M2  M3_M2_9422
timestamp 1745462530
transform 1 0 836 0 1 2265
box -3 -3 3 3
use M3_M2  M3_M2_9423
timestamp 1745462530
transform 1 0 836 0 1 2185
box -3 -3 3 3
use M3_M2  M3_M2_9424
timestamp 1745462530
transform 1 0 804 0 1 2185
box -3 -3 3 3
use M3_M2  M3_M2_9425
timestamp 1745462530
transform 1 0 804 0 1 2125
box -3 -3 3 3
use M3_M2  M3_M2_9426
timestamp 1745462530
transform 1 0 740 0 1 2185
box -3 -3 3 3
use M3_M2  M3_M2_9427
timestamp 1745462530
transform 1 0 660 0 1 2125
box -3 -3 3 3
use M3_M2  M3_M2_9428
timestamp 1745462530
transform 1 0 604 0 1 2125
box -3 -3 3 3
use M3_M2  M3_M2_9429
timestamp 1745462530
transform 1 0 940 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_9430
timestamp 1745462530
transform 1 0 908 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_9431
timestamp 1745462530
transform 1 0 804 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_9432
timestamp 1745462530
transform 1 0 788 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_9433
timestamp 1745462530
transform 1 0 740 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_9434
timestamp 1745462530
transform 1 0 684 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_9435
timestamp 1745462530
transform 1 0 652 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_9436
timestamp 1745462530
transform 1 0 1100 0 1 1975
box -3 -3 3 3
use M3_M2  M3_M2_9437
timestamp 1745462530
transform 1 0 932 0 1 1975
box -3 -3 3 3
use M3_M2  M3_M2_9438
timestamp 1745462530
transform 1 0 860 0 1 1975
box -3 -3 3 3
use M3_M2  M3_M2_9439
timestamp 1745462530
transform 1 0 796 0 1 1975
box -3 -3 3 3
use M3_M2  M3_M2_9440
timestamp 1745462530
transform 1 0 740 0 1 1975
box -3 -3 3 3
use M3_M2  M3_M2_9441
timestamp 1745462530
transform 1 0 668 0 1 1975
box -3 -3 3 3
use M3_M2  M3_M2_9442
timestamp 1745462530
transform 1 0 476 0 1 1975
box -3 -3 3 3
use M3_M2  M3_M2_9443
timestamp 1745462530
transform 1 0 1988 0 1 2415
box -3 -3 3 3
use M3_M2  M3_M2_9444
timestamp 1745462530
transform 1 0 1948 0 1 2415
box -3 -3 3 3
use M3_M2  M3_M2_9445
timestamp 1745462530
transform 1 0 2012 0 1 2355
box -3 -3 3 3
use M3_M2  M3_M2_9446
timestamp 1745462530
transform 1 0 1924 0 1 2355
box -3 -3 3 3
use M3_M2  M3_M2_9447
timestamp 1745462530
transform 1 0 1940 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_9448
timestamp 1745462530
transform 1 0 1724 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_9449
timestamp 1745462530
transform 1 0 1772 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_9450
timestamp 1745462530
transform 1 0 1708 0 1 2385
box -3 -3 3 3
use M3_M2  M3_M2_9451
timestamp 1745462530
transform 1 0 1708 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_9452
timestamp 1745462530
transform 1 0 1540 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_9453
timestamp 1745462530
transform 1 0 1324 0 1 2375
box -3 -3 3 3
use M3_M2  M3_M2_9454
timestamp 1745462530
transform 1 0 1180 0 1 2375
box -3 -3 3 3
use M3_M2  M3_M2_9455
timestamp 1745462530
transform 1 0 1124 0 1 2385
box -3 -3 3 3
use M3_M2  M3_M2_9456
timestamp 1745462530
transform 1 0 1036 0 1 2385
box -3 -3 3 3
use M3_M2  M3_M2_9457
timestamp 1745462530
transform 1 0 2076 0 1 2385
box -3 -3 3 3
use M3_M2  M3_M2_9458
timestamp 1745462530
transform 1 0 1812 0 1 2375
box -3 -3 3 3
use M3_M2  M3_M2_9459
timestamp 1745462530
transform 1 0 1748 0 1 2375
box -3 -3 3 3
use M3_M2  M3_M2_9460
timestamp 1745462530
transform 1 0 1732 0 1 2285
box -3 -3 3 3
use M3_M2  M3_M2_9461
timestamp 1745462530
transform 1 0 1596 0 1 2285
box -3 -3 3 3
use M3_M2  M3_M2_9462
timestamp 1745462530
transform 1 0 1420 0 1 2285
box -3 -3 3 3
use M3_M2  M3_M2_9463
timestamp 1745462530
transform 1 0 1388 0 1 2285
box -3 -3 3 3
use M3_M2  M3_M2_9464
timestamp 1745462530
transform 1 0 1236 0 1 2295
box -3 -3 3 3
use M3_M2  M3_M2_9465
timestamp 1745462530
transform 1 0 1156 0 1 2295
box -3 -3 3 3
use M3_M2  M3_M2_9466
timestamp 1745462530
transform 1 0 2108 0 1 2365
box -3 -3 3 3
use M3_M2  M3_M2_9467
timestamp 1745462530
transform 1 0 1980 0 1 2365
box -3 -3 3 3
use M3_M2  M3_M2_9468
timestamp 1745462530
transform 1 0 1844 0 1 2365
box -3 -3 3 3
use M3_M2  M3_M2_9469
timestamp 1745462530
transform 1 0 1652 0 1 2375
box -3 -3 3 3
use M3_M2  M3_M2_9470
timestamp 1745462530
transform 1 0 1652 0 1 2315
box -3 -3 3 3
use M3_M2  M3_M2_9471
timestamp 1745462530
transform 1 0 1500 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_9472
timestamp 1745462530
transform 1 0 1500 0 1 2315
box -3 -3 3 3
use M3_M2  M3_M2_9473
timestamp 1745462530
transform 1 0 1444 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_9474
timestamp 1745462530
transform 1 0 1420 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_9475
timestamp 1745462530
transform 1 0 1412 0 1 2445
box -3 -3 3 3
use M3_M2  M3_M2_9476
timestamp 1745462530
transform 1 0 1380 0 1 2445
box -3 -3 3 3
use M3_M2  M3_M2_9477
timestamp 1745462530
transform 1 0 1212 0 1 2445
box -3 -3 3 3
use M3_M2  M3_M2_9478
timestamp 1745462530
transform 1 0 2124 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_9479
timestamp 1745462530
transform 1 0 2028 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_9480
timestamp 1745462530
transform 1 0 1924 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_9481
timestamp 1745462530
transform 1 0 1860 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_9482
timestamp 1745462530
transform 1 0 1860 0 1 2265
box -3 -3 3 3
use M3_M2  M3_M2_9483
timestamp 1745462530
transform 1 0 1692 0 1 2265
box -3 -3 3 3
use M3_M2  M3_M2_9484
timestamp 1745462530
transform 1 0 1484 0 1 2265
box -3 -3 3 3
use M3_M2  M3_M2_9485
timestamp 1745462530
transform 1 0 1476 0 1 2245
box -3 -3 3 3
use M3_M2  M3_M2_9486
timestamp 1745462530
transform 1 0 1388 0 1 2245
box -3 -3 3 3
use M3_M2  M3_M2_9487
timestamp 1745462530
transform 1 0 1308 0 1 2245
box -3 -3 3 3
use M3_M2  M3_M2_9488
timestamp 1745462530
transform 1 0 2396 0 1 2875
box -3 -3 3 3
use M3_M2  M3_M2_9489
timestamp 1745462530
transform 1 0 2220 0 1 2875
box -3 -3 3 3
use M3_M2  M3_M2_9490
timestamp 1745462530
transform 1 0 1980 0 1 2875
box -3 -3 3 3
use M3_M2  M3_M2_9491
timestamp 1745462530
transform 1 0 1908 0 1 2875
box -3 -3 3 3
use M3_M2  M3_M2_9492
timestamp 1745462530
transform 1 0 1652 0 1 2875
box -3 -3 3 3
use M3_M2  M3_M2_9493
timestamp 1745462530
transform 1 0 1500 0 1 2885
box -3 -3 3 3
use M3_M2  M3_M2_9494
timestamp 1745462530
transform 1 0 1444 0 1 2885
box -3 -3 3 3
use M3_M2  M3_M2_9495
timestamp 1745462530
transform 1 0 2068 0 1 2755
box -3 -3 3 3
use M3_M2  M3_M2_9496
timestamp 1745462530
transform 1 0 2012 0 1 2755
box -3 -3 3 3
use M3_M2  M3_M2_9497
timestamp 1745462530
transform 1 0 2004 0 1 2915
box -3 -3 3 3
use M3_M2  M3_M2_9498
timestamp 1745462530
transform 1 0 1948 0 1 2915
box -3 -3 3 3
use M3_M2  M3_M2_9499
timestamp 1745462530
transform 1 0 1692 0 1 2915
box -3 -3 3 3
use M3_M2  M3_M2_9500
timestamp 1745462530
transform 1 0 1516 0 1 2915
box -3 -3 3 3
use M3_M2  M3_M2_9501
timestamp 1745462530
transform 1 0 1460 0 1 2915
box -3 -3 3 3
use M3_M2  M3_M2_9502
timestamp 1745462530
transform 1 0 2140 0 1 2455
box -3 -3 3 3
use M3_M2  M3_M2_9503
timestamp 1745462530
transform 1 0 1972 0 1 2445
box -3 -3 3 3
use M3_M2  M3_M2_9504
timestamp 1745462530
transform 1 0 1972 0 1 2375
box -3 -3 3 3
use M3_M2  M3_M2_9505
timestamp 1745462530
transform 1 0 1924 0 1 2375
box -3 -3 3 3
use M3_M2  M3_M2_9506
timestamp 1745462530
transform 1 0 1628 0 1 2445
box -3 -3 3 3
use M3_M2  M3_M2_9507
timestamp 1745462530
transform 1 0 1628 0 1 2375
box -3 -3 3 3
use M3_M2  M3_M2_9508
timestamp 1745462530
transform 1 0 1516 0 1 2365
box -3 -3 3 3
use M3_M2  M3_M2_9509
timestamp 1745462530
transform 1 0 1508 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_9510
timestamp 1745462530
transform 1 0 1412 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_9511
timestamp 1745462530
transform 1 0 1404 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_9512
timestamp 1745462530
transform 1 0 1332 0 1 2405
box -3 -3 3 3
use M3_M2  M3_M2_9513
timestamp 1745462530
transform 1 0 1316 0 1 2405
box -3 -3 3 3
use M3_M2  M3_M2_9514
timestamp 1745462530
transform 1 0 1308 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_9515
timestamp 1745462530
transform 1 0 1196 0 1 2405
box -3 -3 3 3
use M3_M2  M3_M2_9516
timestamp 1745462530
transform 1 0 2156 0 1 2405
box -3 -3 3 3
use M3_M2  M3_M2_9517
timestamp 1745462530
transform 1 0 1980 0 1 2405
box -3 -3 3 3
use M3_M2  M3_M2_9518
timestamp 1745462530
transform 1 0 1916 0 1 2405
box -3 -3 3 3
use M3_M2  M3_M2_9519
timestamp 1745462530
transform 1 0 1748 0 1 2475
box -3 -3 3 3
use M3_M2  M3_M2_9520
timestamp 1745462530
transform 1 0 1748 0 1 2405
box -3 -3 3 3
use M3_M2  M3_M2_9521
timestamp 1745462530
transform 1 0 1684 0 1 2475
box -3 -3 3 3
use M3_M2  M3_M2_9522
timestamp 1745462530
transform 1 0 1572 0 1 2475
box -3 -3 3 3
use M3_M2  M3_M2_9523
timestamp 1745462530
transform 1 0 1452 0 1 2475
box -3 -3 3 3
use M3_M2  M3_M2_9524
timestamp 1745462530
transform 1 0 1372 0 1 2475
box -3 -3 3 3
use M3_M2  M3_M2_9525
timestamp 1745462530
transform 1 0 1204 0 1 2475
box -3 -3 3 3
use M3_M2  M3_M2_9526
timestamp 1745462530
transform 1 0 1620 0 1 1045
box -3 -3 3 3
use M3_M2  M3_M2_9527
timestamp 1745462530
transform 1 0 708 0 1 1045
box -3 -3 3 3
use M3_M2  M3_M2_9528
timestamp 1745462530
transform 1 0 1676 0 1 1035
box -3 -3 3 3
use M3_M2  M3_M2_9529
timestamp 1745462530
transform 1 0 1636 0 1 1035
box -3 -3 3 3
use M3_M2  M3_M2_9530
timestamp 1745462530
transform 1 0 1644 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_9531
timestamp 1745462530
transform 1 0 1620 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_9532
timestamp 1745462530
transform 1 0 1980 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_9533
timestamp 1745462530
transform 1 0 1924 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_9534
timestamp 1745462530
transform 1 0 1788 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_9535
timestamp 1745462530
transform 1 0 1668 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_9536
timestamp 1745462530
transform 1 0 1500 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_9537
timestamp 1745462530
transform 1 0 1420 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_9538
timestamp 1745462530
transform 1 0 1308 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_9539
timestamp 1745462530
transform 1 0 1308 0 1 575
box -3 -3 3 3
use M3_M2  M3_M2_9540
timestamp 1745462530
transform 1 0 1244 0 1 575
box -3 -3 3 3
use M3_M2  M3_M2_9541
timestamp 1745462530
transform 1 0 1972 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_9542
timestamp 1745462530
transform 1 0 1884 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_9543
timestamp 1745462530
transform 1 0 1828 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_9544
timestamp 1745462530
transform 1 0 1716 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_9545
timestamp 1745462530
transform 1 0 1580 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_9546
timestamp 1745462530
transform 1 0 1580 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_9547
timestamp 1745462530
transform 1 0 1452 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_9548
timestamp 1745462530
transform 1 0 1348 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_9549
timestamp 1745462530
transform 1 0 1348 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_9550
timestamp 1745462530
transform 1 0 1300 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_9551
timestamp 1745462530
transform 1 0 1900 0 1 495
box -3 -3 3 3
use M3_M2  M3_M2_9552
timestamp 1745462530
transform 1 0 1836 0 1 495
box -3 -3 3 3
use M3_M2  M3_M2_9553
timestamp 1745462530
transform 1 0 1588 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_9554
timestamp 1745462530
transform 1 0 1348 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_9555
timestamp 1745462530
transform 1 0 1268 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_9556
timestamp 1745462530
transform 1 0 1164 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_9557
timestamp 1745462530
transform 1 0 1164 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_9558
timestamp 1745462530
transform 1 0 1092 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_9559
timestamp 1745462530
transform 1 0 1956 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_9560
timestamp 1745462530
transform 1 0 1900 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_9561
timestamp 1745462530
transform 1 0 1636 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_9562
timestamp 1745462530
transform 1 0 1636 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_9563
timestamp 1745462530
transform 1 0 1564 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_9564
timestamp 1745462530
transform 1 0 1380 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_9565
timestamp 1745462530
transform 1 0 1196 0 1 575
box -3 -3 3 3
use M3_M2  M3_M2_9566
timestamp 1745462530
transform 1 0 1196 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_9567
timestamp 1745462530
transform 1 0 1132 0 1 575
box -3 -3 3 3
use M3_M2  M3_M2_9568
timestamp 1745462530
transform 1 0 1956 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_9569
timestamp 1745462530
transform 1 0 1900 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_9570
timestamp 1745462530
transform 1 0 1636 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_9571
timestamp 1745462530
transform 1 0 1628 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_9572
timestamp 1745462530
transform 1 0 1476 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_9573
timestamp 1745462530
transform 1 0 1460 0 1 1065
box -3 -3 3 3
use M3_M2  M3_M2_9574
timestamp 1745462530
transform 1 0 1460 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_9575
timestamp 1745462530
transform 1 0 1228 0 1 1065
box -3 -3 3 3
use M3_M2  M3_M2_9576
timestamp 1745462530
transform 1 0 1972 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_9577
timestamp 1745462530
transform 1 0 1916 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_9578
timestamp 1745462530
transform 1 0 1916 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_9579
timestamp 1745462530
transform 1 0 1676 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_9580
timestamp 1745462530
transform 1 0 1492 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_9581
timestamp 1745462530
transform 1 0 1380 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_9582
timestamp 1745462530
transform 1 0 1244 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_9583
timestamp 1745462530
transform 1 0 2068 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_9584
timestamp 1745462530
transform 1 0 1900 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_9585
timestamp 1745462530
transform 1 0 1876 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_9586
timestamp 1745462530
transform 1 0 1644 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_9587
timestamp 1745462530
transform 1 0 1508 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_9588
timestamp 1745462530
transform 1 0 1452 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_9589
timestamp 1745462530
transform 1 0 1260 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_9590
timestamp 1745462530
transform 1 0 2292 0 1 1265
box -3 -3 3 3
use M3_M2  M3_M2_9591
timestamp 1745462530
transform 1 0 2124 0 1 1265
box -3 -3 3 3
use M3_M2  M3_M2_9592
timestamp 1745462530
transform 1 0 2124 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_9593
timestamp 1745462530
transform 1 0 2084 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_9594
timestamp 1745462530
transform 1 0 1916 0 1 1265
box -3 -3 3 3
use M3_M2  M3_M2_9595
timestamp 1745462530
transform 1 0 1668 0 1 1265
box -3 -3 3 3
use M3_M2  M3_M2_9596
timestamp 1745462530
transform 1 0 1532 0 1 1265
box -3 -3 3 3
use M3_M2  M3_M2_9597
timestamp 1745462530
transform 1 0 1532 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_9598
timestamp 1745462530
transform 1 0 1508 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_9599
timestamp 1745462530
transform 1 0 1324 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_9600
timestamp 1745462530
transform 1 0 700 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_9601
timestamp 1745462530
transform 1 0 428 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_9602
timestamp 1745462530
transform 1 0 412 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_9603
timestamp 1745462530
transform 1 0 340 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_9604
timestamp 1745462530
transform 1 0 484 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_9605
timestamp 1745462530
transform 1 0 468 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_9606
timestamp 1745462530
transform 1 0 836 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_9607
timestamp 1745462530
transform 1 0 508 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_9608
timestamp 1745462530
transform 1 0 452 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_9609
timestamp 1745462530
transform 1 0 356 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_9610
timestamp 1745462530
transform 1 0 308 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_9611
timestamp 1745462530
transform 1 0 916 0 1 655
box -3 -3 3 3
use M3_M2  M3_M2_9612
timestamp 1745462530
transform 1 0 540 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_9613
timestamp 1745462530
transform 1 0 540 0 1 575
box -3 -3 3 3
use M3_M2  M3_M2_9614
timestamp 1745462530
transform 1 0 500 0 1 575
box -3 -3 3 3
use M3_M2  M3_M2_9615
timestamp 1745462530
transform 1 0 412 0 1 575
box -3 -3 3 3
use M3_M2  M3_M2_9616
timestamp 1745462530
transform 1 0 388 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_9617
timestamp 1745462530
transform 1 0 348 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_9618
timestamp 1745462530
transform 1 0 836 0 1 775
box -3 -3 3 3
use M3_M2  M3_M2_9619
timestamp 1745462530
transform 1 0 468 0 1 775
box -3 -3 3 3
use M3_M2  M3_M2_9620
timestamp 1745462530
transform 1 0 404 0 1 775
box -3 -3 3 3
use M3_M2  M3_M2_9621
timestamp 1745462530
transform 1 0 308 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_9622
timestamp 1745462530
transform 1 0 300 0 1 775
box -3 -3 3 3
use M3_M2  M3_M2_9623
timestamp 1745462530
transform 1 0 276 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_9624
timestamp 1745462530
transform 1 0 900 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_9625
timestamp 1745462530
transform 1 0 516 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_9626
timestamp 1745462530
transform 1 0 516 0 1 815
box -3 -3 3 3
use M3_M2  M3_M2_9627
timestamp 1745462530
transform 1 0 436 0 1 815
box -3 -3 3 3
use M3_M2  M3_M2_9628
timestamp 1745462530
transform 1 0 428 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_9629
timestamp 1745462530
transform 1 0 364 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_9630
timestamp 1745462530
transform 1 0 356 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_9631
timestamp 1745462530
transform 1 0 348 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_9632
timestamp 1745462530
transform 1 0 340 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_9633
timestamp 1745462530
transform 1 0 324 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_9634
timestamp 1745462530
transform 1 0 972 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_9635
timestamp 1745462530
transform 1 0 916 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_9636
timestamp 1745462530
transform 1 0 892 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_9637
timestamp 1745462530
transform 1 0 892 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_9638
timestamp 1745462530
transform 1 0 868 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_9639
timestamp 1745462530
transform 1 0 860 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_9640
timestamp 1745462530
transform 1 0 764 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_9641
timestamp 1745462530
transform 1 0 1020 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_9642
timestamp 1745462530
transform 1 0 964 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_9643
timestamp 1745462530
transform 1 0 956 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_9644
timestamp 1745462530
transform 1 0 940 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_9645
timestamp 1745462530
transform 1 0 916 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_9646
timestamp 1745462530
transform 1 0 908 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_9647
timestamp 1745462530
transform 1 0 804 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_9648
timestamp 1745462530
transform 1 0 764 0 1 725
box -3 -3 3 3
use M3_M2  M3_M2_9649
timestamp 1745462530
transform 1 0 716 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_9650
timestamp 1745462530
transform 1 0 700 0 1 725
box -3 -3 3 3
use M3_M2  M3_M2_9651
timestamp 1745462530
transform 1 0 1124 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_9652
timestamp 1745462530
transform 1 0 1100 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_9653
timestamp 1745462530
transform 1 0 1100 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_9654
timestamp 1745462530
transform 1 0 1036 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_9655
timestamp 1745462530
transform 1 0 988 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_9656
timestamp 1745462530
transform 1 0 804 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_9657
timestamp 1745462530
transform 1 0 804 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_9658
timestamp 1745462530
transform 1 0 748 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_9659
timestamp 1745462530
transform 1 0 676 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_9660
timestamp 1745462530
transform 1 0 676 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_9661
timestamp 1745462530
transform 1 0 628 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_9662
timestamp 1745462530
transform 1 0 1164 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_9663
timestamp 1745462530
transform 1 0 1084 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_9664
timestamp 1745462530
transform 1 0 1028 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_9665
timestamp 1745462530
transform 1 0 964 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_9666
timestamp 1745462530
transform 1 0 964 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_9667
timestamp 1745462530
transform 1 0 836 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_9668
timestamp 1745462530
transform 1 0 764 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_9669
timestamp 1745462530
transform 1 0 700 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_9670
timestamp 1745462530
transform 1 0 700 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_9671
timestamp 1745462530
transform 1 0 668 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_9672
timestamp 1745462530
transform 1 0 2564 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_9673
timestamp 1745462530
transform 1 0 1660 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_9674
timestamp 1745462530
transform 1 0 1652 0 1 1655
box -3 -3 3 3
use M3_M2  M3_M2_9675
timestamp 1745462530
transform 1 0 1620 0 1 1655
box -3 -3 3 3
use M3_M2  M3_M2_9676
timestamp 1745462530
transform 1 0 1492 0 1 1835
box -3 -3 3 3
use M3_M2  M3_M2_9677
timestamp 1745462530
transform 1 0 1412 0 1 1835
box -3 -3 3 3
use M3_M2  M3_M2_9678
timestamp 1745462530
transform 1 0 3044 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_9679
timestamp 1745462530
transform 1 0 1484 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_9680
timestamp 1745462530
transform 1 0 3156 0 1 1055
box -3 -3 3 3
use M3_M2  M3_M2_9681
timestamp 1745462530
transform 1 0 3020 0 1 1055
box -3 -3 3 3
use M3_M2  M3_M2_9682
timestamp 1745462530
transform 1 0 3140 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_9683
timestamp 1745462530
transform 1 0 3028 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_9684
timestamp 1745462530
transform 1 0 3308 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_9685
timestamp 1745462530
transform 1 0 3164 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_9686
timestamp 1745462530
transform 1 0 3332 0 1 865
box -3 -3 3 3
use M3_M2  M3_M2_9687
timestamp 1745462530
transform 1 0 3268 0 1 865
box -3 -3 3 3
use M3_M2  M3_M2_9688
timestamp 1745462530
transform 1 0 3324 0 1 845
box -3 -3 3 3
use M3_M2  M3_M2_9689
timestamp 1745462530
transform 1 0 3276 0 1 845
box -3 -3 3 3
use M3_M2  M3_M2_9690
timestamp 1745462530
transform 1 0 3332 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_9691
timestamp 1745462530
transform 1 0 3292 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_9692
timestamp 1745462530
transform 1 0 3060 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_9693
timestamp 1745462530
transform 1 0 3012 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_9694
timestamp 1745462530
transform 1 0 2996 0 1 675
box -3 -3 3 3
use M3_M2  M3_M2_9695
timestamp 1745462530
transform 1 0 2852 0 1 675
box -3 -3 3 3
use M3_M2  M3_M2_9696
timestamp 1745462530
transform 1 0 3108 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_9697
timestamp 1745462530
transform 1 0 3044 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_9698
timestamp 1745462530
transform 1 0 3156 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_9699
timestamp 1745462530
transform 1 0 3084 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_9700
timestamp 1745462530
transform 1 0 3124 0 1 2775
box -3 -3 3 3
use M3_M2  M3_M2_9701
timestamp 1745462530
transform 1 0 3020 0 1 2785
box -3 -3 3 3
use M3_M2  M3_M2_9702
timestamp 1745462530
transform 1 0 3068 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_9703
timestamp 1745462530
transform 1 0 2932 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_9704
timestamp 1745462530
transform 1 0 3204 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_9705
timestamp 1745462530
transform 1 0 3092 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_9706
timestamp 1745462530
transform 1 0 3356 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_9707
timestamp 1745462530
transform 1 0 3092 0 1 1695
box -3 -3 3 3
use M3_M2  M3_M2_9708
timestamp 1745462530
transform 1 0 3420 0 1 1455
box -3 -3 3 3
use M3_M2  M3_M2_9709
timestamp 1745462530
transform 1 0 3372 0 1 1455
box -3 -3 3 3
use M3_M2  M3_M2_9710
timestamp 1745462530
transform 1 0 3484 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_9711
timestamp 1745462530
transform 1 0 3388 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_9712
timestamp 1745462530
transform 1 0 1452 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_9713
timestamp 1745462530
transform 1 0 1420 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_9714
timestamp 1745462530
transform 1 0 1436 0 1 2085
box -3 -3 3 3
use M3_M2  M3_M2_9715
timestamp 1745462530
transform 1 0 772 0 1 2085
box -3 -3 3 3
use M3_M2  M3_M2_9716
timestamp 1745462530
transform 1 0 796 0 1 2095
box -3 -3 3 3
use M3_M2  M3_M2_9717
timestamp 1745462530
transform 1 0 724 0 1 2095
box -3 -3 3 3
use M3_M2  M3_M2_9718
timestamp 1745462530
transform 1 0 740 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_9719
timestamp 1745462530
transform 1 0 652 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_9720
timestamp 1745462530
transform 1 0 748 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_9721
timestamp 1745462530
transform 1 0 708 0 1 2745
box -3 -3 3 3
use M3_M2  M3_M2_9722
timestamp 1745462530
transform 1 0 684 0 1 2745
box -3 -3 3 3
use M3_M2  M3_M2_9723
timestamp 1745462530
transform 1 0 676 0 1 2775
box -3 -3 3 3
use M3_M2  M3_M2_9724
timestamp 1745462530
transform 1 0 540 0 1 2775
box -3 -3 3 3
use M3_M2  M3_M2_9725
timestamp 1745462530
transform 1 0 540 0 1 2705
box -3 -3 3 3
use M3_M2  M3_M2_9726
timestamp 1745462530
transform 1 0 516 0 1 2705
box -3 -3 3 3
use M3_M2  M3_M2_9727
timestamp 1745462530
transform 1 0 516 0 1 2675
box -3 -3 3 3
use M3_M2  M3_M2_9728
timestamp 1745462530
transform 1 0 492 0 1 2535
box -3 -3 3 3
use M3_M2  M3_M2_9729
timestamp 1745462530
transform 1 0 492 0 1 2175
box -3 -3 3 3
use M3_M2  M3_M2_9730
timestamp 1745462530
transform 1 0 484 0 1 2675
box -3 -3 3 3
use M3_M2  M3_M2_9731
timestamp 1745462530
transform 1 0 468 0 1 2535
box -3 -3 3 3
use M3_M2  M3_M2_9732
timestamp 1745462530
transform 1 0 1388 0 1 2405
box -3 -3 3 3
use M3_M2  M3_M2_9733
timestamp 1745462530
transform 1 0 1364 0 1 2405
box -3 -3 3 3
use M3_M2  M3_M2_9734
timestamp 1745462530
transform 1 0 1436 0 1 2805
box -3 -3 3 3
use M3_M2  M3_M2_9735
timestamp 1745462530
transform 1 0 1420 0 1 2805
box -3 -3 3 3
use M3_M2  M3_M2_9736
timestamp 1745462530
transform 1 0 1420 0 1 2385
box -3 -3 3 3
use M3_M2  M3_M2_9737
timestamp 1745462530
transform 1 0 1316 0 1 2385
box -3 -3 3 3
use M3_M2  M3_M2_9738
timestamp 1745462530
transform 1 0 1324 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_9739
timestamp 1745462530
transform 1 0 1204 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_9740
timestamp 1745462530
transform 1 0 1524 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_9741
timestamp 1745462530
transform 1 0 1500 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_9742
timestamp 1745462530
transform 1 0 1500 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_9743
timestamp 1745462530
transform 1 0 708 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_9744
timestamp 1745462530
transform 1 0 1460 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_9745
timestamp 1745462530
transform 1 0 1364 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_9746
timestamp 1745462530
transform 1 0 1492 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_9747
timestamp 1745462530
transform 1 0 1436 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_9748
timestamp 1745462530
transform 1 0 668 0 1 815
box -3 -3 3 3
use M3_M2  M3_M2_9749
timestamp 1745462530
transform 1 0 556 0 1 815
box -3 -3 3 3
use M3_M2  M3_M2_9750
timestamp 1745462530
transform 1 0 516 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_9751
timestamp 1745462530
transform 1 0 500 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_9752
timestamp 1745462530
transform 1 0 540 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_9753
timestamp 1745462530
transform 1 0 388 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_9754
timestamp 1745462530
transform 1 0 2164 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_9755
timestamp 1745462530
transform 1 0 1772 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_9756
timestamp 1745462530
transform 1 0 1644 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_9757
timestamp 1745462530
transform 1 0 1684 0 1 1655
box -3 -3 3 3
use M3_M2  M3_M2_9758
timestamp 1745462530
transform 1 0 1596 0 1 1975
box -3 -3 3 3
use M3_M2  M3_M2_9759
timestamp 1745462530
transform 1 0 1596 0 1 1665
box -3 -3 3 3
use M3_M2  M3_M2_9760
timestamp 1745462530
transform 1 0 1580 0 1 1975
box -3 -3 3 3
use M3_M2  M3_M2_9761
timestamp 1745462530
transform 1 0 3076 0 1 1495
box -3 -3 3 3
use M3_M2  M3_M2_9762
timestamp 1745462530
transform 1 0 1772 0 1 1525
box -3 -3 3 3
use M3_M2  M3_M2_9763
timestamp 1745462530
transform 1 0 1772 0 1 1495
box -3 -3 3 3
use M3_M2  M3_M2_9764
timestamp 1745462530
transform 1 0 1732 0 1 1525
box -3 -3 3 3
use M3_M2  M3_M2_9765
timestamp 1745462530
transform 1 0 3452 0 1 1615
box -3 -3 3 3
use M3_M2  M3_M2_9766
timestamp 1745462530
transform 1 0 3060 0 1 1615
box -3 -3 3 3
use M3_M2  M3_M2_9767
timestamp 1745462530
transform 1 0 3188 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_9768
timestamp 1745462530
transform 1 0 3148 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_9769
timestamp 1745462530
transform 1 0 3132 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_9770
timestamp 1745462530
transform 1 0 3076 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_9771
timestamp 1745462530
transform 1 0 3148 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_9772
timestamp 1745462530
transform 1 0 2436 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_9773
timestamp 1745462530
transform 1 0 3876 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_9774
timestamp 1745462530
transform 1 0 3188 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_9775
timestamp 1745462530
transform 1 0 3924 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_9776
timestamp 1745462530
transform 1 0 3876 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_9777
timestamp 1745462530
transform 1 0 2444 0 1 1215
box -3 -3 3 3
use M3_M2  M3_M2_9778
timestamp 1745462530
transform 1 0 2404 0 1 1215
box -3 -3 3 3
use M3_M2  M3_M2_9779
timestamp 1745462530
transform 1 0 2484 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_9780
timestamp 1745462530
transform 1 0 2428 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_9781
timestamp 1745462530
transform 1 0 2420 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_9782
timestamp 1745462530
transform 1 0 2268 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_9783
timestamp 1745462530
transform 1 0 2452 0 1 605
box -3 -3 3 3
use M3_M2  M3_M2_9784
timestamp 1745462530
transform 1 0 2404 0 1 605
box -3 -3 3 3
use M3_M2  M3_M2_9785
timestamp 1745462530
transform 1 0 4444 0 1 2615
box -3 -3 3 3
use M3_M2  M3_M2_9786
timestamp 1745462530
transform 1 0 4444 0 1 1875
box -3 -3 3 3
use M3_M2  M3_M2_9787
timestamp 1745462530
transform 1 0 4060 0 1 2615
box -3 -3 3 3
use M3_M2  M3_M2_9788
timestamp 1745462530
transform 1 0 3476 0 1 1875
box -3 -3 3 3
use M3_M2  M3_M2_9789
timestamp 1745462530
transform 1 0 4156 0 1 2525
box -3 -3 3 3
use M3_M2  M3_M2_9790
timestamp 1745462530
transform 1 0 4084 0 1 2525
box -3 -3 3 3
use M3_M2  M3_M2_9791
timestamp 1745462530
transform 1 0 3380 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_9792
timestamp 1745462530
transform 1 0 2868 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_9793
timestamp 1745462530
transform 1 0 3420 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_9794
timestamp 1745462530
transform 1 0 3356 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_9795
timestamp 1745462530
transform 1 0 3516 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_9796
timestamp 1745462530
transform 1 0 3428 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_9797
timestamp 1745462530
transform 1 0 3588 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_9798
timestamp 1745462530
transform 1 0 3548 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_9799
timestamp 1745462530
transform 1 0 3636 0 1 1485
box -3 -3 3 3
use M3_M2  M3_M2_9800
timestamp 1745462530
transform 1 0 3620 0 1 1485
box -3 -3 3 3
use M3_M2  M3_M2_9801
timestamp 1745462530
transform 1 0 1628 0 1 2185
box -3 -3 3 3
use M3_M2  M3_M2_9802
timestamp 1745462530
transform 1 0 1580 0 1 2185
box -3 -3 3 3
use M3_M2  M3_M2_9803
timestamp 1745462530
transform 1 0 1580 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_9804
timestamp 1745462530
transform 1 0 740 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_9805
timestamp 1745462530
transform 1 0 676 0 1 2055
box -3 -3 3 3
use M3_M2  M3_M2_9806
timestamp 1745462530
transform 1 0 652 0 1 2055
box -3 -3 3 3
use M3_M2  M3_M2_9807
timestamp 1745462530
transform 1 0 692 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_9808
timestamp 1745462530
transform 1 0 596 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_9809
timestamp 1745462530
transform 1 0 700 0 1 2235
box -3 -3 3 3
use M3_M2  M3_M2_9810
timestamp 1745462530
transform 1 0 684 0 1 2235
box -3 -3 3 3
use M3_M2  M3_M2_9811
timestamp 1745462530
transform 1 0 732 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_9812
timestamp 1745462530
transform 1 0 700 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_9813
timestamp 1745462530
transform 1 0 1668 0 1 2405
box -3 -3 3 3
use M3_M2  M3_M2_9814
timestamp 1745462530
transform 1 0 1596 0 1 2405
box -3 -3 3 3
use M3_M2  M3_M2_9815
timestamp 1745462530
transform 1 0 1668 0 1 2885
box -3 -3 3 3
use M3_M2  M3_M2_9816
timestamp 1745462530
transform 1 0 1644 0 1 2885
box -3 -3 3 3
use M3_M2  M3_M2_9817
timestamp 1745462530
transform 1 0 1668 0 1 2365
box -3 -3 3 3
use M3_M2  M3_M2_9818
timestamp 1745462530
transform 1 0 1612 0 1 2365
box -3 -3 3 3
use M3_M2  M3_M2_9819
timestamp 1745462530
transform 1 0 1628 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_9820
timestamp 1745462530
transform 1 0 1572 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_9821
timestamp 1745462530
transform 1 0 1708 0 1 875
box -3 -3 3 3
use M3_M2  M3_M2_9822
timestamp 1745462530
transform 1 0 772 0 1 875
box -3 -3 3 3
use M3_M2  M3_M2_9823
timestamp 1745462530
transform 1 0 1876 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_9824
timestamp 1745462530
transform 1 0 1732 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_9825
timestamp 1745462530
transform 1 0 1900 0 1 1215
box -3 -3 3 3
use M3_M2  M3_M2_9826
timestamp 1745462530
transform 1 0 1804 0 1 1215
box -3 -3 3 3
use M3_M2  M3_M2_9827
timestamp 1745462530
transform 1 0 1908 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_9828
timestamp 1745462530
transform 1 0 1852 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_9829
timestamp 1745462530
transform 1 0 1876 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_9830
timestamp 1745462530
transform 1 0 1836 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_9831
timestamp 1745462530
transform 1 0 716 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_9832
timestamp 1745462530
transform 1 0 492 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_9833
timestamp 1745462530
transform 1 0 476 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_9834
timestamp 1745462530
transform 1 0 372 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_9835
timestamp 1745462530
transform 1 0 2140 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_9836
timestamp 1745462530
transform 1 0 1844 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_9837
timestamp 1745462530
transform 1 0 1908 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_9838
timestamp 1745462530
transform 1 0 1900 0 1 1275
box -3 -3 3 3
use M3_M2  M3_M2_9839
timestamp 1745462530
transform 1 0 1868 0 1 1275
box -3 -3 3 3
use M3_M2  M3_M2_9840
timestamp 1745462530
transform 1 0 1868 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_9841
timestamp 1745462530
transform 1 0 3588 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_9842
timestamp 1745462530
transform 1 0 3372 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_9843
timestamp 1745462530
transform 1 0 3340 0 1 1525
box -3 -3 3 3
use M3_M2  M3_M2_9844
timestamp 1745462530
transform 1 0 1876 0 1 1525
box -3 -3 3 3
use M3_M2  M3_M2_9845
timestamp 1745462530
transform 1 0 3748 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_9846
timestamp 1745462530
transform 1 0 3556 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_9847
timestamp 1745462530
transform 1 0 3548 0 1 775
box -3 -3 3 3
use M3_M2  M3_M2_9848
timestamp 1745462530
transform 1 0 2580 0 1 775
box -3 -3 3 3
use M3_M2  M3_M2_9849
timestamp 1745462530
transform 1 0 3772 0 1 815
box -3 -3 3 3
use M3_M2  M3_M2_9850
timestamp 1745462530
transform 1 0 3572 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_9851
timestamp 1745462530
transform 1 0 3748 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_9852
timestamp 1745462530
transform 1 0 3684 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_9853
timestamp 1745462530
transform 1 0 3876 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_9854
timestamp 1745462530
transform 1 0 3740 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_9855
timestamp 1745462530
transform 1 0 3764 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_9856
timestamp 1745462530
transform 1 0 3668 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_9857
timestamp 1745462530
transform 1 0 3660 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_9858
timestamp 1745462530
transform 1 0 3620 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_9859
timestamp 1745462530
transform 1 0 3724 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_9860
timestamp 1745462530
transform 1 0 3708 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_9861
timestamp 1745462530
transform 1 0 2540 0 1 845
box -3 -3 3 3
use M3_M2  M3_M2_9862
timestamp 1745462530
transform 1 0 2516 0 1 845
box -3 -3 3 3
use M3_M2  M3_M2_9863
timestamp 1745462530
transform 1 0 2556 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_9864
timestamp 1745462530
transform 1 0 2484 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_9865
timestamp 1745462530
transform 1 0 2588 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_9866
timestamp 1745462530
transform 1 0 2540 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_9867
timestamp 1745462530
transform 1 0 3812 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_9868
timestamp 1745462530
transform 1 0 3788 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_9869
timestamp 1745462530
transform 1 0 3796 0 1 2625
box -3 -3 3 3
use M3_M2  M3_M2_9870
timestamp 1745462530
transform 1 0 3748 0 1 2625
box -3 -3 3 3
use M3_M2  M3_M2_9871
timestamp 1745462530
transform 1 0 3844 0 1 2615
box -3 -3 3 3
use M3_M2  M3_M2_9872
timestamp 1745462530
transform 1 0 3804 0 1 2615
box -3 -3 3 3
use M3_M2  M3_M2_9873
timestamp 1745462530
transform 1 0 3924 0 1 2575
box -3 -3 3 3
use M3_M2  M3_M2_9874
timestamp 1745462530
transform 1 0 3852 0 1 2575
box -3 -3 3 3
use M3_M2  M3_M2_9875
timestamp 1745462530
transform 1 0 3732 0 1 1685
box -3 -3 3 3
use M3_M2  M3_M2_9876
timestamp 1745462530
transform 1 0 2996 0 1 1685
box -3 -3 3 3
use M3_M2  M3_M2_9877
timestamp 1745462530
transform 1 0 3804 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_9878
timestamp 1745462530
transform 1 0 3748 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_9879
timestamp 1745462530
transform 1 0 3812 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_9880
timestamp 1745462530
transform 1 0 3772 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_9881
timestamp 1745462530
transform 1 0 3892 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_9882
timestamp 1745462530
transform 1 0 3820 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_9883
timestamp 1745462530
transform 1 0 1940 0 1 2185
box -3 -3 3 3
use M3_M2  M3_M2_9884
timestamp 1745462530
transform 1 0 1908 0 1 2375
box -3 -3 3 3
use M3_M2  M3_M2_9885
timestamp 1745462530
transform 1 0 1884 0 1 2375
box -3 -3 3 3
use M3_M2  M3_M2_9886
timestamp 1745462530
transform 1 0 1868 0 1 2185
box -3 -3 3 3
use M3_M2  M3_M2_9887
timestamp 1745462530
transform 1 0 1884 0 1 2095
box -3 -3 3 3
use M3_M2  M3_M2_9888
timestamp 1745462530
transform 1 0 860 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_9889
timestamp 1745462530
transform 1 0 852 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_9890
timestamp 1745462530
transform 1 0 836 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_9891
timestamp 1745462530
transform 1 0 844 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_9892
timestamp 1745462530
transform 1 0 796 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_9893
timestamp 1745462530
transform 1 0 820 0 1 2835
box -3 -3 3 3
use M3_M2  M3_M2_9894
timestamp 1745462530
transform 1 0 796 0 1 2835
box -3 -3 3 3
use M3_M2  M3_M2_9895
timestamp 1745462530
transform 1 0 1908 0 1 2415
box -3 -3 3 3
use M3_M2  M3_M2_9896
timestamp 1745462530
transform 1 0 1852 0 1 2415
box -3 -3 3 3
use M3_M2  M3_M2_9897
timestamp 1745462530
transform 1 0 1932 0 1 2835
box -3 -3 3 3
use M3_M2  M3_M2_9898
timestamp 1745462530
transform 1 0 1860 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_9899
timestamp 1745462530
transform 1 0 1796 0 1 2835
box -3 -3 3 3
use M3_M2  M3_M2_9900
timestamp 1745462530
transform 1 0 1796 0 1 2535
box -3 -3 3 3
use M3_M2  M3_M2_9901
timestamp 1745462530
transform 1 0 1876 0 1 2355
box -3 -3 3 3
use M3_M2  M3_M2_9902
timestamp 1745462530
transform 1 0 1828 0 1 2355
box -3 -3 3 3
use M3_M2  M3_M2_9903
timestamp 1745462530
transform 1 0 1844 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_9904
timestamp 1745462530
transform 1 0 1788 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_9905
timestamp 1745462530
transform 1 0 1916 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_9906
timestamp 1745462530
transform 1 0 908 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_9907
timestamp 1745462530
transform 1 0 2028 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_9908
timestamp 1745462530
transform 1 0 1940 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_9909
timestamp 1745462530
transform 1 0 2076 0 1 1015
box -3 -3 3 3
use M3_M2  M3_M2_9910
timestamp 1745462530
transform 1 0 1996 0 1 1015
box -3 -3 3 3
use M3_M2  M3_M2_9911
timestamp 1745462530
transform 1 0 2020 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_9912
timestamp 1745462530
transform 1 0 1940 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_9913
timestamp 1745462530
transform 1 0 2060 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_9914
timestamp 1745462530
transform 1 0 1956 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_9915
timestamp 1745462530
transform 1 0 932 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_9916
timestamp 1745462530
transform 1 0 860 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_9917
timestamp 1745462530
transform 1 0 836 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_9918
timestamp 1745462530
transform 1 0 396 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_9919
timestamp 1745462530
transform 1 0 340 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_9920
timestamp 1745462530
transform 1 0 324 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_9921
timestamp 1745462530
transform 1 0 372 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_9922
timestamp 1745462530
transform 1 0 324 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_9923
timestamp 1745462530
transform 1 0 2364 0 1 1975
box -3 -3 3 3
use M3_M2  M3_M2_9924
timestamp 1745462530
transform 1 0 2332 0 1 1975
box -3 -3 3 3
use M3_M2  M3_M2_9925
timestamp 1745462530
transform 1 0 2332 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_9926
timestamp 1745462530
transform 1 0 1244 0 1 2155
box -3 -3 3 3
use M3_M2  M3_M2_9927
timestamp 1745462530
transform 1 0 1244 0 1 2055
box -3 -3 3 3
use M3_M2  M3_M2_9928
timestamp 1745462530
transform 1 0 1220 0 1 2055
box -3 -3 3 3
use M3_M2  M3_M2_9929
timestamp 1745462530
transform 1 0 1212 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_9930
timestamp 1745462530
transform 1 0 1148 0 1 2155
box -3 -3 3 3
use M3_M2  M3_M2_9931
timestamp 1745462530
transform 1 0 1228 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_9932
timestamp 1745462530
transform 1 0 1164 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_9933
timestamp 1745462530
transform 1 0 1164 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_9934
timestamp 1745462530
transform 1 0 1132 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_9935
timestamp 1745462530
transform 1 0 1124 0 1 2165
box -3 -3 3 3
use M3_M2  M3_M2_9936
timestamp 1745462530
transform 1 0 1108 0 1 2165
box -3 -3 3 3
use M3_M2  M3_M2_9937
timestamp 1745462530
transform 1 0 3252 0 1 2155
box -3 -3 3 3
use M3_M2  M3_M2_9938
timestamp 1745462530
transform 1 0 1284 0 1 2245
box -3 -3 3 3
use M3_M2  M3_M2_9939
timestamp 1745462530
transform 1 0 1284 0 1 2155
box -3 -3 3 3
use M3_M2  M3_M2_9940
timestamp 1745462530
transform 1 0 1108 0 1 2245
box -3 -3 3 3
use M3_M2  M3_M2_9941
timestamp 1745462530
transform 1 0 3260 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_9942
timestamp 1745462530
transform 1 0 3204 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_9943
timestamp 1745462530
transform 1 0 3260 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_9944
timestamp 1745462530
transform 1 0 3260 0 1 1855
box -3 -3 3 3
use M3_M2  M3_M2_9945
timestamp 1745462530
transform 1 0 3244 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_9946
timestamp 1745462530
transform 1 0 3220 0 1 1855
box -3 -3 3 3
use M3_M2  M3_M2_9947
timestamp 1745462530
transform 1 0 3220 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_9948
timestamp 1745462530
transform 1 0 3212 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_9949
timestamp 1745462530
transform 1 0 3244 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_9950
timestamp 1745462530
transform 1 0 2620 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_9951
timestamp 1745462530
transform 1 0 3460 0 1 815
box -3 -3 3 3
use M3_M2  M3_M2_9952
timestamp 1745462530
transform 1 0 3276 0 1 815
box -3 -3 3 3
use M3_M2  M3_M2_9953
timestamp 1745462530
transform 1 0 3548 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_9954
timestamp 1745462530
transform 1 0 3420 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_9955
timestamp 1745462530
transform 1 0 3500 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_9956
timestamp 1745462530
transform 1 0 3444 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_9957
timestamp 1745462530
transform 1 0 3572 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_9958
timestamp 1745462530
transform 1 0 3508 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_9959
timestamp 1745462530
transform 1 0 2660 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_9960
timestamp 1745462530
transform 1 0 2652 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_9961
timestamp 1745462530
transform 1 0 2588 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_9962
timestamp 1745462530
transform 1 0 2516 0 1 1205
box -3 -3 3 3
use M3_M2  M3_M2_9963
timestamp 1745462530
transform 1 0 2636 0 1 845
box -3 -3 3 3
use M3_M2  M3_M2_9964
timestamp 1745462530
transform 1 0 2588 0 1 845
box -3 -3 3 3
use M3_M2  M3_M2_9965
timestamp 1745462530
transform 1 0 2604 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_9966
timestamp 1745462530
transform 1 0 2524 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_9967
timestamp 1745462530
transform 1 0 2524 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_9968
timestamp 1745462530
transform 1 0 2500 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_9969
timestamp 1745462530
transform 1 0 2452 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_9970
timestamp 1745462530
transform 1 0 2332 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_9971
timestamp 1745462530
transform 1 0 3324 0 1 2065
box -3 -3 3 3
use M3_M2  M3_M2_9972
timestamp 1745462530
transform 1 0 3228 0 1 2065
box -3 -3 3 3
use M3_M2  M3_M2_9973
timestamp 1745462530
transform 1 0 3364 0 1 2625
box -3 -3 3 3
use M3_M2  M3_M2_9974
timestamp 1745462530
transform 1 0 3324 0 1 2625
box -3 -3 3 3
use M3_M2  M3_M2_9975
timestamp 1745462530
transform 1 0 3380 0 1 2725
box -3 -3 3 3
use M3_M2  M3_M2_9976
timestamp 1745462530
transform 1 0 3340 0 1 2725
box -3 -3 3 3
use M3_M2  M3_M2_9977
timestamp 1745462530
transform 1 0 3356 0 1 2695
box -3 -3 3 3
use M3_M2  M3_M2_9978
timestamp 1745462530
transform 1 0 3340 0 1 2695
box -3 -3 3 3
use M3_M2  M3_M2_9979
timestamp 1745462530
transform 1 0 3292 0 1 2085
box -3 -3 3 3
use M3_M2  M3_M2_9980
timestamp 1745462530
transform 1 0 2948 0 1 2085
box -3 -3 3 3
use M3_M2  M3_M2_9981
timestamp 1745462530
transform 1 0 3452 0 1 2085
box -3 -3 3 3
use M3_M2  M3_M2_9982
timestamp 1745462530
transform 1 0 3308 0 1 2085
box -3 -3 3 3
use M3_M2  M3_M2_9983
timestamp 1745462530
transform 1 0 3476 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_9984
timestamp 1745462530
transform 1 0 3316 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_9985
timestamp 1745462530
transform 1 0 3532 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_9986
timestamp 1745462530
transform 1 0 3468 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_9987
timestamp 1745462530
transform 1 0 3660 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_9988
timestamp 1745462530
transform 1 0 3484 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_9989
timestamp 1745462530
transform 1 0 1092 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_9990
timestamp 1745462530
transform 1 0 908 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_9991
timestamp 1745462530
transform 1 0 948 0 1 2165
box -3 -3 3 3
use M3_M2  M3_M2_9992
timestamp 1745462530
transform 1 0 948 0 1 2065
box -3 -3 3 3
use M3_M2  M3_M2_9993
timestamp 1745462530
transform 1 0 924 0 1 2065
box -3 -3 3 3
use M3_M2  M3_M2_9994
timestamp 1745462530
transform 1 0 860 0 1 2165
box -3 -3 3 3
use M3_M2  M3_M2_9995
timestamp 1745462530
transform 1 0 852 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_9996
timestamp 1745462530
transform 1 0 828 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_9997
timestamp 1745462530
transform 1 0 892 0 1 2575
box -3 -3 3 3
use M3_M2  M3_M2_9998
timestamp 1745462530
transform 1 0 860 0 1 2575
box -3 -3 3 3
use M3_M2  M3_M2_9999
timestamp 1745462530
transform 1 0 1196 0 1 2445
box -3 -3 3 3
use M3_M2  M3_M2_10000
timestamp 1745462530
transform 1 0 1092 0 1 2445
box -3 -3 3 3
use M3_M2  M3_M2_10001
timestamp 1745462530
transform 1 0 1452 0 1 2865
box -3 -3 3 3
use M3_M2  M3_M2_10002
timestamp 1745462530
transform 1 0 1116 0 1 2865
box -3 -3 3 3
use M3_M2  M3_M2_10003
timestamp 1745462530
transform 1 0 1244 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_10004
timestamp 1745462530
transform 1 0 1140 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_10005
timestamp 1745462530
transform 1 0 1156 0 1 2385
box -3 -3 3 3
use M3_M2  M3_M2_10006
timestamp 1745462530
transform 1 0 1140 0 1 2385
box -3 -3 3 3
use M3_M2  M3_M2_10007
timestamp 1745462530
transform 1 0 1172 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_10008
timestamp 1745462530
transform 1 0 852 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_10009
timestamp 1745462530
transform 1 0 1252 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_10010
timestamp 1745462530
transform 1 0 1212 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_10011
timestamp 1745462530
transform 1 0 1324 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_10012
timestamp 1745462530
transform 1 0 1244 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_10013
timestamp 1745462530
transform 1 0 996 0 1 1065
box -3 -3 3 3
use M3_M2  M3_M2_10014
timestamp 1745462530
transform 1 0 820 0 1 1065
box -3 -3 3 3
use M3_M2  M3_M2_10015
timestamp 1745462530
transform 1 0 900 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_10016
timestamp 1745462530
transform 1 0 820 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_10017
timestamp 1745462530
transform 1 0 804 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_10018
timestamp 1745462530
transform 1 0 348 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_10019
timestamp 1745462530
transform 1 0 2196 0 1 2005
box -3 -3 3 3
use M3_M2  M3_M2_10020
timestamp 1745462530
transform 1 0 1508 0 1 2005
box -3 -3 3 3
use M3_M2  M3_M2_10021
timestamp 1745462530
transform 1 0 1476 0 1 2005
box -3 -3 3 3
use M3_M2  M3_M2_10022
timestamp 1745462530
transform 1 0 1484 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_10023
timestamp 1745462530
transform 1 0 1132 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_10024
timestamp 1745462530
transform 1 0 3140 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_10025
timestamp 1745462530
transform 1 0 1596 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_10026
timestamp 1745462530
transform 1 0 1596 0 1 2085
box -3 -3 3 3
use M3_M2  M3_M2_10027
timestamp 1745462530
transform 1 0 1508 0 1 2085
box -3 -3 3 3
use M3_M2  M3_M2_10028
timestamp 1745462530
transform 1 0 3476 0 1 2235
box -3 -3 3 3
use M3_M2  M3_M2_10029
timestamp 1745462530
transform 1 0 3116 0 1 2235
box -3 -3 3 3
use M3_M2  M3_M2_10030
timestamp 1745462530
transform 1 0 3196 0 1 1875
box -3 -3 3 3
use M3_M2  M3_M2_10031
timestamp 1745462530
transform 1 0 3124 0 1 1875
box -3 -3 3 3
use M3_M2  M3_M2_10032
timestamp 1745462530
transform 1 0 3196 0 1 885
box -3 -3 3 3
use M3_M2  M3_M2_10033
timestamp 1745462530
transform 1 0 2884 0 1 885
box -3 -3 3 3
use M3_M2  M3_M2_10034
timestamp 1745462530
transform 1 0 3604 0 1 885
box -3 -3 3 3
use M3_M2  M3_M2_10035
timestamp 1745462530
transform 1 0 3244 0 1 885
box -3 -3 3 3
use M3_M2  M3_M2_10036
timestamp 1745462530
transform 1 0 3644 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_10037
timestamp 1745462530
transform 1 0 3588 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_10038
timestamp 1745462530
transform 1 0 3612 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_10039
timestamp 1745462530
transform 1 0 3580 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_10040
timestamp 1745462530
transform 1 0 3268 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_10041
timestamp 1745462530
transform 1 0 3236 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_10042
timestamp 1745462530
transform 1 0 3236 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_10043
timestamp 1745462530
transform 1 0 3196 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_10044
timestamp 1745462530
transform 1 0 3188 0 1 1375
box -3 -3 3 3
use M3_M2  M3_M2_10045
timestamp 1745462530
transform 1 0 2756 0 1 1865
box -3 -3 3 3
use M3_M2  M3_M2_10046
timestamp 1745462530
transform 1 0 2748 0 1 1375
box -3 -3 3 3
use M3_M2  M3_M2_10047
timestamp 1745462530
transform 1 0 2676 0 1 1375
box -3 -3 3 3
use M3_M2  M3_M2_10048
timestamp 1745462530
transform 1 0 2372 0 1 2055
box -3 -3 3 3
use M3_M2  M3_M2_10049
timestamp 1745462530
transform 1 0 2372 0 1 1865
box -3 -3 3 3
use M3_M2  M3_M2_10050
timestamp 1745462530
transform 1 0 2260 0 1 2055
box -3 -3 3 3
use M3_M2  M3_M2_10051
timestamp 1745462530
transform 1 0 3228 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_10052
timestamp 1745462530
transform 1 0 3188 0 1 1855
box -3 -3 3 3
use M3_M2  M3_M2_10053
timestamp 1745462530
transform 1 0 2732 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_10054
timestamp 1745462530
transform 1 0 2316 0 1 1975
box -3 -3 3 3
use M3_M2  M3_M2_10055
timestamp 1745462530
transform 1 0 2300 0 1 2215
box -3 -3 3 3
use M3_M2  M3_M2_10056
timestamp 1745462530
transform 1 0 2212 0 1 2215
box -3 -3 3 3
use M3_M2  M3_M2_10057
timestamp 1745462530
transform 1 0 2172 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_10058
timestamp 1745462530
transform 1 0 2172 0 1 1855
box -3 -3 3 3
use M3_M2  M3_M2_10059
timestamp 1745462530
transform 1 0 2172 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_10060
timestamp 1745462530
transform 1 0 1404 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_10061
timestamp 1745462530
transform 1 0 1404 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_10062
timestamp 1745462530
transform 1 0 1052 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_10063
timestamp 1745462530
transform 1 0 1044 0 1 1135
box -3 -3 3 3
use M3_M2  M3_M2_10064
timestamp 1745462530
transform 1 0 1004 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_10065
timestamp 1745462530
transform 1 0 988 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_10066
timestamp 1745462530
transform 1 0 988 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_10067
timestamp 1745462530
transform 1 0 3324 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_10068
timestamp 1745462530
transform 1 0 3308 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_10069
timestamp 1745462530
transform 1 0 3268 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_10070
timestamp 1745462530
transform 1 0 3260 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_10071
timestamp 1745462530
transform 1 0 3260 0 1 1075
box -3 -3 3 3
use M3_M2  M3_M2_10072
timestamp 1745462530
transform 1 0 2700 0 1 1075
box -3 -3 3 3
use M3_M2  M3_M2_10073
timestamp 1745462530
transform 1 0 2324 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_10074
timestamp 1745462530
transform 1 0 2324 0 1 2255
box -3 -3 3 3
use M3_M2  M3_M2_10075
timestamp 1745462530
transform 1 0 2228 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_10076
timestamp 1745462530
transform 1 0 1964 0 1 2255
box -3 -3 3 3
use M3_M2  M3_M2_10077
timestamp 1745462530
transform 1 0 1964 0 1 1075
box -3 -3 3 3
use M3_M2  M3_M2_10078
timestamp 1745462530
transform 1 0 1964 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_10079
timestamp 1745462530
transform 1 0 1604 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_10080
timestamp 1745462530
transform 1 0 980 0 1 2255
box -3 -3 3 3
use M3_M2  M3_M2_10081
timestamp 1745462530
transform 1 0 980 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_10082
timestamp 1745462530
transform 1 0 3252 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_10083
timestamp 1745462530
transform 1 0 3212 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_10084
timestamp 1745462530
transform 1 0 3164 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_10085
timestamp 1745462530
transform 1 0 3156 0 1 1895
box -3 -3 3 3
use M3_M2  M3_M2_10086
timestamp 1745462530
transform 1 0 2956 0 1 1895
box -3 -3 3 3
use M3_M2  M3_M2_10087
timestamp 1745462530
transform 1 0 2308 0 1 1895
box -3 -3 3 3
use M3_M2  M3_M2_10088
timestamp 1745462530
transform 1 0 3228 0 1 1295
box -3 -3 3 3
use M3_M2  M3_M2_10089
timestamp 1745462530
transform 1 0 2932 0 1 2455
box -3 -3 3 3
use M3_M2  M3_M2_10090
timestamp 1745462530
transform 1 0 2684 0 1 1295
box -3 -3 3 3
use M3_M2  M3_M2_10091
timestamp 1745462530
transform 1 0 2300 0 1 1295
box -3 -3 3 3
use M3_M2  M3_M2_10092
timestamp 1745462530
transform 1 0 2284 0 1 2465
box -3 -3 3 3
use M3_M2  M3_M2_10093
timestamp 1745462530
transform 1 0 2252 0 1 1295
box -3 -3 3 3
use M3_M2  M3_M2_10094
timestamp 1745462530
transform 1 0 2244 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_10095
timestamp 1745462530
transform 1 0 1276 0 1 2465
box -3 -3 3 3
use M3_M2  M3_M2_10096
timestamp 1745462530
transform 1 0 1268 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_10097
timestamp 1745462530
transform 1 0 1268 0 1 2285
box -3 -3 3 3
use M3_M2  M3_M2_10098
timestamp 1745462530
transform 1 0 1268 0 1 2005
box -3 -3 3 3
use M3_M2  M3_M2_10099
timestamp 1745462530
transform 1 0 1268 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_10100
timestamp 1745462530
transform 1 0 1252 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_10101
timestamp 1745462530
transform 1 0 1220 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_10102
timestamp 1745462530
transform 1 0 1220 0 1 2285
box -3 -3 3 3
use M3_M2  M3_M2_10103
timestamp 1745462530
transform 1 0 1220 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_10104
timestamp 1745462530
transform 1 0 1108 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_10105
timestamp 1745462530
transform 1 0 1060 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_10106
timestamp 1745462530
transform 1 0 3204 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_10107
timestamp 1745462530
transform 1 0 2972 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_10108
timestamp 1745462530
transform 1 0 2940 0 1 2175
box -3 -3 3 3
use M3_M2  M3_M2_10109
timestamp 1745462530
transform 1 0 2924 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_10110
timestamp 1745462530
transform 1 0 2900 0 1 2295
box -3 -3 3 3
use M3_M2  M3_M2_10111
timestamp 1745462530
transform 1 0 2900 0 1 2175
box -3 -3 3 3
use M3_M2  M3_M2_10112
timestamp 1745462530
transform 1 0 2876 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_10113
timestamp 1745462530
transform 1 0 2444 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_10114
timestamp 1745462530
transform 1 0 2380 0 1 2295
box -3 -3 3 3
use M3_M2  M3_M2_10115
timestamp 1745462530
transform 1 0 2052 0 1 2275
box -3 -3 3 3
use M3_M2  M3_M2_10116
timestamp 1745462530
transform 1 0 1236 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_10117
timestamp 1745462530
transform 1 0 1236 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_10118
timestamp 1745462530
transform 1 0 1148 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_10119
timestamp 1745462530
transform 1 0 956 0 1 2185
box -3 -3 3 3
use M3_M2  M3_M2_10120
timestamp 1745462530
transform 1 0 884 0 1 2275
box -3 -3 3 3
use M3_M2  M3_M2_10121
timestamp 1745462530
transform 1 0 876 0 1 2185
box -3 -3 3 3
use M3_M2  M3_M2_10122
timestamp 1745462530
transform 1 0 2988 0 1 1065
box -3 -3 3 3
use M3_M2  M3_M2_10123
timestamp 1745462530
transform 1 0 2956 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_10124
timestamp 1745462530
transform 1 0 2828 0 1 1055
box -3 -3 3 3
use M3_M2  M3_M2_10125
timestamp 1745462530
transform 1 0 2796 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_10126
timestamp 1745462530
transform 1 0 2836 0 1 535
box -3 -3 3 3
use M3_M2  M3_M2_10127
timestamp 1745462530
transform 1 0 2716 0 1 535
box -3 -3 3 3
use M3_M2  M3_M2_10128
timestamp 1745462530
transform 1 0 2724 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_10129
timestamp 1745462530
transform 1 0 2708 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_10130
timestamp 1745462530
transform 1 0 2676 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_10131
timestamp 1745462530
transform 1 0 2668 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_10132
timestamp 1745462530
transform 1 0 2404 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_10133
timestamp 1745462530
transform 1 0 2292 0 1 1375
box -3 -3 3 3
use M3_M2  M3_M2_10134
timestamp 1745462530
transform 1 0 2276 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_10135
timestamp 1745462530
transform 1 0 2236 0 1 1375
box -3 -3 3 3
use M3_M2  M3_M2_10136
timestamp 1745462530
transform 1 0 3532 0 1 2055
box -3 -3 3 3
use M3_M2  M3_M2_10137
timestamp 1745462530
transform 1 0 3500 0 1 2055
box -3 -3 3 3
use M3_M2  M3_M2_10138
timestamp 1745462530
transform 1 0 3548 0 1 2475
box -3 -3 3 3
use M3_M2  M3_M2_10139
timestamp 1745462530
transform 1 0 3516 0 1 2475
box -3 -3 3 3
use M3_M2  M3_M2_10140
timestamp 1745462530
transform 1 0 3556 0 1 2695
box -3 -3 3 3
use M3_M2  M3_M2_10141
timestamp 1745462530
transform 1 0 3524 0 1 2695
box -3 -3 3 3
use M3_M2  M3_M2_10142
timestamp 1745462530
transform 1 0 3588 0 1 2625
box -3 -3 3 3
use M3_M2  M3_M2_10143
timestamp 1745462530
transform 1 0 3516 0 1 2625
box -3 -3 3 3
use M3_M2  M3_M2_10144
timestamp 1745462530
transform 1 0 3540 0 1 2615
box -3 -3 3 3
use M3_M2  M3_M2_10145
timestamp 1745462530
transform 1 0 3524 0 1 2615
box -3 -3 3 3
use M3_M2  M3_M2_10146
timestamp 1745462530
transform 1 0 3540 0 1 2565
box -3 -3 3 3
use M3_M2  M3_M2_10147
timestamp 1745462530
transform 1 0 3516 0 1 2565
box -3 -3 3 3
use M3_M2  M3_M2_10148
timestamp 1745462530
transform 1 0 2916 0 1 2335
box -3 -3 3 3
use M3_M2  M3_M2_10149
timestamp 1745462530
transform 1 0 2908 0 1 2365
box -3 -3 3 3
use M3_M2  M3_M2_10150
timestamp 1745462530
transform 1 0 2876 0 1 2335
box -3 -3 3 3
use M3_M2  M3_M2_10151
timestamp 1745462530
transform 1 0 2652 0 1 2365
box -3 -3 3 3
use M3_M2  M3_M2_10152
timestamp 1745462530
transform 1 0 2628 0 1 2365
box -3 -3 3 3
use M3_M2  M3_M2_10153
timestamp 1745462530
transform 1 0 2612 0 1 2365
box -3 -3 3 3
use M3_M2  M3_M2_10154
timestamp 1745462530
transform 1 0 2284 0 1 2365
box -3 -3 3 3
use M3_M2  M3_M2_10155
timestamp 1745462530
transform 1 0 2692 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_10156
timestamp 1745462530
transform 1 0 2284 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_10157
timestamp 1745462530
transform 1 0 2228 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_10158
timestamp 1745462530
transform 1 0 2084 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_10159
timestamp 1745462530
transform 1 0 2724 0 1 2545
box -3 -3 3 3
use M3_M2  M3_M2_10160
timestamp 1745462530
transform 1 0 2636 0 1 2545
box -3 -3 3 3
use M3_M2  M3_M2_10161
timestamp 1745462530
transform 1 0 2332 0 1 2545
box -3 -3 3 3
use M3_M2  M3_M2_10162
timestamp 1745462530
transform 1 0 2212 0 1 2535
box -3 -3 3 3
use M3_M2  M3_M2_10163
timestamp 1745462530
transform 1 0 2692 0 1 2405
box -3 -3 3 3
use M3_M2  M3_M2_10164
timestamp 1745462530
transform 1 0 2556 0 1 2405
box -3 -3 3 3
use M3_M2  M3_M2_10165
timestamp 1745462530
transform 1 0 2332 0 1 2405
box -3 -3 3 3
use M3_M2  M3_M2_10166
timestamp 1745462530
transform 1 0 2188 0 1 2405
box -3 -3 3 3
use M3_M2  M3_M2_10167
timestamp 1745462530
transform 1 0 2652 0 1 2435
box -3 -3 3 3
use M3_M2  M3_M2_10168
timestamp 1745462530
transform 1 0 2532 0 1 2435
box -3 -3 3 3
use M3_M2  M3_M2_10169
timestamp 1745462530
transform 1 0 2388 0 1 2435
box -3 -3 3 3
use M3_M2  M3_M2_10170
timestamp 1745462530
transform 1 0 2388 0 1 2375
box -3 -3 3 3
use M3_M2  M3_M2_10171
timestamp 1745462530
transform 1 0 2140 0 1 2375
box -3 -3 3 3
use M3_M2  M3_M2_10172
timestamp 1745462530
transform 1 0 3508 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_10173
timestamp 1745462530
transform 1 0 3012 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_10174
timestamp 1745462530
transform 1 0 3556 0 1 2085
box -3 -3 3 3
use M3_M2  M3_M2_10175
timestamp 1745462530
transform 1 0 3508 0 1 2085
box -3 -3 3 3
use M3_M2  M3_M2_10176
timestamp 1745462530
transform 1 0 3684 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_10177
timestamp 1745462530
transform 1 0 3524 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_10178
timestamp 1745462530
transform 1 0 3772 0 1 1855
box -3 -3 3 3
use M3_M2  M3_M2_10179
timestamp 1745462530
transform 1 0 3708 0 1 1855
box -3 -3 3 3
use M3_M2  M3_M2_10180
timestamp 1745462530
transform 1 0 3756 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_10181
timestamp 1745462530
transform 1 0 3724 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_10182
timestamp 1745462530
transform 1 0 1508 0 1 2185
box -3 -3 3 3
use M3_M2  M3_M2_10183
timestamp 1745462530
transform 1 0 796 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_10184
timestamp 1745462530
transform 1 0 788 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_10185
timestamp 1745462530
transform 1 0 772 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_10186
timestamp 1745462530
transform 1 0 748 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_10187
timestamp 1745462530
transform 1 0 724 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_10188
timestamp 1745462530
transform 1 0 764 0 1 2645
box -3 -3 3 3
use M3_M2  M3_M2_10189
timestamp 1745462530
transform 1 0 684 0 1 2645
box -3 -3 3 3
use M3_M2  M3_M2_10190
timestamp 1745462530
transform 1 0 660 0 1 2745
box -3 -3 3 3
use M3_M2  M3_M2_10191
timestamp 1745462530
transform 1 0 644 0 1 2745
box -3 -3 3 3
use M3_M2  M3_M2_10192
timestamp 1745462530
transform 1 0 716 0 1 2685
box -3 -3 3 3
use M3_M2  M3_M2_10193
timestamp 1745462530
transform 1 0 692 0 1 2685
box -3 -3 3 3
use M3_M2  M3_M2_10194
timestamp 1745462530
transform 1 0 2180 0 1 2235
box -3 -3 3 3
use M3_M2  M3_M2_10195
timestamp 1745462530
transform 1 0 996 0 1 2235
box -3 -3 3 3
use M3_M2  M3_M2_10196
timestamp 1745462530
transform 1 0 956 0 1 2235
box -3 -3 3 3
use M3_M2  M3_M2_10197
timestamp 1745462530
transform 1 0 2180 0 1 2065
box -3 -3 3 3
use M3_M2  M3_M2_10198
timestamp 1745462530
transform 1 0 2028 0 1 2065
box -3 -3 3 3
use M3_M2  M3_M2_10199
timestamp 1745462530
transform 1 0 2028 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_10200
timestamp 1745462530
transform 1 0 1092 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_10201
timestamp 1745462530
transform 1 0 1092 0 1 1265
box -3 -3 3 3
use M3_M2  M3_M2_10202
timestamp 1745462530
transform 1 0 1036 0 1 1265
box -3 -3 3 3
use M3_M2  M3_M2_10203
timestamp 1745462530
transform 1 0 964 0 1 1005
box -3 -3 3 3
use M3_M2  M3_M2_10204
timestamp 1745462530
transform 1 0 876 0 1 1265
box -3 -3 3 3
use M3_M2  M3_M2_10205
timestamp 1745462530
transform 1 0 868 0 1 1005
box -3 -3 3 3
use M3_M2  M3_M2_10206
timestamp 1745462530
transform 1 0 1556 0 1 2405
box -3 -3 3 3
use M3_M2  M3_M2_10207
timestamp 1745462530
transform 1 0 1468 0 1 2405
box -3 -3 3 3
use M3_M2  M3_M2_10208
timestamp 1745462530
transform 1 0 1452 0 1 2405
box -3 -3 3 3
use M3_M2  M3_M2_10209
timestamp 1745462530
transform 1 0 1404 0 1 2405
box -3 -3 3 3
use M3_M2  M3_M2_10210
timestamp 1745462530
transform 1 0 1460 0 1 2365
box -3 -3 3 3
use M3_M2  M3_M2_10211
timestamp 1745462530
transform 1 0 1412 0 1 2365
box -3 -3 3 3
use M3_M2  M3_M2_10212
timestamp 1745462530
transform 1 0 1428 0 1 2315
box -3 -3 3 3
use M3_M2  M3_M2_10213
timestamp 1745462530
transform 1 0 1364 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_10214
timestamp 1745462530
transform 1 0 2212 0 1 2455
box -3 -3 3 3
use M3_M2  M3_M2_10215
timestamp 1745462530
transform 1 0 2188 0 1 2355
box -3 -3 3 3
use M3_M2  M3_M2_10216
timestamp 1745462530
transform 1 0 2164 0 1 2455
box -3 -3 3 3
use M3_M2  M3_M2_10217
timestamp 1745462530
transform 1 0 2164 0 1 2355
box -3 -3 3 3
use M3_M2  M3_M2_10218
timestamp 1745462530
transform 1 0 2100 0 1 2355
box -3 -3 3 3
use M3_M2  M3_M2_10219
timestamp 1745462530
transform 1 0 2060 0 1 2355
box -3 -3 3 3
use M3_M2  M3_M2_10220
timestamp 1745462530
transform 1 0 1116 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_10221
timestamp 1745462530
transform 1 0 772 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_10222
timestamp 1745462530
transform 1 0 1300 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_10223
timestamp 1745462530
transform 1 0 1276 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_10224
timestamp 1745462530
transform 1 0 1260 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_10225
timestamp 1745462530
transform 1 0 1164 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_10226
timestamp 1745462530
transform 1 0 1236 0 1 975
box -3 -3 3 3
use M3_M2  M3_M2_10227
timestamp 1745462530
transform 1 0 1172 0 1 975
box -3 -3 3 3
use M3_M2  M3_M2_10228
timestamp 1745462530
transform 1 0 1156 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_10229
timestamp 1745462530
transform 1 0 1108 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_10230
timestamp 1745462530
transform 1 0 1260 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_10231
timestamp 1745462530
transform 1 0 1196 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_10232
timestamp 1745462530
transform 1 0 2100 0 1 1675
box -3 -3 3 3
use M3_M2  M3_M2_10233
timestamp 1745462530
transform 1 0 2044 0 1 1535
box -3 -3 3 3
use M3_M2  M3_M2_10234
timestamp 1745462530
transform 1 0 2036 0 1 1675
box -3 -3 3 3
use M3_M2  M3_M2_10235
timestamp 1745462530
transform 1 0 1996 0 1 1535
box -3 -3 3 3
use M3_M2  M3_M2_10236
timestamp 1745462530
transform 1 0 1996 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_10237
timestamp 1745462530
transform 1 0 1972 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_10238
timestamp 1745462530
transform 1 0 1972 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_10239
timestamp 1745462530
transform 1 0 1636 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_10240
timestamp 1745462530
transform 1 0 1612 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_10241
timestamp 1745462530
transform 1 0 1572 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_10242
timestamp 1745462530
transform 1 0 1396 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_10243
timestamp 1745462530
transform 1 0 1380 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_10244
timestamp 1745462530
transform 1 0 1284 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_10245
timestamp 1745462530
transform 1 0 1284 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_10246
timestamp 1745462530
transform 1 0 1220 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_10247
timestamp 1745462530
transform 1 0 1220 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_10248
timestamp 1745462530
transform 1 0 1164 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_10249
timestamp 1745462530
transform 1 0 820 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_10250
timestamp 1745462530
transform 1 0 772 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_10251
timestamp 1745462530
transform 1 0 772 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_10252
timestamp 1745462530
transform 1 0 740 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_10253
timestamp 1745462530
transform 1 0 804 0 1 845
box -3 -3 3 3
use M3_M2  M3_M2_10254
timestamp 1745462530
transform 1 0 748 0 1 845
box -3 -3 3 3
use M3_M2  M3_M2_10255
timestamp 1745462530
transform 1 0 708 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_10256
timestamp 1745462530
transform 1 0 540 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_10257
timestamp 1745462530
transform 1 0 2284 0 1 2865
box -3 -3 3 3
use M3_M2  M3_M2_10258
timestamp 1745462530
transform 1 0 2204 0 1 2865
box -3 -3 3 3
use M3_M2  M3_M2_10259
timestamp 1745462530
transform 1 0 2108 0 1 2865
box -3 -3 3 3
use M3_M2  M3_M2_10260
timestamp 1745462530
transform 1 0 2332 0 1 2845
box -3 -3 3 3
use M3_M2  M3_M2_10261
timestamp 1745462530
transform 1 0 2180 0 1 2845
box -3 -3 3 3
use M3_M2  M3_M2_10262
timestamp 1745462530
transform 1 0 2148 0 1 2845
box -3 -3 3 3
use M3_M2  M3_M2_10263
timestamp 1745462530
transform 1 0 2100 0 1 2945
box -3 -3 3 3
use M3_M2  M3_M2_10264
timestamp 1745462530
transform 1 0 2100 0 1 2845
box -3 -3 3 3
use M3_M2  M3_M2_10265
timestamp 1745462530
transform 1 0 2036 0 1 2945
box -3 -3 3 3
use M3_M2  M3_M2_10266
timestamp 1745462530
transform 1 0 2252 0 1 2885
box -3 -3 3 3
use M3_M2  M3_M2_10267
timestamp 1745462530
transform 1 0 2172 0 1 2885
box -3 -3 3 3
use M3_M2  M3_M2_10268
timestamp 1745462530
transform 1 0 2244 0 1 3045
box -3 -3 3 3
use M3_M2  M3_M2_10269
timestamp 1745462530
transform 1 0 2076 0 1 3045
box -3 -3 3 3
use M3_M2  M3_M2_10270
timestamp 1745462530
transform 1 0 1132 0 1 3185
box -3 -3 3 3
use M3_M2  M3_M2_10271
timestamp 1745462530
transform 1 0 988 0 1 3185
box -3 -3 3 3
use M3_M2  M3_M2_10272
timestamp 1745462530
transform 1 0 516 0 1 3215
box -3 -3 3 3
use M3_M2  M3_M2_10273
timestamp 1745462530
transform 1 0 452 0 1 3215
box -3 -3 3 3
use M3_M2  M3_M2_10274
timestamp 1745462530
transform 1 0 356 0 1 3215
box -3 -3 3 3
use M3_M2  M3_M2_10275
timestamp 1745462530
transform 1 0 244 0 1 3215
box -3 -3 3 3
use M3_M2  M3_M2_10276
timestamp 1745462530
transform 1 0 252 0 1 3115
box -3 -3 3 3
use M3_M2  M3_M2_10277
timestamp 1745462530
transform 1 0 220 0 1 3115
box -3 -3 3 3
use M3_M2  M3_M2_10278
timestamp 1745462530
transform 1 0 1532 0 1 3105
box -3 -3 3 3
use M3_M2  M3_M2_10279
timestamp 1745462530
transform 1 0 1268 0 1 3165
box -3 -3 3 3
use M3_M2  M3_M2_10280
timestamp 1745462530
transform 1 0 1268 0 1 3105
box -3 -3 3 3
use M3_M2  M3_M2_10281
timestamp 1745462530
transform 1 0 1100 0 1 3165
box -3 -3 3 3
use M3_M2  M3_M2_10282
timestamp 1745462530
transform 1 0 1316 0 1 2805
box -3 -3 3 3
use M3_M2  M3_M2_10283
timestamp 1745462530
transform 1 0 1276 0 1 2805
box -3 -3 3 3
use M3_M2  M3_M2_10284
timestamp 1745462530
transform 1 0 1052 0 1 3445
box -3 -3 3 3
use M3_M2  M3_M2_10285
timestamp 1745462530
transform 1 0 956 0 1 3445
box -3 -3 3 3
use M3_M2  M3_M2_10286
timestamp 1745462530
transform 1 0 1084 0 1 3415
box -3 -3 3 3
use M3_M2  M3_M2_10287
timestamp 1745462530
transform 1 0 964 0 1 3415
box -3 -3 3 3
use M3_M2  M3_M2_10288
timestamp 1745462530
transform 1 0 1132 0 1 3445
box -3 -3 3 3
use M3_M2  M3_M2_10289
timestamp 1745462530
transform 1 0 1076 0 1 3445
box -3 -3 3 3
use M3_M2  M3_M2_10290
timestamp 1745462530
transform 1 0 1220 0 1 3505
box -3 -3 3 3
use M3_M2  M3_M2_10291
timestamp 1745462530
transform 1 0 1044 0 1 3505
box -3 -3 3 3
use M3_M2  M3_M2_10292
timestamp 1745462530
transform 1 0 1508 0 1 3605
box -3 -3 3 3
use M3_M2  M3_M2_10293
timestamp 1745462530
transform 1 0 1404 0 1 3605
box -3 -3 3 3
use M3_M2  M3_M2_10294
timestamp 1745462530
transform 1 0 1556 0 1 3555
box -3 -3 3 3
use M3_M2  M3_M2_10295
timestamp 1745462530
transform 1 0 1492 0 1 3555
box -3 -3 3 3
use M3_M2  M3_M2_10296
timestamp 1745462530
transform 1 0 1444 0 1 3555
box -3 -3 3 3
use M3_M2  M3_M2_10297
timestamp 1745462530
transform 1 0 1340 0 1 3555
box -3 -3 3 3
use M3_M2  M3_M2_10298
timestamp 1745462530
transform 1 0 1276 0 1 3555
box -3 -3 3 3
use M3_M2  M3_M2_10299
timestamp 1745462530
transform 1 0 1524 0 1 3655
box -3 -3 3 3
use M3_M2  M3_M2_10300
timestamp 1745462530
transform 1 0 1300 0 1 3655
box -3 -3 3 3
use M3_M2  M3_M2_10301
timestamp 1745462530
transform 1 0 1428 0 1 3715
box -3 -3 3 3
use M3_M2  M3_M2_10302
timestamp 1745462530
transform 1 0 1364 0 1 3775
box -3 -3 3 3
use M3_M2  M3_M2_10303
timestamp 1745462530
transform 1 0 1364 0 1 3715
box -3 -3 3 3
use M3_M2  M3_M2_10304
timestamp 1745462530
transform 1 0 1308 0 1 3775
box -3 -3 3 3
use M3_M2  M3_M2_10305
timestamp 1745462530
transform 1 0 1228 0 1 3775
box -3 -3 3 3
use M3_M2  M3_M2_10306
timestamp 1745462530
transform 1 0 1468 0 1 3595
box -3 -3 3 3
use M3_M2  M3_M2_10307
timestamp 1745462530
transform 1 0 1412 0 1 3595
box -3 -3 3 3
use M3_M2  M3_M2_10308
timestamp 1745462530
transform 1 0 1580 0 1 3705
box -3 -3 3 3
use M3_M2  M3_M2_10309
timestamp 1745462530
transform 1 0 1484 0 1 3725
box -3 -3 3 3
use M3_M2  M3_M2_10310
timestamp 1745462530
transform 1 0 1436 0 1 3725
box -3 -3 3 3
use M3_M2  M3_M2_10311
timestamp 1745462530
transform 1 0 1436 0 1 3495
box -3 -3 3 3
use M3_M2  M3_M2_10312
timestamp 1745462530
transform 1 0 1396 0 1 3495
box -3 -3 3 3
use M3_M2  M3_M2_10313
timestamp 1745462530
transform 1 0 1356 0 1 3725
box -3 -3 3 3
use M3_M2  M3_M2_10314
timestamp 1745462530
transform 1 0 1356 0 1 3755
box -3 -3 3 3
use M3_M2  M3_M2_10315
timestamp 1745462530
transform 1 0 1260 0 1 3755
box -3 -3 3 3
use M3_M2  M3_M2_10316
timestamp 1745462530
transform 1 0 1612 0 1 3745
box -3 -3 3 3
use M3_M2  M3_M2_10317
timestamp 1745462530
transform 1 0 1316 0 1 3745
box -3 -3 3 3
use M3_M2  M3_M2_10318
timestamp 1745462530
transform 1 0 1292 0 1 3745
box -3 -3 3 3
use M3_M2  M3_M2_10319
timestamp 1745462530
transform 1 0 1460 0 1 3535
box -3 -3 3 3
use M3_M2  M3_M2_10320
timestamp 1745462530
transform 1 0 1420 0 1 3535
box -3 -3 3 3
use M3_M2  M3_M2_10321
timestamp 1745462530
transform 1 0 1492 0 1 3515
box -3 -3 3 3
use M3_M2  M3_M2_10322
timestamp 1745462530
transform 1 0 1476 0 1 3515
box -3 -3 3 3
use M3_M2  M3_M2_10323
timestamp 1745462530
transform 1 0 1476 0 1 3495
box -3 -3 3 3
use M3_M2  M3_M2_10324
timestamp 1745462530
transform 1 0 1404 0 1 3585
box -3 -3 3 3
use M3_M2  M3_M2_10325
timestamp 1745462530
transform 1 0 1404 0 1 3485
box -3 -3 3 3
use M3_M2  M3_M2_10326
timestamp 1745462530
transform 1 0 1204 0 1 3585
box -3 -3 3 3
use M3_M2  M3_M2_10327
timestamp 1745462530
transform 1 0 1516 0 1 3465
box -3 -3 3 3
use M3_M2  M3_M2_10328
timestamp 1745462530
transform 1 0 1380 0 1 3365
box -3 -3 3 3
use M3_M2  M3_M2_10329
timestamp 1745462530
transform 1 0 1364 0 1 3465
box -3 -3 3 3
use M3_M2  M3_M2_10330
timestamp 1745462530
transform 1 0 1316 0 1 3365
box -3 -3 3 3
use M3_M2  M3_M2_10331
timestamp 1745462530
transform 1 0 1508 0 1 3375
box -3 -3 3 3
use M3_M2  M3_M2_10332
timestamp 1745462530
transform 1 0 1476 0 1 3375
box -3 -3 3 3
use M3_M2  M3_M2_10333
timestamp 1745462530
transform 1 0 1484 0 1 3305
box -3 -3 3 3
use M3_M2  M3_M2_10334
timestamp 1745462530
transform 1 0 1420 0 1 3305
box -3 -3 3 3
use M3_M2  M3_M2_10335
timestamp 1745462530
transform 1 0 1500 0 1 3685
box -3 -3 3 3
use M3_M2  M3_M2_10336
timestamp 1745462530
transform 1 0 1396 0 1 3355
box -3 -3 3 3
use M3_M2  M3_M2_10337
timestamp 1745462530
transform 1 0 1356 0 1 3355
box -3 -3 3 3
use M3_M2  M3_M2_10338
timestamp 1745462530
transform 1 0 1348 0 1 3685
box -3 -3 3 3
use M3_M2  M3_M2_10339
timestamp 1745462530
transform 1 0 1564 0 1 3445
box -3 -3 3 3
use M3_M2  M3_M2_10340
timestamp 1745462530
transform 1 0 1420 0 1 3445
box -3 -3 3 3
use M3_M2  M3_M2_10341
timestamp 1745462530
transform 1 0 1612 0 1 3375
box -3 -3 3 3
use M3_M2  M3_M2_10342
timestamp 1745462530
transform 1 0 1580 0 1 3375
box -3 -3 3 3
use M3_M2  M3_M2_10343
timestamp 1745462530
transform 1 0 996 0 1 3755
box -3 -3 3 3
use M3_M2  M3_M2_10344
timestamp 1745462530
transform 1 0 916 0 1 3755
box -3 -3 3 3
use M3_M2  M3_M2_10345
timestamp 1745462530
transform 1 0 1156 0 1 3795
box -3 -3 3 3
use M3_M2  M3_M2_10346
timestamp 1745462530
transform 1 0 1044 0 1 3795
box -3 -3 3 3
use M3_M2  M3_M2_10347
timestamp 1745462530
transform 1 0 3132 0 1 3825
box -3 -3 3 3
use M3_M2  M3_M2_10348
timestamp 1745462530
transform 1 0 3068 0 1 3825
box -3 -3 3 3
use M3_M2  M3_M2_10349
timestamp 1745462530
transform 1 0 3356 0 1 3805
box -3 -3 3 3
use M3_M2  M3_M2_10350
timestamp 1745462530
transform 1 0 3300 0 1 3805
box -3 -3 3 3
use M3_M2  M3_M2_10351
timestamp 1745462530
transform 1 0 2484 0 1 3945
box -3 -3 3 3
use M3_M2  M3_M2_10352
timestamp 1745462530
transform 1 0 2396 0 1 3945
box -3 -3 3 3
use M3_M2  M3_M2_10353
timestamp 1745462530
transform 1 0 2852 0 1 3975
box -3 -3 3 3
use M3_M2  M3_M2_10354
timestamp 1745462530
transform 1 0 2772 0 1 3975
box -3 -3 3 3
use M3_M2  M3_M2_10355
timestamp 1745462530
transform 1 0 3868 0 1 3795
box -3 -3 3 3
use M3_M2  M3_M2_10356
timestamp 1745462530
transform 1 0 3644 0 1 3795
box -3 -3 3 3
use M3_M2  M3_M2_10357
timestamp 1745462530
transform 1 0 3684 0 1 4005
box -3 -3 3 3
use M3_M2  M3_M2_10358
timestamp 1745462530
transform 1 0 3612 0 1 4005
box -3 -3 3 3
use M3_M2  M3_M2_10359
timestamp 1745462530
transform 1 0 3756 0 1 3825
box -3 -3 3 3
use M3_M2  M3_M2_10360
timestamp 1745462530
transform 1 0 3604 0 1 3825
box -3 -3 3 3
use M3_M2  M3_M2_10361
timestamp 1745462530
transform 1 0 3316 0 1 4185
box -3 -3 3 3
use M3_M2  M3_M2_10362
timestamp 1745462530
transform 1 0 3244 0 1 4185
box -3 -3 3 3
use M3_M2  M3_M2_10363
timestamp 1745462530
transform 1 0 2484 0 1 4045
box -3 -3 3 3
use M3_M2  M3_M2_10364
timestamp 1745462530
transform 1 0 2388 0 1 4045
box -3 -3 3 3
use M3_M2  M3_M2_10365
timestamp 1745462530
transform 1 0 2276 0 1 3975
box -3 -3 3 3
use M3_M2  M3_M2_10366
timestamp 1745462530
transform 1 0 2228 0 1 3975
box -3 -3 3 3
use M3_M2  M3_M2_10367
timestamp 1745462530
transform 1 0 2836 0 1 4115
box -3 -3 3 3
use M3_M2  M3_M2_10368
timestamp 1745462530
transform 1 0 2756 0 1 4115
box -3 -3 3 3
use M3_M2  M3_M2_10369
timestamp 1745462530
transform 1 0 3116 0 1 4185
box -3 -3 3 3
use M3_M2  M3_M2_10370
timestamp 1745462530
transform 1 0 3028 0 1 4185
box -3 -3 3 3
use M3_M2  M3_M2_10371
timestamp 1745462530
transform 1 0 3564 0 1 4185
box -3 -3 3 3
use M3_M2  M3_M2_10372
timestamp 1745462530
transform 1 0 3500 0 1 4185
box -3 -3 3 3
use M3_M2  M3_M2_10373
timestamp 1745462530
transform 1 0 3660 0 1 3985
box -3 -3 3 3
use M3_M2  M3_M2_10374
timestamp 1745462530
transform 1 0 3516 0 1 3985
box -3 -3 3 3
use M3_M2  M3_M2_10375
timestamp 1745462530
transform 1 0 3220 0 1 4185
box -3 -3 3 3
use M3_M2  M3_M2_10376
timestamp 1745462530
transform 1 0 3188 0 1 4185
box -3 -3 3 3
use M3_M2  M3_M2_10377
timestamp 1745462530
transform 1 0 2188 0 1 4145
box -3 -3 3 3
use M3_M2  M3_M2_10378
timestamp 1745462530
transform 1 0 2172 0 1 4145
box -3 -3 3 3
use M3_M2  M3_M2_10379
timestamp 1745462530
transform 1 0 2164 0 1 4195
box -3 -3 3 3
use M3_M2  M3_M2_10380
timestamp 1745462530
transform 1 0 2084 0 1 4205
box -3 -3 3 3
use M3_M2  M3_M2_10381
timestamp 1745462530
transform 1 0 2756 0 1 4185
box -3 -3 3 3
use M3_M2  M3_M2_10382
timestamp 1745462530
transform 1 0 2660 0 1 4185
box -3 -3 3 3
use M3_M2  M3_M2_10383
timestamp 1745462530
transform 1 0 2996 0 1 4105
box -3 -3 3 3
use M3_M2  M3_M2_10384
timestamp 1745462530
transform 1 0 2956 0 1 4105
box -3 -3 3 3
use M3_M2  M3_M2_10385
timestamp 1745462530
transform 1 0 3868 0 1 4005
box -3 -3 3 3
use M3_M2  M3_M2_10386
timestamp 1745462530
transform 1 0 3780 0 1 4005
box -3 -3 3 3
use M3_M2  M3_M2_10387
timestamp 1745462530
transform 1 0 3948 0 1 4185
box -3 -3 3 3
use M3_M2  M3_M2_10388
timestamp 1745462530
transform 1 0 3868 0 1 4185
box -3 -3 3 3
use M3_M2  M3_M2_10389
timestamp 1745462530
transform 1 0 3788 0 1 3915
box -3 -3 3 3
use M3_M2  M3_M2_10390
timestamp 1745462530
transform 1 0 3700 0 1 3915
box -3 -3 3 3
use M3_M2  M3_M2_10391
timestamp 1745462530
transform 1 0 3756 0 1 4275
box -3 -3 3 3
use M3_M2  M3_M2_10392
timestamp 1745462530
transform 1 0 3700 0 1 4275
box -3 -3 3 3
use M3_M2  M3_M2_10393
timestamp 1745462530
transform 1 0 4308 0 1 3865
box -3 -3 3 3
use M3_M2  M3_M2_10394
timestamp 1745462530
transform 1 0 4228 0 1 3865
box -3 -3 3 3
use M3_M2  M3_M2_10395
timestamp 1745462530
transform 1 0 4316 0 1 3625
box -3 -3 3 3
use M3_M2  M3_M2_10396
timestamp 1745462530
transform 1 0 4244 0 1 3625
box -3 -3 3 3
use M3_M2  M3_M2_10397
timestamp 1745462530
transform 1 0 1996 0 1 3795
box -3 -3 3 3
use M3_M2  M3_M2_10398
timestamp 1745462530
transform 1 0 1948 0 1 3795
box -3 -3 3 3
use M3_M2  M3_M2_10399
timestamp 1745462530
transform 1 0 2692 0 1 3945
box -3 -3 3 3
use M3_M2  M3_M2_10400
timestamp 1745462530
transform 1 0 2628 0 1 3945
box -3 -3 3 3
use M3_M2  M3_M2_10401
timestamp 1745462530
transform 1 0 2940 0 1 3805
box -3 -3 3 3
use M3_M2  M3_M2_10402
timestamp 1745462530
transform 1 0 2868 0 1 3805
box -3 -3 3 3
use M3_M2  M3_M2_10403
timestamp 1745462530
transform 1 0 4188 0 1 3515
box -3 -3 3 3
use M3_M2  M3_M2_10404
timestamp 1745462530
transform 1 0 4084 0 1 3515
box -3 -3 3 3
use M3_M2  M3_M2_10405
timestamp 1745462530
transform 1 0 4140 0 1 3625
box -3 -3 3 3
use M3_M2  M3_M2_10406
timestamp 1745462530
transform 1 0 4060 0 1 3625
box -3 -3 3 3
use M3_M2  M3_M2_10407
timestamp 1745462530
transform 1 0 4308 0 1 3455
box -3 -3 3 3
use M3_M2  M3_M2_10408
timestamp 1745462530
transform 1 0 4148 0 1 3455
box -3 -3 3 3
use M3_M2  M3_M2_10409
timestamp 1745462530
transform 1 0 4076 0 1 3425
box -3 -3 3 3
use M3_M2  M3_M2_10410
timestamp 1745462530
transform 1 0 3980 0 1 3425
box -3 -3 3 3
use M3_M2  M3_M2_10411
timestamp 1745462530
transform 1 0 2020 0 1 3575
box -3 -3 3 3
use M3_M2  M3_M2_10412
timestamp 1745462530
transform 1 0 1964 0 1 3575
box -3 -3 3 3
use M3_M2  M3_M2_10413
timestamp 1745462530
transform 1 0 1964 0 1 3985
box -3 -3 3 3
use M3_M2  M3_M2_10414
timestamp 1745462530
transform 1 0 1940 0 1 3985
box -3 -3 3 3
use M3_M2  M3_M2_10415
timestamp 1745462530
transform 1 0 4316 0 1 3315
box -3 -3 3 3
use M3_M2  M3_M2_10416
timestamp 1745462530
transform 1 0 4236 0 1 3315
box -3 -3 3 3
use M3_M2  M3_M2_10417
timestamp 1745462530
transform 1 0 4316 0 1 3405
box -3 -3 3 3
use M3_M2  M3_M2_10418
timestamp 1745462530
transform 1 0 4236 0 1 3405
box -3 -3 3 3
use M3_M2  M3_M2_10419
timestamp 1745462530
transform 1 0 4124 0 1 3205
box -3 -3 3 3
use M3_M2  M3_M2_10420
timestamp 1745462530
transform 1 0 4052 0 1 3205
box -3 -3 3 3
use M3_M2  M3_M2_10421
timestamp 1745462530
transform 1 0 1676 0 1 3885
box -3 -3 3 3
use M3_M2  M3_M2_10422
timestamp 1745462530
transform 1 0 1564 0 1 3885
box -3 -3 3 3
use M3_M2  M3_M2_10423
timestamp 1745462530
transform 1 0 1652 0 1 3935
box -3 -3 3 3
use M3_M2  M3_M2_10424
timestamp 1745462530
transform 1 0 1436 0 1 3935
box -3 -3 3 3
use M3_M2  M3_M2_10425
timestamp 1745462530
transform 1 0 1700 0 1 3995
box -3 -3 3 3
use M3_M2  M3_M2_10426
timestamp 1745462530
transform 1 0 1548 0 1 3995
box -3 -3 3 3
use M3_M2  M3_M2_10427
timestamp 1745462530
transform 1 0 4308 0 1 3135
box -3 -3 3 3
use M3_M2  M3_M2_10428
timestamp 1745462530
transform 1 0 4228 0 1 3135
box -3 -3 3 3
use M3_M2  M3_M2_10429
timestamp 1745462530
transform 1 0 4308 0 1 3205
box -3 -3 3 3
use M3_M2  M3_M2_10430
timestamp 1745462530
transform 1 0 4236 0 1 3205
box -3 -3 3 3
use M3_M2  M3_M2_10431
timestamp 1745462530
transform 1 0 4140 0 1 3335
box -3 -3 3 3
use M3_M2  M3_M2_10432
timestamp 1745462530
transform 1 0 4052 0 1 3335
box -3 -3 3 3
use M3_M2  M3_M2_10433
timestamp 1745462530
transform 1 0 3932 0 1 3715
box -3 -3 3 3
use M3_M2  M3_M2_10434
timestamp 1745462530
transform 1 0 3836 0 1 3715
box -3 -3 3 3
use M3_M2  M3_M2_10435
timestamp 1745462530
transform 1 0 1572 0 1 3795
box -3 -3 3 3
use M3_M2  M3_M2_10436
timestamp 1745462530
transform 1 0 1508 0 1 3795
box -3 -3 3 3
use M3_M2  M3_M2_10437
timestamp 1745462530
transform 1 0 1604 0 1 3775
box -3 -3 3 3
use M3_M2  M3_M2_10438
timestamp 1745462530
transform 1 0 1396 0 1 3775
box -3 -3 3 3
use M3_M2  M3_M2_10439
timestamp 1745462530
transform 1 0 828 0 1 3535
box -3 -3 3 3
use M3_M2  M3_M2_10440
timestamp 1745462530
transform 1 0 740 0 1 3535
box -3 -3 3 3
use M3_M2  M3_M2_10441
timestamp 1745462530
transform 1 0 876 0 1 3605
box -3 -3 3 3
use M3_M2  M3_M2_10442
timestamp 1745462530
transform 1 0 812 0 1 3605
box -3 -3 3 3
use M3_M2  M3_M2_10443
timestamp 1745462530
transform 1 0 1012 0 1 3605
box -3 -3 3 3
use M3_M2  M3_M2_10444
timestamp 1745462530
transform 1 0 948 0 1 3605
box -3 -3 3 3
use M3_M2  M3_M2_10445
timestamp 1745462530
transform 1 0 860 0 1 3395
box -3 -3 3 3
use M3_M2  M3_M2_10446
timestamp 1745462530
transform 1 0 764 0 1 3395
box -3 -3 3 3
use M3_M2  M3_M2_10447
timestamp 1745462530
transform 1 0 1268 0 1 3205
box -3 -3 3 3
use M3_M2  M3_M2_10448
timestamp 1745462530
transform 1 0 1196 0 1 3205
box -3 -3 3 3
use M3_M2  M3_M2_10449
timestamp 1745462530
transform 1 0 1580 0 1 3115
box -3 -3 3 3
use M3_M2  M3_M2_10450
timestamp 1745462530
transform 1 0 1516 0 1 3115
box -3 -3 3 3
use M3_M2  M3_M2_10451
timestamp 1745462530
transform 1 0 1428 0 1 3205
box -3 -3 3 3
use M3_M2  M3_M2_10452
timestamp 1745462530
transform 1 0 1380 0 1 3195
box -3 -3 3 3
use M3_M2  M3_M2_10453
timestamp 1745462530
transform 1 0 1940 0 1 3095
box -3 -3 3 3
use M3_M2  M3_M2_10454
timestamp 1745462530
transform 1 0 1628 0 1 3095
box -3 -3 3 3
use M3_M2  M3_M2_10455
timestamp 1745462530
transform 1 0 1964 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_10456
timestamp 1745462530
transform 1 0 1892 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_10457
timestamp 1745462530
transform 1 0 2076 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_10458
timestamp 1745462530
transform 1 0 1988 0 1 2215
box -3 -3 3 3
use M3_M2  M3_M2_10459
timestamp 1745462530
transform 1 0 2052 0 1 2565
box -3 -3 3 3
use M3_M2  M3_M2_10460
timestamp 1745462530
transform 1 0 1908 0 1 2565
box -3 -3 3 3
use M3_M2  M3_M2_10461
timestamp 1745462530
transform 1 0 2108 0 1 2055
box -3 -3 3 3
use M3_M2  M3_M2_10462
timestamp 1745462530
transform 1 0 1892 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_10463
timestamp 1745462530
transform 1 0 1892 0 1 2055
box -3 -3 3 3
use M3_M2  M3_M2_10464
timestamp 1745462530
transform 1 0 1804 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_10465
timestamp 1745462530
transform 1 0 1772 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_10466
timestamp 1745462530
transform 1 0 1732 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_10467
timestamp 1745462530
transform 1 0 372 0 1 2535
box -3 -3 3 3
use M3_M2  M3_M2_10468
timestamp 1745462530
transform 1 0 308 0 1 2535
box -3 -3 3 3
use M3_M2  M3_M2_10469
timestamp 1745462530
transform 1 0 588 0 1 2485
box -3 -3 3 3
use M3_M2  M3_M2_10470
timestamp 1745462530
transform 1 0 548 0 1 2485
box -3 -3 3 3
use M3_M2  M3_M2_10471
timestamp 1745462530
transform 1 0 220 0 1 2545
box -3 -3 3 3
use M3_M2  M3_M2_10472
timestamp 1745462530
transform 1 0 140 0 1 2545
box -3 -3 3 3
use M3_M2  M3_M2_10473
timestamp 1745462530
transform 1 0 292 0 1 2185
box -3 -3 3 3
use M3_M2  M3_M2_10474
timestamp 1745462530
transform 1 0 260 0 1 2185
box -3 -3 3 3
use M3_M2  M3_M2_10475
timestamp 1745462530
transform 1 0 620 0 1 1895
box -3 -3 3 3
use M3_M2  M3_M2_10476
timestamp 1745462530
transform 1 0 580 0 1 1895
box -3 -3 3 3
use M3_M2  M3_M2_10477
timestamp 1745462530
transform 1 0 356 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_10478
timestamp 1745462530
transform 1 0 252 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_10479
timestamp 1745462530
transform 1 0 252 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_10480
timestamp 1745462530
transform 1 0 148 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_10481
timestamp 1745462530
transform 1 0 260 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_10482
timestamp 1745462530
transform 1 0 188 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_10483
timestamp 1745462530
transform 1 0 596 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_10484
timestamp 1745462530
transform 1 0 476 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_10485
timestamp 1745462530
transform 1 0 708 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_10486
timestamp 1745462530
transform 1 0 620 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_10487
timestamp 1745462530
transform 1 0 852 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_10488
timestamp 1745462530
transform 1 0 780 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_10489
timestamp 1745462530
transform 1 0 580 0 1 1335
box -3 -3 3 3
use M3_M2  M3_M2_10490
timestamp 1745462530
transform 1 0 500 0 1 1335
box -3 -3 3 3
use M3_M2  M3_M2_10491
timestamp 1745462530
transform 1 0 724 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_10492
timestamp 1745462530
transform 1 0 692 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_10493
timestamp 1745462530
transform 1 0 1500 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_10494
timestamp 1745462530
transform 1 0 1404 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_10495
timestamp 1745462530
transform 1 0 1772 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_10496
timestamp 1745462530
transform 1 0 1684 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_10497
timestamp 1745462530
transform 1 0 1660 0 1 405
box -3 -3 3 3
use M3_M2  M3_M2_10498
timestamp 1745462530
transform 1 0 1572 0 1 405
box -3 -3 3 3
use M3_M2  M3_M2_10499
timestamp 1745462530
transform 1 0 1740 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_10500
timestamp 1745462530
transform 1 0 1716 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_10501
timestamp 1745462530
transform 1 0 1844 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_10502
timestamp 1745462530
transform 1 0 1756 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_10503
timestamp 1745462530
transform 1 0 1844 0 1 1335
box -3 -3 3 3
use M3_M2  M3_M2_10504
timestamp 1745462530
transform 1 0 1764 0 1 1335
box -3 -3 3 3
use M3_M2  M3_M2_10505
timestamp 1745462530
transform 1 0 3124 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_10506
timestamp 1745462530
transform 1 0 3036 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_10507
timestamp 1745462530
transform 1 0 3028 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_10508
timestamp 1745462530
transform 1 0 2940 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_10509
timestamp 1745462530
transform 1 0 2988 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_10510
timestamp 1745462530
transform 1 0 2916 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_10511
timestamp 1745462530
transform 1 0 3028 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_10512
timestamp 1745462530
transform 1 0 2860 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_10513
timestamp 1745462530
transform 1 0 2916 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_10514
timestamp 1745462530
transform 1 0 2812 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_10515
timestamp 1745462530
transform 1 0 3372 0 1 205
box -3 -3 3 3
use M3_M2  M3_M2_10516
timestamp 1745462530
transform 1 0 3324 0 1 205
box -3 -3 3 3
use M3_M2  M3_M2_10517
timestamp 1745462530
transform 1 0 4060 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_10518
timestamp 1745462530
transform 1 0 3996 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_10519
timestamp 1745462530
transform 1 0 4220 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_10520
timestamp 1745462530
transform 1 0 4140 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_10521
timestamp 1745462530
transform 1 0 4116 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_10522
timestamp 1745462530
transform 1 0 3884 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_10523
timestamp 1745462530
transform 1 0 4188 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_10524
timestamp 1745462530
transform 1 0 4116 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_10525
timestamp 1745462530
transform 1 0 3988 0 1 1775
box -3 -3 3 3
use M3_M2  M3_M2_10526
timestamp 1745462530
transform 1 0 3836 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_10527
timestamp 1745462530
transform 1 0 4324 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_10528
timestamp 1745462530
transform 1 0 4188 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_10529
timestamp 1745462530
transform 1 0 4036 0 1 2005
box -3 -3 3 3
use M3_M2  M3_M2_10530
timestamp 1745462530
transform 1 0 3868 0 1 2005
box -3 -3 3 3
use M3_M2  M3_M2_10531
timestamp 1745462530
transform 1 0 3980 0 1 2205
box -3 -3 3 3
use M3_M2  M3_M2_10532
timestamp 1745462530
transform 1 0 3868 0 1 2205
box -3 -3 3 3
use M3_M2  M3_M2_10533
timestamp 1745462530
transform 1 0 3220 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_10534
timestamp 1745462530
transform 1 0 3124 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_10535
timestamp 1745462530
transform 1 0 3028 0 1 2235
box -3 -3 3 3
use M3_M2  M3_M2_10536
timestamp 1745462530
transform 1 0 2940 0 1 2235
box -3 -3 3 3
use M3_M2  M3_M2_10537
timestamp 1745462530
transform 1 0 4268 0 1 2735
box -3 -3 3 3
use M3_M2  M3_M2_10538
timestamp 1745462530
transform 1 0 4204 0 1 2735
box -3 -3 3 3
use M3_M2  M3_M2_10539
timestamp 1745462530
transform 1 0 4020 0 1 3025
box -3 -3 3 3
use M3_M2  M3_M2_10540
timestamp 1745462530
transform 1 0 3924 0 1 3025
box -3 -3 3 3
use M3_M2  M3_M2_10541
timestamp 1745462530
transform 1 0 4212 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_10542
timestamp 1745462530
transform 1 0 4092 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_10543
timestamp 1745462530
transform 1 0 4276 0 1 3025
box -3 -3 3 3
use M3_M2  M3_M2_10544
timestamp 1745462530
transform 1 0 4180 0 1 3025
box -3 -3 3 3
use M3_M2  M3_M2_10545
timestamp 1745462530
transform 1 0 4308 0 1 2545
box -3 -3 3 3
use M3_M2  M3_M2_10546
timestamp 1745462530
transform 1 0 4220 0 1 2545
box -3 -3 3 3
use M3_M2  M3_M2_10547
timestamp 1745462530
transform 1 0 4316 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_10548
timestamp 1745462530
transform 1 0 4236 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_10549
timestamp 1745462530
transform 1 0 2812 0 1 2835
box -3 -3 3 3
use M3_M2  M3_M2_10550
timestamp 1745462530
transform 1 0 2780 0 1 2835
box -3 -3 3 3
use M3_M2  M3_M2_10551
timestamp 1745462530
transform 1 0 1372 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_10552
timestamp 1745462530
transform 1 0 1308 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_10553
timestamp 1745462530
transform 1 0 1284 0 1 2765
box -3 -3 3 3
use M3_M2  M3_M2_10554
timestamp 1745462530
transform 1 0 1260 0 1 2765
box -3 -3 3 3
use M3_M2  M3_M2_10555
timestamp 1745462530
transform 1 0 1340 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_10556
timestamp 1745462530
transform 1 0 1236 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_10557
timestamp 1745462530
transform 1 0 300 0 1 2905
box -3 -3 3 3
use M3_M2  M3_M2_10558
timestamp 1745462530
transform 1 0 236 0 1 2905
box -3 -3 3 3
use M3_M2  M3_M2_10559
timestamp 1745462530
transform 1 0 1148 0 1 2885
box -3 -3 3 3
use M3_M2  M3_M2_10560
timestamp 1745462530
transform 1 0 964 0 1 2885
box -3 -3 3 3
use M3_M2  M3_M2_10561
timestamp 1745462530
transform 1 0 444 0 1 2405
box -3 -3 3 3
use M3_M2  M3_M2_10562
timestamp 1745462530
transform 1 0 412 0 1 2405
box -3 -3 3 3
use M3_M2  M3_M2_10563
timestamp 1745462530
transform 1 0 500 0 1 2005
box -3 -3 3 3
use M3_M2  M3_M2_10564
timestamp 1745462530
transform 1 0 436 0 1 2005
box -3 -3 3 3
use M3_M2  M3_M2_10565
timestamp 1745462530
transform 1 0 828 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_10566
timestamp 1745462530
transform 1 0 724 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_10567
timestamp 1745462530
transform 1 0 500 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_10568
timestamp 1745462530
transform 1 0 388 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_10569
timestamp 1745462530
transform 1 0 716 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_10570
timestamp 1745462530
transform 1 0 644 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_10571
timestamp 1745462530
transform 1 0 476 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_10572
timestamp 1745462530
transform 1 0 388 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_10573
timestamp 1745462530
transform 1 0 708 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_10574
timestamp 1745462530
transform 1 0 620 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_10575
timestamp 1745462530
transform 1 0 1172 0 1 165
box -3 -3 3 3
use M3_M2  M3_M2_10576
timestamp 1745462530
transform 1 0 1084 0 1 165
box -3 -3 3 3
use M3_M2  M3_M2_10577
timestamp 1745462530
transform 1 0 1532 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_10578
timestamp 1745462530
transform 1 0 1436 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_10579
timestamp 1745462530
transform 1 0 1460 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_10580
timestamp 1745462530
transform 1 0 1420 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_10581
timestamp 1745462530
transform 1 0 1428 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_10582
timestamp 1745462530
transform 1 0 1332 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_10583
timestamp 1745462530
transform 1 0 1596 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_10584
timestamp 1745462530
transform 1 0 1500 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_10585
timestamp 1745462530
transform 1 0 1660 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_10586
timestamp 1745462530
transform 1 0 1588 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_10587
timestamp 1745462530
transform 1 0 3188 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_10588
timestamp 1745462530
transform 1 0 3092 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_10589
timestamp 1745462530
transform 1 0 2748 0 1 335
box -3 -3 3 3
use M3_M2  M3_M2_10590
timestamp 1745462530
transform 1 0 2684 0 1 335
box -3 -3 3 3
use M3_M2  M3_M2_10591
timestamp 1745462530
transform 1 0 3108 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_10592
timestamp 1745462530
transform 1 0 3012 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_10593
timestamp 1745462530
transform 1 0 3060 0 1 335
box -3 -3 3 3
use M3_M2  M3_M2_10594
timestamp 1745462530
transform 1 0 2980 0 1 335
box -3 -3 3 3
use M3_M2  M3_M2_10595
timestamp 1745462530
transform 1 0 2940 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_10596
timestamp 1745462530
transform 1 0 2908 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_10597
timestamp 1745462530
transform 1 0 2916 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_10598
timestamp 1745462530
transform 1 0 2844 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_10599
timestamp 1745462530
transform 1 0 2948 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_10600
timestamp 1745462530
transform 1 0 2852 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_10601
timestamp 1745462530
transform 1 0 3268 0 1 335
box -3 -3 3 3
use M3_M2  M3_M2_10602
timestamp 1745462530
transform 1 0 3188 0 1 335
box -3 -3 3 3
use M3_M2  M3_M2_10603
timestamp 1745462530
transform 1 0 3364 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_10604
timestamp 1745462530
transform 1 0 3164 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_10605
timestamp 1745462530
transform 1 0 4140 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_10606
timestamp 1745462530
transform 1 0 4084 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_10607
timestamp 1745462530
transform 1 0 4228 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_10608
timestamp 1745462530
transform 1 0 4156 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_10609
timestamp 1745462530
transform 1 0 4068 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_10610
timestamp 1745462530
transform 1 0 4036 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_10611
timestamp 1745462530
transform 1 0 3396 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_10612
timestamp 1745462530
transform 1 0 3308 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_10613
timestamp 1745462530
transform 1 0 3380 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_10614
timestamp 1745462530
transform 1 0 3276 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_10615
timestamp 1745462530
transform 1 0 3540 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_10616
timestamp 1745462530
transform 1 0 3516 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_10617
timestamp 1745462530
transform 1 0 4140 0 1 1535
box -3 -3 3 3
use M3_M2  M3_M2_10618
timestamp 1745462530
transform 1 0 4084 0 1 1535
box -3 -3 3 3
use M3_M2  M3_M2_10619
timestamp 1745462530
transform 1 0 3572 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_10620
timestamp 1745462530
transform 1 0 3500 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_10621
timestamp 1745462530
transform 1 0 4252 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_10622
timestamp 1745462530
transform 1 0 4180 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_10623
timestamp 1745462530
transform 1 0 2828 0 1 1665
box -3 -3 3 3
use M3_M2  M3_M2_10624
timestamp 1745462530
transform 1 0 2780 0 1 1665
box -3 -3 3 3
use M3_M2  M3_M2_10625
timestamp 1745462530
transform 1 0 3276 0 1 2705
box -3 -3 3 3
use M3_M2  M3_M2_10626
timestamp 1745462530
transform 1 0 3212 0 1 2705
box -3 -3 3 3
use M3_M2  M3_M2_10627
timestamp 1745462530
transform 1 0 3004 0 1 2935
box -3 -3 3 3
use M3_M2  M3_M2_10628
timestamp 1745462530
transform 1 0 2932 0 1 2935
box -3 -3 3 3
use M3_M2  M3_M2_10629
timestamp 1745462530
transform 1 0 3260 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_10630
timestamp 1745462530
transform 1 0 3116 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_10631
timestamp 1745462530
transform 1 0 3204 0 1 3005
box -3 -3 3 3
use M3_M2  M3_M2_10632
timestamp 1745462530
transform 1 0 3132 0 1 3005
box -3 -3 3 3
use M3_M2  M3_M2_10633
timestamp 1745462530
transform 1 0 3260 0 1 2205
box -3 -3 3 3
use M3_M2  M3_M2_10634
timestamp 1745462530
transform 1 0 3196 0 1 2335
box -3 -3 3 3
use M3_M2  M3_M2_10635
timestamp 1745462530
transform 1 0 3196 0 1 2275
box -3 -3 3 3
use M3_M2  M3_M2_10636
timestamp 1745462530
transform 1 0 3180 0 1 2335
box -3 -3 3 3
use M3_M2  M3_M2_10637
timestamp 1745462530
transform 1 0 3148 0 1 2275
box -3 -3 3 3
use M3_M2  M3_M2_10638
timestamp 1745462530
transform 1 0 3148 0 1 2205
box -3 -3 3 3
use M3_M2  M3_M2_10639
timestamp 1745462530
transform 1 0 3180 0 1 2935
box -3 -3 3 3
use M3_M2  M3_M2_10640
timestamp 1745462530
transform 1 0 3108 0 1 2935
box -3 -3 3 3
use M3_M2  M3_M2_10641
timestamp 1745462530
transform 1 0 2780 0 1 2645
box -3 -3 3 3
use M3_M2  M3_M2_10642
timestamp 1745462530
transform 1 0 2732 0 1 2645
box -3 -3 3 3
use M3_M2  M3_M2_10643
timestamp 1745462530
transform 1 0 1748 0 1 2755
box -3 -3 3 3
use M3_M2  M3_M2_10644
timestamp 1745462530
transform 1 0 1692 0 1 2755
box -3 -3 3 3
use M3_M2  M3_M2_10645
timestamp 1745462530
transform 1 0 1700 0 1 1975
box -3 -3 3 3
use M3_M2  M3_M2_10646
timestamp 1745462530
transform 1 0 1612 0 1 1975
box -3 -3 3 3
use M3_M2  M3_M2_10647
timestamp 1745462530
transform 1 0 1644 0 1 2535
box -3 -3 3 3
use M3_M2  M3_M2_10648
timestamp 1745462530
transform 1 0 1540 0 1 2535
box -3 -3 3 3
use M3_M2  M3_M2_10649
timestamp 1745462530
transform 1 0 436 0 1 2745
box -3 -3 3 3
use M3_M2  M3_M2_10650
timestamp 1745462530
transform 1 0 356 0 1 2745
box -3 -3 3 3
use M3_M2  M3_M2_10651
timestamp 1745462530
transform 1 0 524 0 1 2635
box -3 -3 3 3
use M3_M2  M3_M2_10652
timestamp 1745462530
transform 1 0 452 0 1 2635
box -3 -3 3 3
use M3_M2  M3_M2_10653
timestamp 1745462530
transform 1 0 348 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_10654
timestamp 1745462530
transform 1 0 260 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_10655
timestamp 1745462530
transform 1 0 1068 0 1 2555
box -3 -3 3 3
use M3_M2  M3_M2_10656
timestamp 1745462530
transform 1 0 964 0 1 2555
box -3 -3 3 3
use M3_M2  M3_M2_10657
timestamp 1745462530
transform 1 0 452 0 1 2335
box -3 -3 3 3
use M3_M2  M3_M2_10658
timestamp 1745462530
transform 1 0 372 0 1 2335
box -3 -3 3 3
use M3_M2  M3_M2_10659
timestamp 1745462530
transform 1 0 380 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_10660
timestamp 1745462530
transform 1 0 316 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_10661
timestamp 1745462530
transform 1 0 548 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_10662
timestamp 1745462530
transform 1 0 476 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_10663
timestamp 1745462530
transform 1 0 772 0 1 1435
box -3 -3 3 3
use M3_M2  M3_M2_10664
timestamp 1745462530
transform 1 0 708 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_10665
timestamp 1745462530
transform 1 0 1844 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_10666
timestamp 1745462530
transform 1 0 1828 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_10667
timestamp 1745462530
transform 1 0 1852 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_10668
timestamp 1745462530
transform 1 0 1836 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_10669
timestamp 1745462530
transform 1 0 2004 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_10670
timestamp 1745462530
transform 1 0 1908 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_10671
timestamp 1745462530
transform 1 0 2036 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_10672
timestamp 1745462530
transform 1 0 1948 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_10673
timestamp 1745462530
transform 1 0 2004 0 1 1215
box -3 -3 3 3
use M3_M2  M3_M2_10674
timestamp 1745462530
transform 1 0 1940 0 1 1215
box -3 -3 3 3
use M3_M2  M3_M2_10675
timestamp 1745462530
transform 1 0 1940 0 1 1335
box -3 -3 3 3
use M3_M2  M3_M2_10676
timestamp 1745462530
transform 1 0 1916 0 1 1335
box -3 -3 3 3
use M3_M2  M3_M2_10677
timestamp 1745462530
transform 1 0 2244 0 1 255
box -3 -3 3 3
use M3_M2  M3_M2_10678
timestamp 1745462530
transform 1 0 2132 0 1 255
box -3 -3 3 3
use M3_M2  M3_M2_10679
timestamp 1745462530
transform 1 0 2204 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_10680
timestamp 1745462530
transform 1 0 2116 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_10681
timestamp 1745462530
transform 1 0 2244 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_10682
timestamp 1745462530
transform 1 0 2148 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_10683
timestamp 1745462530
transform 1 0 2508 0 1 125
box -3 -3 3 3
use M3_M2  M3_M2_10684
timestamp 1745462530
transform 1 0 2404 0 1 115
box -3 -3 3 3
use M3_M2  M3_M2_10685
timestamp 1745462530
transform 1 0 2356 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_10686
timestamp 1745462530
transform 1 0 2220 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_10687
timestamp 1745462530
transform 1 0 2308 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_10688
timestamp 1745462530
transform 1 0 2236 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_10689
timestamp 1745462530
transform 1 0 2372 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_10690
timestamp 1745462530
transform 1 0 2268 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_10691
timestamp 1745462530
transform 1 0 4300 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_10692
timestamp 1745462530
transform 1 0 4228 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_10693
timestamp 1745462530
transform 1 0 4076 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_10694
timestamp 1745462530
transform 1 0 3996 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_10695
timestamp 1745462530
transform 1 0 4316 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_10696
timestamp 1745462530
transform 1 0 4252 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_10697
timestamp 1745462530
transform 1 0 4316 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_10698
timestamp 1745462530
transform 1 0 4228 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_10699
timestamp 1745462530
transform 1 0 4028 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_10700
timestamp 1745462530
transform 1 0 3932 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_10701
timestamp 1745462530
transform 1 0 4308 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_10702
timestamp 1745462530
transform 1 0 4220 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_10703
timestamp 1745462530
transform 1 0 4316 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_10704
timestamp 1745462530
transform 1 0 4228 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_10705
timestamp 1745462530
transform 1 0 3668 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_10706
timestamp 1745462530
transform 1 0 3636 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_10707
timestamp 1745462530
transform 1 0 4324 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_10708
timestamp 1745462530
transform 1 0 4300 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_10709
timestamp 1745462530
transform 1 0 3308 0 1 1855
box -3 -3 3 3
use M3_M2  M3_M2_10710
timestamp 1745462530
transform 1 0 3284 0 1 1855
box -3 -3 3 3
use M3_M2  M3_M2_10711
timestamp 1745462530
transform 1 0 2676 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_10712
timestamp 1745462530
transform 1 0 2596 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_10713
timestamp 1745462530
transform 1 0 4276 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_10714
timestamp 1745462530
transform 1 0 4204 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_10715
timestamp 1745462530
transform 1 0 3988 0 1 2915
box -3 -3 3 3
use M3_M2  M3_M2_10716
timestamp 1745462530
transform 1 0 3908 0 1 2915
box -3 -3 3 3
use M3_M2  M3_M2_10717
timestamp 1745462530
transform 1 0 4316 0 1 2805
box -3 -3 3 3
use M3_M2  M3_M2_10718
timestamp 1745462530
transform 1 0 4164 0 1 2805
box -3 -3 3 3
use M3_M2  M3_M2_10719
timestamp 1745462530
transform 1 0 4316 0 1 2915
box -3 -3 3 3
use M3_M2  M3_M2_10720
timestamp 1745462530
transform 1 0 4236 0 1 2915
box -3 -3 3 3
use M3_M2  M3_M2_10721
timestamp 1745462530
transform 1 0 4300 0 1 2425
box -3 -3 3 3
use M3_M2  M3_M2_10722
timestamp 1745462530
transform 1 0 4228 0 1 2425
box -3 -3 3 3
use M3_M2  M3_M2_10723
timestamp 1745462530
transform 1 0 4140 0 1 2915
box -3 -3 3 3
use M3_M2  M3_M2_10724
timestamp 1745462530
transform 1 0 4068 0 1 2915
box -3 -3 3 3
use M3_M2  M3_M2_10725
timestamp 1745462530
transform 1 0 2620 0 1 2905
box -3 -3 3 3
use M3_M2  M3_M2_10726
timestamp 1745462530
transform 1 0 2556 0 1 2905
box -3 -3 3 3
use M3_M2  M3_M2_10727
timestamp 1745462530
transform 1 0 1876 0 1 2675
box -3 -3 3 3
use M3_M2  M3_M2_10728
timestamp 1745462530
transform 1 0 1836 0 1 2675
box -3 -3 3 3
use M3_M2  M3_M2_10729
timestamp 1745462530
transform 1 0 2012 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_10730
timestamp 1745462530
transform 1 0 1844 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_10731
timestamp 1745462530
transform 1 0 1908 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_10732
timestamp 1745462530
transform 1 0 1812 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_10733
timestamp 1745462530
transform 1 0 1036 0 1 2915
box -3 -3 3 3
use M3_M2  M3_M2_10734
timestamp 1745462530
transform 1 0 916 0 1 2915
box -3 -3 3 3
use M3_M2  M3_M2_10735
timestamp 1745462530
transform 1 0 380 0 1 2165
box -3 -3 3 3
use M3_M2  M3_M2_10736
timestamp 1745462530
transform 1 0 332 0 1 2175
box -3 -3 3 3
use M3_M2  M3_M2_10737
timestamp 1745462530
transform 1 0 364 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_10738
timestamp 1745462530
transform 1 0 300 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_10739
timestamp 1745462530
transform 1 0 788 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_10740
timestamp 1745462530
transform 1 0 668 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_10741
timestamp 1745462530
transform 1 0 364 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_10742
timestamp 1745462530
transform 1 0 260 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_10743
timestamp 1745462530
transform 1 0 212 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_10744
timestamp 1745462530
transform 1 0 140 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_10745
timestamp 1745462530
transform 1 0 212 0 1 245
box -3 -3 3 3
use M3_M2  M3_M2_10746
timestamp 1745462530
transform 1 0 148 0 1 245
box -3 -3 3 3
use M3_M2  M3_M2_10747
timestamp 1745462530
transform 1 0 212 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_10748
timestamp 1745462530
transform 1 0 148 0 1 405
box -3 -3 3 3
use M3_M2  M3_M2_10749
timestamp 1745462530
transform 1 0 812 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_10750
timestamp 1745462530
transform 1 0 724 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_10751
timestamp 1745462530
transform 1 0 204 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_10752
timestamp 1745462530
transform 1 0 164 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_10753
timestamp 1745462530
transform 1 0 2020 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_10754
timestamp 1745462530
transform 1 0 1932 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_10755
timestamp 1745462530
transform 1 0 2004 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_10756
timestamp 1745462530
transform 1 0 1900 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_10757
timestamp 1745462530
transform 1 0 2020 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_10758
timestamp 1745462530
transform 1 0 1900 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_10759
timestamp 1745462530
transform 1 0 2012 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_10760
timestamp 1745462530
transform 1 0 1908 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_10761
timestamp 1745462530
transform 1 0 2084 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_10762
timestamp 1745462530
transform 1 0 2012 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_10763
timestamp 1745462530
transform 1 0 2180 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_10764
timestamp 1745462530
transform 1 0 2012 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_10765
timestamp 1745462530
transform 1 0 2116 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_10766
timestamp 1745462530
transform 1 0 2004 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_10767
timestamp 1745462530
transform 1 0 2356 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_10768
timestamp 1745462530
transform 1 0 2292 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_10769
timestamp 1745462530
transform 1 0 2380 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_10770
timestamp 1745462530
transform 1 0 2308 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_10771
timestamp 1745462530
transform 1 0 2292 0 1 875
box -3 -3 3 3
use M3_M2  M3_M2_10772
timestamp 1745462530
transform 1 0 2204 0 1 875
box -3 -3 3 3
use M3_M2  M3_M2_10773
timestamp 1745462530
transform 1 0 3460 0 1 335
box -3 -3 3 3
use M3_M2  M3_M2_10774
timestamp 1745462530
transform 1 0 3396 0 1 335
box -3 -3 3 3
use M3_M2  M3_M2_10775
timestamp 1745462530
transform 1 0 4308 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_10776
timestamp 1745462530
transform 1 0 4228 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_10777
timestamp 1745462530
transform 1 0 3868 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_10778
timestamp 1745462530
transform 1 0 3788 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_10779
timestamp 1745462530
transform 1 0 4316 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_10780
timestamp 1745462530
transform 1 0 4228 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_10781
timestamp 1745462530
transform 1 0 3788 0 1 1135
box -3 -3 3 3
use M3_M2  M3_M2_10782
timestamp 1745462530
transform 1 0 3748 0 1 1135
box -3 -3 3 3
use M3_M2  M3_M2_10783
timestamp 1745462530
transform 1 0 4308 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_10784
timestamp 1745462530
transform 1 0 4220 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_10785
timestamp 1745462530
transform 1 0 3900 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_10786
timestamp 1745462530
transform 1 0 3820 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_10787
timestamp 1745462530
transform 1 0 3972 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_10788
timestamp 1745462530
transform 1 0 3884 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_10789
timestamp 1745462530
transform 1 0 3084 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_10790
timestamp 1745462530
transform 1 0 2980 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_10791
timestamp 1745462530
transform 1 0 2708 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_10792
timestamp 1745462530
transform 1 0 2588 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_10793
timestamp 1745462530
transform 1 0 3772 0 1 3015
box -3 -3 3 3
use M3_M2  M3_M2_10794
timestamp 1745462530
transform 1 0 3684 0 1 3015
box -3 -3 3 3
use M3_M2  M3_M2_10795
timestamp 1745462530
transform 1 0 3932 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_10796
timestamp 1745462530
transform 1 0 3868 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_10797
timestamp 1745462530
transform 1 0 3820 0 1 2945
box -3 -3 3 3
use M3_M2  M3_M2_10798
timestamp 1745462530
transform 1 0 3740 0 1 2945
box -3 -3 3 3
use M3_M2  M3_M2_10799
timestamp 1745462530
transform 1 0 3916 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_10800
timestamp 1745462530
transform 1 0 3844 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_10801
timestamp 1745462530
transform 1 0 4004 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_10802
timestamp 1745462530
transform 1 0 3940 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_10803
timestamp 1745462530
transform 1 0 3092 0 1 2405
box -3 -3 3 3
use M3_M2  M3_M2_10804
timestamp 1745462530
transform 1 0 2988 0 1 2405
box -3 -3 3 3
use M3_M2  M3_M2_10805
timestamp 1745462530
transform 1 0 2508 0 1 2845
box -3 -3 3 3
use M3_M2  M3_M2_10806
timestamp 1745462530
transform 1 0 2444 0 1 2845
box -3 -3 3 3
use M3_M2  M3_M2_10807
timestamp 1745462530
transform 1 0 1244 0 1 2945
box -3 -3 3 3
use M3_M2  M3_M2_10808
timestamp 1745462530
transform 1 0 1100 0 1 2945
box -3 -3 3 3
use M3_M2  M3_M2_10809
timestamp 1745462530
transform 1 0 1228 0 1 2205
box -3 -3 3 3
use M3_M2  M3_M2_10810
timestamp 1745462530
transform 1 0 1060 0 1 2205
box -3 -3 3 3
use M3_M2  M3_M2_10811
timestamp 1745462530
transform 1 0 1236 0 1 2765
box -3 -3 3 3
use M3_M2  M3_M2_10812
timestamp 1745462530
transform 1 0 1140 0 1 2765
box -3 -3 3 3
use M3_M2  M3_M2_10813
timestamp 1745462530
transform 1 0 1212 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_10814
timestamp 1745462530
transform 1 0 1020 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_10815
timestamp 1745462530
transform 1 0 1188 0 1 2535
box -3 -3 3 3
use M3_M2  M3_M2_10816
timestamp 1745462530
transform 1 0 1100 0 1 2535
box -3 -3 3 3
use M3_M2  M3_M2_10817
timestamp 1745462530
transform 1 0 1172 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_10818
timestamp 1745462530
transform 1 0 1156 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_10819
timestamp 1745462530
transform 1 0 836 0 1 2535
box -3 -3 3 3
use M3_M2  M3_M2_10820
timestamp 1745462530
transform 1 0 796 0 1 2535
box -3 -3 3 3
use M3_M2  M3_M2_10821
timestamp 1745462530
transform 1 0 228 0 1 2715
box -3 -3 3 3
use M3_M2  M3_M2_10822
timestamp 1745462530
transform 1 0 124 0 1 2715
box -3 -3 3 3
use M3_M2  M3_M2_10823
timestamp 1745462530
transform 1 0 204 0 1 2355
box -3 -3 3 3
use M3_M2  M3_M2_10824
timestamp 1745462530
transform 1 0 140 0 1 2355
box -3 -3 3 3
use M3_M2  M3_M2_10825
timestamp 1745462530
transform 1 0 220 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_10826
timestamp 1745462530
transform 1 0 140 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_10827
timestamp 1745462530
transform 1 0 220 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_10828
timestamp 1745462530
transform 1 0 140 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_10829
timestamp 1745462530
transform 1 0 820 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_10830
timestamp 1745462530
transform 1 0 692 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_10831
timestamp 1745462530
transform 1 0 228 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_10832
timestamp 1745462530
transform 1 0 132 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_10833
timestamp 1745462530
transform 1 0 212 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_10834
timestamp 1745462530
transform 1 0 116 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_10835
timestamp 1745462530
transform 1 0 244 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_10836
timestamp 1745462530
transform 1 0 148 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_10837
timestamp 1745462530
transform 1 0 212 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_10838
timestamp 1745462530
transform 1 0 140 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_10839
timestamp 1745462530
transform 1 0 220 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_10840
timestamp 1745462530
transform 1 0 124 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_10841
timestamp 1745462530
transform 1 0 1044 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_10842
timestamp 1745462530
transform 1 0 956 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_10843
timestamp 1745462530
transform 1 0 1132 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_10844
timestamp 1745462530
transform 1 0 1028 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_10845
timestamp 1745462530
transform 1 0 1164 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_10846
timestamp 1745462530
transform 1 0 1060 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_10847
timestamp 1745462530
transform 1 0 1332 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_10848
timestamp 1745462530
transform 1 0 1244 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_10849
timestamp 1745462530
transform 1 0 1356 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_10850
timestamp 1745462530
transform 1 0 1220 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_10851
timestamp 1745462530
transform 1 0 1420 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_10852
timestamp 1745462530
transform 1 0 1292 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_10853
timestamp 1745462530
transform 1 0 1420 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_10854
timestamp 1745462530
transform 1 0 1332 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_10855
timestamp 1745462530
transform 1 0 1476 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_10856
timestamp 1745462530
transform 1 0 1348 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_10857
timestamp 1745462530
transform 1 0 1532 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_10858
timestamp 1745462530
transform 1 0 1452 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_10859
timestamp 1745462530
transform 1 0 2308 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_10860
timestamp 1745462530
transform 1 0 2148 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_10861
timestamp 1745462530
transform 1 0 2204 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_10862
timestamp 1745462530
transform 1 0 2124 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_10863
timestamp 1745462530
transform 1 0 2308 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_10864
timestamp 1745462530
transform 1 0 2140 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_10865
timestamp 1745462530
transform 1 0 2300 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_10866
timestamp 1745462530
transform 1 0 2156 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_10867
timestamp 1745462530
transform 1 0 2628 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_10868
timestamp 1745462530
transform 1 0 2564 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_10869
timestamp 1745462530
transform 1 0 3532 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_10870
timestamp 1745462530
transform 1 0 3460 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_10871
timestamp 1745462530
transform 1 0 4100 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_10872
timestamp 1745462530
transform 1 0 4004 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_10873
timestamp 1745462530
transform 1 0 3964 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_10874
timestamp 1745462530
transform 1 0 3908 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_10875
timestamp 1745462530
transform 1 0 3500 0 1 1275
box -3 -3 3 3
use M3_M2  M3_M2_10876
timestamp 1745462530
transform 1 0 3460 0 1 1275
box -3 -3 3 3
use M3_M2  M3_M2_10877
timestamp 1745462530
transform 1 0 4092 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_10878
timestamp 1745462530
transform 1 0 3972 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_10879
timestamp 1745462530
transform 1 0 3484 0 1 1855
box -3 -3 3 3
use M3_M2  M3_M2_10880
timestamp 1745462530
transform 1 0 3412 0 1 1855
box -3 -3 3 3
use M3_M2  M3_M2_10881
timestamp 1745462530
transform 1 0 3460 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_10882
timestamp 1745462530
transform 1 0 3396 0 1 2205
box -3 -3 3 3
use M3_M2  M3_M2_10883
timestamp 1745462530
transform 1 0 2796 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_10884
timestamp 1745462530
transform 1 0 2724 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_10885
timestamp 1745462530
transform 1 0 2636 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_10886
timestamp 1745462530
transform 1 0 2540 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_10887
timestamp 1745462530
transform 1 0 3484 0 1 2775
box -3 -3 3 3
use M3_M2  M3_M2_10888
timestamp 1745462530
transform 1 0 3452 0 1 2775
box -3 -3 3 3
use M3_M2  M3_M2_10889
timestamp 1745462530
transform 1 0 3388 0 1 2985
box -3 -3 3 3
use M3_M2  M3_M2_10890
timestamp 1745462530
transform 1 0 3300 0 1 2985
box -3 -3 3 3
use M3_M2  M3_M2_10891
timestamp 1745462530
transform 1 0 3468 0 1 2455
box -3 -3 3 3
use M3_M2  M3_M2_10892
timestamp 1745462530
transform 1 0 3436 0 1 2455
box -3 -3 3 3
use M3_M2  M3_M2_10893
timestamp 1745462530
transform 1 0 3436 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_10894
timestamp 1745462530
transform 1 0 3380 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_10895
timestamp 1745462530
transform 1 0 3204 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_10896
timestamp 1745462530
transform 1 0 2892 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_10897
timestamp 1745462530
transform 1 0 1436 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_10898
timestamp 1745462530
transform 1 0 1420 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_10899
timestamp 1745462530
transform 1 0 1396 0 1 2535
box -3 -3 3 3
use M3_M2  M3_M2_10900
timestamp 1745462530
transform 1 0 1340 0 1 2535
box -3 -3 3 3
use M3_M2  M3_M2_10901
timestamp 1745462530
transform 1 0 276 0 1 2745
box -3 -3 3 3
use M3_M2  M3_M2_10902
timestamp 1745462530
transform 1 0 124 0 1 2745
box -3 -3 3 3
use M3_M2  M3_M2_10903
timestamp 1745462530
transform 1 0 588 0 1 2745
box -3 -3 3 3
use M3_M2  M3_M2_10904
timestamp 1745462530
transform 1 0 524 0 1 2745
box -3 -3 3 3
use M3_M2  M3_M2_10905
timestamp 1745462530
transform 1 0 228 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_10906
timestamp 1745462530
transform 1 0 140 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_10907
timestamp 1745462530
transform 1 0 1004 0 1 2755
box -3 -3 3 3
use M3_M2  M3_M2_10908
timestamp 1745462530
transform 1 0 948 0 1 2755
box -3 -3 3 3
use M3_M2  M3_M2_10909
timestamp 1745462530
transform 1 0 220 0 1 2425
box -3 -3 3 3
use M3_M2  M3_M2_10910
timestamp 1745462530
transform 1 0 140 0 1 2425
box -3 -3 3 3
use M3_M2  M3_M2_10911
timestamp 1745462530
transform 1 0 204 0 1 2005
box -3 -3 3 3
use M3_M2  M3_M2_10912
timestamp 1745462530
transform 1 0 108 0 1 2005
box -3 -3 3 3
use M3_M2  M3_M2_10913
timestamp 1745462530
transform 1 0 180 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_10914
timestamp 1745462530
transform 1 0 140 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_10915
timestamp 1745462530
transform 1 0 300 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_10916
timestamp 1745462530
transform 1 0 132 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_10917
timestamp 1745462530
transform 1 0 380 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_10918
timestamp 1745462530
transform 1 0 308 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_10919
timestamp 1745462530
transform 1 0 484 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_10920
timestamp 1745462530
transform 1 0 404 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_10921
timestamp 1745462530
transform 1 0 540 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_10922
timestamp 1745462530
transform 1 0 492 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_10923
timestamp 1745462530
transform 1 0 828 0 1 245
box -3 -3 3 3
use M3_M2  M3_M2_10924
timestamp 1745462530
transform 1 0 764 0 1 245
box -3 -3 3 3
use M3_M2  M3_M2_10925
timestamp 1745462530
transform 1 0 868 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_10926
timestamp 1745462530
transform 1 0 788 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_10927
timestamp 1745462530
transform 1 0 1108 0 1 205
box -3 -3 3 3
use M3_M2  M3_M2_10928
timestamp 1745462530
transform 1 0 1028 0 1 205
box -3 -3 3 3
use M3_M2  M3_M2_10929
timestamp 1745462530
transform 1 0 1036 0 1 575
box -3 -3 3 3
use M3_M2  M3_M2_10930
timestamp 1745462530
transform 1 0 1004 0 1 575
box -3 -3 3 3
use M3_M2  M3_M2_10931
timestamp 1745462530
transform 1 0 1372 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_10932
timestamp 1745462530
transform 1 0 1300 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_10933
timestamp 1745462530
transform 1 0 1268 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_10934
timestamp 1745462530
transform 1 0 1156 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_10935
timestamp 1745462530
transform 1 0 1324 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_10936
timestamp 1745462530
transform 1 0 1220 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_10937
timestamp 1745462530
transform 1 0 1428 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_10938
timestamp 1745462530
transform 1 0 1332 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_10939
timestamp 1745462530
transform 1 0 1420 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_10940
timestamp 1745462530
transform 1 0 1340 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_10941
timestamp 1745462530
transform 1 0 2852 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_10942
timestamp 1745462530
transform 1 0 2756 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_10943
timestamp 1745462530
transform 1 0 2692 0 1 1485
box -3 -3 3 3
use M3_M2  M3_M2_10944
timestamp 1745462530
transform 1 0 2660 0 1 1485
box -3 -3 3 3
use M3_M2  M3_M2_10945
timestamp 1745462530
transform 1 0 4308 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_10946
timestamp 1745462530
transform 1 0 4236 0 1 815
box -3 -3 3 3
use M3_M2  M3_M2_10947
timestamp 1745462530
transform 1 0 4308 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_10948
timestamp 1745462530
transform 1 0 4228 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_10949
timestamp 1745462530
transform 1 0 3684 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_10950
timestamp 1745462530
transform 1 0 3596 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_10951
timestamp 1745462530
transform 1 0 4316 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_10952
timestamp 1745462530
transform 1 0 4228 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_10953
timestamp 1745462530
transform 1 0 3788 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_10954
timestamp 1745462530
transform 1 0 3748 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_10955
timestamp 1745462530
transform 1 0 3668 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_10956
timestamp 1745462530
transform 1 0 3588 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_10957
timestamp 1745462530
transform 1 0 3708 0 1 2985
box -3 -3 3 3
use M3_M2  M3_M2_10958
timestamp 1745462530
transform 1 0 3620 0 1 2985
box -3 -3 3 3
use M3_M2  M3_M2_10959
timestamp 1745462530
transform 1 0 3708 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_10960
timestamp 1745462530
transform 1 0 3636 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_10961
timestamp 1745462530
transform 1 0 3628 0 1 2945
box -3 -3 3 3
use M3_M2  M3_M2_10962
timestamp 1745462530
transform 1 0 3540 0 1 2945
box -3 -3 3 3
use M3_M2  M3_M2_10963
timestamp 1745462530
transform 1 0 3740 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_10964
timestamp 1745462530
transform 1 0 3668 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_10965
timestamp 1745462530
transform 1 0 3700 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_10966
timestamp 1745462530
transform 1 0 3628 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_10967
timestamp 1745462530
transform 1 0 2988 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_10968
timestamp 1745462530
transform 1 0 2876 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_10969
timestamp 1745462530
transform 1 0 2636 0 1 2755
box -3 -3 3 3
use M3_M2  M3_M2_10970
timestamp 1745462530
transform 1 0 2572 0 1 2755
box -3 -3 3 3
use M3_M2  M3_M2_10971
timestamp 1745462530
transform 1 0 2404 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_10972
timestamp 1745462530
transform 1 0 2340 0 1 2815
box -3 -3 3 3
use M3_M2  M3_M2_10973
timestamp 1745462530
transform 1 0 2308 0 1 2915
box -3 -3 3 3
use M3_M2  M3_M2_10974
timestamp 1745462530
transform 1 0 2244 0 1 2915
box -3 -3 3 3
use M3_M2  M3_M2_10975
timestamp 1745462530
transform 1 0 2228 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_10976
timestamp 1745462530
transform 1 0 2172 0 1 2815
box -3 -3 3 3
use M3_M2  M3_M2_10977
timestamp 1745462530
transform 1 0 2076 0 1 2775
box -3 -3 3 3
use M3_M2  M3_M2_10978
timestamp 1745462530
transform 1 0 2028 0 1 2775
box -3 -3 3 3
use M3_M2  M3_M2_10979
timestamp 1745462530
transform 1 0 2284 0 1 3045
box -3 -3 3 3
use M3_M2  M3_M2_10980
timestamp 1745462530
transform 1 0 2260 0 1 3045
box -3 -3 3 3
use M3_M2  M3_M2_10981
timestamp 1745462530
transform 1 0 1324 0 1 3155
box -3 -3 3 3
use M3_M2  M3_M2_10982
timestamp 1745462530
transform 1 0 1228 0 1 3155
box -3 -3 3 3
use M3_M2  M3_M2_10983
timestamp 1745462530
transform 1 0 1132 0 1 4145
box -3 -3 3 3
use M3_M2  M3_M2_10984
timestamp 1745462530
transform 1 0 1068 0 1 4145
box -3 -3 3 3
use M3_M2  M3_M2_10985
timestamp 1745462530
transform 1 0 1004 0 1 4145
box -3 -3 3 3
use M3_M2  M3_M2_10986
timestamp 1745462530
transform 1 0 1116 0 1 4195
box -3 -3 3 3
use M3_M2  M3_M2_10987
timestamp 1745462530
transform 1 0 1020 0 1 4195
box -3 -3 3 3
use M3_M2  M3_M2_10988
timestamp 1745462530
transform 1 0 908 0 1 4195
box -3 -3 3 3
use M3_M2  M3_M2_10989
timestamp 1745462530
transform 1 0 4036 0 1 4125
box -3 -3 3 3
use M3_M2  M3_M2_10990
timestamp 1745462530
transform 1 0 4028 0 1 4225
box -3 -3 3 3
use M3_M2  M3_M2_10991
timestamp 1745462530
transform 1 0 3996 0 1 4225
box -3 -3 3 3
use M3_M2  M3_M2_10992
timestamp 1745462530
transform 1 0 3996 0 1 4175
box -3 -3 3 3
use M3_M2  M3_M2_10993
timestamp 1745462530
transform 1 0 3996 0 1 4125
box -3 -3 3 3
use M3_M2  M3_M2_10994
timestamp 1745462530
transform 1 0 2964 0 1 4175
box -3 -3 3 3
use M3_M2  M3_M2_10995
timestamp 1745462530
transform 1 0 2596 0 1 4175
box -3 -3 3 3
use M3_M2  M3_M2_10996
timestamp 1745462530
transform 1 0 2068 0 1 4235
box -3 -3 3 3
use M3_M2  M3_M2_10997
timestamp 1745462530
transform 1 0 2068 0 1 4175
box -3 -3 3 3
use M3_M2  M3_M2_10998
timestamp 1745462530
transform 1 0 2020 0 1 4235
box -3 -3 3 3
use M3_M2  M3_M2_10999
timestamp 1745462530
transform 1 0 1852 0 1 4235
box -3 -3 3 3
use M3_M2  M3_M2_11000
timestamp 1745462530
transform 1 0 1692 0 1 4235
box -3 -3 3 3
use M3_M2  M3_M2_11001
timestamp 1745462530
transform 1 0 1692 0 1 4045
box -3 -3 3 3
use M3_M2  M3_M2_11002
timestamp 1745462530
transform 1 0 1300 0 1 4035
box -3 -3 3 3
use M3_M2  M3_M2_11003
timestamp 1745462530
transform 1 0 1212 0 1 4035
box -3 -3 3 3
use M3_M2  M3_M2_11004
timestamp 1745462530
transform 1 0 1092 0 1 4035
box -3 -3 3 3
use M3_M2  M3_M2_11005
timestamp 1745462530
transform 1 0 1036 0 1 4035
box -3 -3 3 3
use M3_M2  M3_M2_11006
timestamp 1745462530
transform 1 0 948 0 1 4095
box -3 -3 3 3
use M3_M2  M3_M2_11007
timestamp 1745462530
transform 1 0 948 0 1 4035
box -3 -3 3 3
use M3_M2  M3_M2_11008
timestamp 1745462530
transform 1 0 868 0 1 4095
box -3 -3 3 3
use M3_M2  M3_M2_11009
timestamp 1745462530
transform 1 0 716 0 1 4205
box -3 -3 3 3
use M3_M2  M3_M2_11010
timestamp 1745462530
transform 1 0 628 0 1 4205
box -3 -3 3 3
use M3_M2  M3_M2_11011
timestamp 1745462530
transform 1 0 572 0 1 4215
box -3 -3 3 3
use M3_M2  M3_M2_11012
timestamp 1745462530
transform 1 0 844 0 1 3945
box -3 -3 3 3
use M3_M2  M3_M2_11013
timestamp 1745462530
transform 1 0 788 0 1 3945
box -3 -3 3 3
use M3_M2  M3_M2_11014
timestamp 1745462530
transform 1 0 732 0 1 3945
box -3 -3 3 3
use M3_M2  M3_M2_11015
timestamp 1745462530
transform 1 0 468 0 1 3945
box -3 -3 3 3
use M3_M2  M3_M2_11016
timestamp 1745462530
transform 1 0 772 0 1 3995
box -3 -3 3 3
use M3_M2  M3_M2_11017
timestamp 1745462530
transform 1 0 492 0 1 3995
box -3 -3 3 3
use M3_M2  M3_M2_11018
timestamp 1745462530
transform 1 0 1140 0 1 4205
box -3 -3 3 3
use M3_M2  M3_M2_11019
timestamp 1745462530
transform 1 0 1068 0 1 4205
box -3 -3 3 3
use M3_M2  M3_M2_11020
timestamp 1745462530
transform 1 0 1748 0 1 4195
box -3 -3 3 3
use M3_M2  M3_M2_11021
timestamp 1745462530
transform 1 0 1676 0 1 4195
box -3 -3 3 3
use M3_M2  M3_M2_11022
timestamp 1745462530
transform 1 0 4316 0 1 4025
box -3 -3 3 3
use M3_M2  M3_M2_11023
timestamp 1745462530
transform 1 0 4268 0 1 4025
box -3 -3 3 3
use M3_M2  M3_M2_11024
timestamp 1745462530
transform 1 0 4308 0 1 4205
box -3 -3 3 3
use M3_M2  M3_M2_11025
timestamp 1745462530
transform 1 0 4268 0 1 4205
box -3 -3 3 3
use M3_M2  M3_M2_11026
timestamp 1745462530
transform 1 0 1492 0 1 4225
box -3 -3 3 3
use M3_M2  M3_M2_11027
timestamp 1745462530
transform 1 0 1444 0 1 4225
box -3 -3 3 3
use M3_M2  M3_M2_11028
timestamp 1745462530
transform 1 0 780 0 1 4165
box -3 -3 3 3
use M3_M2  M3_M2_11029
timestamp 1745462530
transform 1 0 636 0 1 4165
box -3 -3 3 3
use M3_M2  M3_M2_11030
timestamp 1745462530
transform 1 0 740 0 1 4125
box -3 -3 3 3
use M3_M2  M3_M2_11031
timestamp 1745462530
transform 1 0 700 0 1 4125
box -3 -3 3 3
use M3_M2  M3_M2_11032
timestamp 1745462530
transform 1 0 676 0 1 4125
box -3 -3 3 3
use M3_M2  M3_M2_11033
timestamp 1745462530
transform 1 0 684 0 1 4225
box -3 -3 3 3
use M3_M2  M3_M2_11034
timestamp 1745462530
transform 1 0 612 0 1 4225
box -3 -3 3 3
use M3_M2  M3_M2_11035
timestamp 1745462530
transform 1 0 900 0 1 4015
box -3 -3 3 3
use M3_M2  M3_M2_11036
timestamp 1745462530
transform 1 0 868 0 1 4015
box -3 -3 3 3
use M3_M2  M3_M2_11037
timestamp 1745462530
transform 1 0 836 0 1 4015
box -3 -3 3 3
use M3_M2  M3_M2_11038
timestamp 1745462530
transform 1 0 716 0 1 4015
box -3 -3 3 3
use M3_M2  M3_M2_11039
timestamp 1745462530
transform 1 0 668 0 1 4015
box -3 -3 3 3
use M3_M2  M3_M2_11040
timestamp 1745462530
transform 1 0 4212 0 1 4095
box -3 -3 3 3
use M3_M2  M3_M2_11041
timestamp 1745462530
transform 1 0 4124 0 1 4185
box -3 -3 3 3
use M3_M2  M3_M2_11042
timestamp 1745462530
transform 1 0 4124 0 1 4095
box -3 -3 3 3
use M3_M2  M3_M2_11043
timestamp 1745462530
transform 1 0 2868 0 1 4305
box -3 -3 3 3
use M3_M2  M3_M2_11044
timestamp 1745462530
transform 1 0 2868 0 1 4205
box -3 -3 3 3
use M3_M2  M3_M2_11045
timestamp 1745462530
transform 1 0 2276 0 1 4295
box -3 -3 3 3
use M3_M2  M3_M2_11046
timestamp 1745462530
transform 1 0 2276 0 1 4165
box -3 -3 3 3
use M3_M2  M3_M2_11047
timestamp 1745462530
transform 1 0 2164 0 1 4165
box -3 -3 3 3
use M3_M2  M3_M2_11048
timestamp 1745462530
transform 1 0 2148 0 1 4125
box -3 -3 3 3
use M3_M2  M3_M2_11049
timestamp 1745462530
transform 1 0 1716 0 1 4135
box -3 -3 3 3
use M3_M2  M3_M2_11050
timestamp 1745462530
transform 1 0 1556 0 1 4145
box -3 -3 3 3
use M3_M2  M3_M2_11051
timestamp 1745462530
transform 1 0 1508 0 1 4145
box -3 -3 3 3
use M3_M2  M3_M2_11052
timestamp 1745462530
transform 1 0 1500 0 1 4075
box -3 -3 3 3
use M3_M2  M3_M2_11053
timestamp 1745462530
transform 1 0 1436 0 1 4075
box -3 -3 3 3
use M3_M2  M3_M2_11054
timestamp 1745462530
transform 1 0 1108 0 1 4135
box -3 -3 3 3
use M3_M2  M3_M2_11055
timestamp 1745462530
transform 1 0 1108 0 1 4075
box -3 -3 3 3
use M3_M2  M3_M2_11056
timestamp 1745462530
transform 1 0 812 0 1 4155
box -3 -3 3 3
use M3_M2  M3_M2_11057
timestamp 1745462530
transform 1 0 764 0 1 4155
box -3 -3 3 3
use M3_M2  M3_M2_11058
timestamp 1745462530
transform 1 0 1372 0 1 4125
box -3 -3 3 3
use M3_M2  M3_M2_11059
timestamp 1745462530
transform 1 0 1028 0 1 4125
box -3 -3 3 3
use M3_M2  M3_M2_11060
timestamp 1745462530
transform 1 0 452 0 1 3995
box -3 -3 3 3
use M3_M2  M3_M2_11061
timestamp 1745462530
transform 1 0 388 0 1 3995
box -3 -3 3 3
use M3_M2  M3_M2_11062
timestamp 1745462530
transform 1 0 364 0 1 4045
box -3 -3 3 3
use M3_M2  M3_M2_11063
timestamp 1745462530
transform 1 0 324 0 1 4045
box -3 -3 3 3
use M3_M2  M3_M2_11064
timestamp 1745462530
transform 1 0 372 0 1 4015
box -3 -3 3 3
use M3_M2  M3_M2_11065
timestamp 1745462530
transform 1 0 300 0 1 4015
box -3 -3 3 3
use M3_M2  M3_M2_11066
timestamp 1745462530
transform 1 0 268 0 1 3945
box -3 -3 3 3
use M3_M2  M3_M2_11067
timestamp 1745462530
transform 1 0 84 0 1 3945
box -3 -3 3 3
use M3_M2  M3_M2_11068
timestamp 1745462530
transform 1 0 588 0 1 3955
box -3 -3 3 3
use M3_M2  M3_M2_11069
timestamp 1745462530
transform 1 0 508 0 1 3955
box -3 -3 3 3
use M3_M2  M3_M2_11070
timestamp 1745462530
transform 1 0 636 0 1 4045
box -3 -3 3 3
use M3_M2  M3_M2_11071
timestamp 1745462530
transform 1 0 612 0 1 4045
box -3 -3 3 3
use M3_M2  M3_M2_11072
timestamp 1745462530
transform 1 0 572 0 1 4045
box -3 -3 3 3
use M3_M2  M3_M2_11073
timestamp 1745462530
transform 1 0 684 0 1 3955
box -3 -3 3 3
use M3_M2  M3_M2_11074
timestamp 1745462530
transform 1 0 628 0 1 3955
box -3 -3 3 3
use M3_M2  M3_M2_11075
timestamp 1745462530
transform 1 0 220 0 1 4105
box -3 -3 3 3
use M3_M2  M3_M2_11076
timestamp 1745462530
transform 1 0 148 0 1 4125
box -3 -3 3 3
use M3_M2  M3_M2_11077
timestamp 1745462530
transform 1 0 148 0 1 4085
box -3 -3 3 3
use M3_M2  M3_M2_11078
timestamp 1745462530
transform 1 0 124 0 1 4085
box -3 -3 3 3
use M3_M2  M3_M2_11079
timestamp 1745462530
transform 1 0 1476 0 1 4135
box -3 -3 3 3
use M3_M2  M3_M2_11080
timestamp 1745462530
transform 1 0 1404 0 1 4135
box -3 -3 3 3
use M3_M2  M3_M2_11081
timestamp 1745462530
transform 1 0 1460 0 1 4115
box -3 -3 3 3
use M3_M2  M3_M2_11082
timestamp 1745462530
transform 1 0 1428 0 1 4115
box -3 -3 3 3
use M3_M2  M3_M2_11083
timestamp 1745462530
transform 1 0 4244 0 1 4105
box -3 -3 3 3
use M3_M2  M3_M2_11084
timestamp 1745462530
transform 1 0 4228 0 1 4105
box -3 -3 3 3
use M3_M2  M3_M2_11085
timestamp 1745462530
transform 1 0 4140 0 1 4125
box -3 -3 3 3
use M3_M2  M3_M2_11086
timestamp 1745462530
transform 1 0 4140 0 1 4105
box -3 -3 3 3
use M3_M2  M3_M2_11087
timestamp 1745462530
transform 1 0 3972 0 1 4225
box -3 -3 3 3
use M3_M2  M3_M2_11088
timestamp 1745462530
transform 1 0 3972 0 1 4135
box -3 -3 3 3
use M3_M2  M3_M2_11089
timestamp 1745462530
transform 1 0 1732 0 1 4125
box -3 -3 3 3
use M3_M2  M3_M2_11090
timestamp 1745462530
transform 1 0 1724 0 1 4225
box -3 -3 3 3
use M3_M2  M3_M2_11091
timestamp 1745462530
transform 1 0 1572 0 1 4125
box -3 -3 3 3
use M3_M2  M3_M2_11092
timestamp 1745462530
transform 1 0 1516 0 1 4125
box -3 -3 3 3
use M3_M2  M3_M2_11093
timestamp 1745462530
transform 1 0 1516 0 1 4065
box -3 -3 3 3
use M3_M2  M3_M2_11094
timestamp 1745462530
transform 1 0 1452 0 1 4065
box -3 -3 3 3
use M3_M2  M3_M2_11095
timestamp 1745462530
transform 1 0 860 0 1 4065
box -3 -3 3 3
use M3_M2  M3_M2_11096
timestamp 1745462530
transform 1 0 4172 0 1 4115
box -3 -3 3 3
use M3_M2  M3_M2_11097
timestamp 1745462530
transform 1 0 4084 0 1 4115
box -3 -3 3 3
use M3_M2  M3_M2_11098
timestamp 1745462530
transform 1 0 4084 0 1 4075
box -3 -3 3 3
use M3_M2  M3_M2_11099
timestamp 1745462530
transform 1 0 1780 0 1 4215
box -3 -3 3 3
use M3_M2  M3_M2_11100
timestamp 1745462530
transform 1 0 1780 0 1 4075
box -3 -3 3 3
use M3_M2  M3_M2_11101
timestamp 1745462530
transform 1 0 1532 0 1 4215
box -3 -3 3 3
use M3_M2  M3_M2_11102
timestamp 1745462530
transform 1 0 1532 0 1 4135
box -3 -3 3 3
use M3_M2  M3_M2_11103
timestamp 1745462530
transform 1 0 1476 0 1 4125
box -3 -3 3 3
use M3_M2  M3_M2_11104
timestamp 1745462530
transform 1 0 1468 0 1 4095
box -3 -3 3 3
use M3_M2  M3_M2_11105
timestamp 1745462530
transform 1 0 1100 0 1 4095
box -3 -3 3 3
use M3_M2  M3_M2_11106
timestamp 1745462530
transform 1 0 1860 0 1 4095
box -3 -3 3 3
use M3_M2  M3_M2_11107
timestamp 1745462530
transform 1 0 1484 0 1 4095
box -3 -3 3 3
use M3_M2  M3_M2_11108
timestamp 1745462530
transform 1 0 1884 0 1 4135
box -3 -3 3 3
use M3_M2  M3_M2_11109
timestamp 1745462530
transform 1 0 1844 0 1 4135
box -3 -3 3 3
use M3_M2  M3_M2_11110
timestamp 1745462530
transform 1 0 1908 0 1 4145
box -3 -3 3 3
use M3_M2  M3_M2_11111
timestamp 1745462530
transform 1 0 1868 0 1 4145
box -3 -3 3 3
use M3_M2  M3_M2_11112
timestamp 1745462530
transform 1 0 2036 0 1 4115
box -3 -3 3 3
use M3_M2  M3_M2_11113
timestamp 1745462530
transform 1 0 1868 0 1 4115
box -3 -3 3 3
use M3_M2  M3_M2_11114
timestamp 1745462530
transform 1 0 1868 0 1 4185
box -3 -3 3 3
use M3_M2  M3_M2_11115
timestamp 1745462530
transform 1 0 1828 0 1 4185
box -3 -3 3 3
use M3_M2  M3_M2_11116
timestamp 1745462530
transform 1 0 2140 0 1 4195
box -3 -3 3 3
use M3_M2  M3_M2_11117
timestamp 1745462530
transform 1 0 1812 0 1 4195
box -3 -3 3 3
use M3_M2  M3_M2_11118
timestamp 1745462530
transform 1 0 1540 0 1 4165
box -3 -3 3 3
use M3_M2  M3_M2_11119
timestamp 1745462530
transform 1 0 1484 0 1 4165
box -3 -3 3 3
use M3_M2  M3_M2_11120
timestamp 1745462530
transform 1 0 1908 0 1 4275
box -3 -3 3 3
use M3_M2  M3_M2_11121
timestamp 1745462530
transform 1 0 1532 0 1 4275
box -3 -3 3 3
use M3_M2  M3_M2_11122
timestamp 1745462530
transform 1 0 2020 0 1 4165
box -3 -3 3 3
use M3_M2  M3_M2_11123
timestamp 1745462530
transform 1 0 1892 0 1 4165
box -3 -3 3 3
use M3_M2  M3_M2_11124
timestamp 1745462530
transform 1 0 2180 0 1 4275
box -3 -3 3 3
use M3_M2  M3_M2_11125
timestamp 1745462530
transform 1 0 1924 0 1 4275
box -3 -3 3 3
use M3_M2  M3_M2_11126
timestamp 1745462530
transform 1 0 2308 0 1 4135
box -3 -3 3 3
use M3_M2  M3_M2_11127
timestamp 1745462530
transform 1 0 1996 0 1 4135
box -3 -3 3 3
use M3_M2  M3_M2_11128
timestamp 1745462530
transform 1 0 4140 0 1 4175
box -3 -3 3 3
use M3_M2  M3_M2_11129
timestamp 1745462530
transform 1 0 4116 0 1 4175
box -3 -3 3 3
use M3_M2  M3_M2_11130
timestamp 1745462530
transform 1 0 4100 0 1 4105
box -3 -3 3 3
use M3_M2  M3_M2_11131
timestamp 1745462530
transform 1 0 4044 0 1 4105
box -3 -3 3 3
use M3_M2  M3_M2_11132
timestamp 1745462530
transform 1 0 4028 0 1 4145
box -3 -3 3 3
use M3_M2  M3_M2_11133
timestamp 1745462530
transform 1 0 4012 0 1 4145
box -3 -3 3 3
use M3_M2  M3_M2_11134
timestamp 1745462530
transform 1 0 4020 0 1 4105
box -3 -3 3 3
use M3_M2  M3_M2_11135
timestamp 1745462530
transform 1 0 4004 0 1 4105
box -3 -3 3 3
use M3_M2  M3_M2_11136
timestamp 1745462530
transform 1 0 3948 0 1 4135
box -3 -3 3 3
use M3_M2  M3_M2_11137
timestamp 1745462530
transform 1 0 3348 0 1 4135
box -3 -3 3 3
use M3_M2  M3_M2_11138
timestamp 1745462530
transform 1 0 4012 0 1 4275
box -3 -3 3 3
use M3_M2  M3_M2_11139
timestamp 1745462530
transform 1 0 3836 0 1 4285
box -3 -3 3 3
use M3_M2  M3_M2_11140
timestamp 1745462530
transform 1 0 4236 0 1 3955
box -3 -3 3 3
use M3_M2  M3_M2_11141
timestamp 1745462530
transform 1 0 4196 0 1 3955
box -3 -3 3 3
use M3_M2  M3_M2_11142
timestamp 1745462530
transform 1 0 4196 0 1 3895
box -3 -3 3 3
use M3_M2  M3_M2_11143
timestamp 1745462530
transform 1 0 4076 0 1 3895
box -3 -3 3 3
use M3_M2  M3_M2_11144
timestamp 1745462530
transform 1 0 4044 0 1 3965
box -3 -3 3 3
use M3_M2  M3_M2_11145
timestamp 1745462530
transform 1 0 4012 0 1 3965
box -3 -3 3 3
use M3_M2  M3_M2_11146
timestamp 1745462530
transform 1 0 4092 0 1 3975
box -3 -3 3 3
use M3_M2  M3_M2_11147
timestamp 1745462530
transform 1 0 3956 0 1 3975
box -3 -3 3 3
use M3_M2  M3_M2_11148
timestamp 1745462530
transform 1 0 3924 0 1 4085
box -3 -3 3 3
use M3_M2  M3_M2_11149
timestamp 1745462530
transform 1 0 3660 0 1 4085
box -3 -3 3 3
use M3_M2  M3_M2_11150
timestamp 1745462530
transform 1 0 4068 0 1 3945
box -3 -3 3 3
use M3_M2  M3_M2_11151
timestamp 1745462530
transform 1 0 3996 0 1 3945
box -3 -3 3 3
use M3_M2  M3_M2_11152
timestamp 1745462530
transform 1 0 3988 0 1 4105
box -3 -3 3 3
use M3_M2  M3_M2_11153
timestamp 1745462530
transform 1 0 3788 0 1 4105
box -3 -3 3 3
use M3_M2  M3_M2_11154
timestamp 1745462530
transform 1 0 4204 0 1 4135
box -3 -3 3 3
use M3_M2  M3_M2_11155
timestamp 1745462530
transform 1 0 4164 0 1 4135
box -3 -3 3 3
use M3_M2  M3_M2_11156
timestamp 1745462530
transform 1 0 4132 0 1 4215
box -3 -3 3 3
use M3_M2  M3_M2_11157
timestamp 1745462530
transform 1 0 4068 0 1 4215
box -3 -3 3 3
use M3_M2  M3_M2_11158
timestamp 1745462530
transform 1 0 4076 0 1 4235
box -3 -3 3 3
use M3_M2  M3_M2_11159
timestamp 1745462530
transform 1 0 3468 0 1 4235
box -3 -3 3 3
use M3_M2  M3_M2_11160
timestamp 1745462530
transform 1 0 4028 0 1 4215
box -3 -3 3 3
use M3_M2  M3_M2_11161
timestamp 1745462530
transform 1 0 3876 0 1 4215
box -3 -3 3 3
use M3_M2  M3_M2_11162
timestamp 1745462530
transform 1 0 4236 0 1 3985
box -3 -3 3 3
use M3_M2  M3_M2_11163
timestamp 1745462530
transform 1 0 4196 0 1 3985
box -3 -3 3 3
use M3_M2  M3_M2_11164
timestamp 1745462530
transform 1 0 4196 0 1 4035
box -3 -3 3 3
use M3_M2  M3_M2_11165
timestamp 1745462530
transform 1 0 4100 0 1 4035
box -3 -3 3 3
use M3_M2  M3_M2_11166
timestamp 1745462530
transform 1 0 4132 0 1 4135
box -3 -3 3 3
use M3_M2  M3_M2_11167
timestamp 1745462530
transform 1 0 4044 0 1 4145
box -3 -3 3 3
use M3_M2  M3_M2_11168
timestamp 1745462530
transform 1 0 4052 0 1 4115
box -3 -3 3 3
use M3_M2  M3_M2_11169
timestamp 1745462530
transform 1 0 3604 0 1 4125
box -3 -3 3 3
use M3_M2  M3_M2_11170
timestamp 1745462530
transform 1 0 4116 0 1 4005
box -3 -3 3 3
use M3_M2  M3_M2_11171
timestamp 1745462530
transform 1 0 4020 0 1 4005
box -3 -3 3 3
use M3_M2  M3_M2_11172
timestamp 1745462530
transform 1 0 4004 0 1 4035
box -3 -3 3 3
use M3_M2  M3_M2_11173
timestamp 1745462530
transform 1 0 3828 0 1 4045
box -3 -3 3 3
use M3_M2  M3_M2_11174
timestamp 1745462530
transform 1 0 1788 0 1 4155
box -3 -3 3 3
use M3_M2  M3_M2_11175
timestamp 1745462530
transform 1 0 1580 0 1 4155
box -3 -3 3 3
use M3_M2  M3_M2_11176
timestamp 1745462530
transform 1 0 2876 0 1 4275
box -3 -3 3 3
use M3_M2  M3_M2_11177
timestamp 1745462530
transform 1 0 2836 0 1 4275
box -3 -3 3 3
use M3_M2  M3_M2_11178
timestamp 1745462530
transform 1 0 2836 0 1 4255
box -3 -3 3 3
use M3_M2  M3_M2_11179
timestamp 1745462530
transform 1 0 1788 0 1 4255
box -3 -3 3 3
use M3_M2  M3_M2_11180
timestamp 1745462530
transform 1 0 2996 0 1 4255
box -3 -3 3 3
use M3_M2  M3_M2_11181
timestamp 1745462530
transform 1 0 2852 0 1 4255
box -3 -3 3 3
use M3_M2  M3_M2_11182
timestamp 1745462530
transform 1 0 3052 0 1 4275
box -3 -3 3 3
use M3_M2  M3_M2_11183
timestamp 1745462530
transform 1 0 2892 0 1 4275
box -3 -3 3 3
use M3_M2  M3_M2_11184
timestamp 1745462530
transform 1 0 3012 0 1 4215
box -3 -3 3 3
use M3_M2  M3_M2_11185
timestamp 1745462530
transform 1 0 2980 0 1 4215
box -3 -3 3 3
use M3_M2  M3_M2_11186
timestamp 1745462530
transform 1 0 1812 0 1 4185
box -3 -3 3 3
use M3_M2  M3_M2_11187
timestamp 1745462530
transform 1 0 1740 0 1 4185
box -3 -3 3 3
use M3_M2  M3_M2_11188
timestamp 1745462530
transform 1 0 2532 0 1 4215
box -3 -3 3 3
use M3_M2  M3_M2_11189
timestamp 1745462530
transform 1 0 1828 0 1 4215
box -3 -3 3 3
use M3_M2  M3_M2_11190
timestamp 1745462530
transform 1 0 2604 0 1 4205
box -3 -3 3 3
use M3_M2  M3_M2_11191
timestamp 1745462530
transform 1 0 2540 0 1 4205
box -3 -3 3 3
use M3_M2  M3_M2_11192
timestamp 1745462530
transform 1 0 2668 0 1 4215
box -3 -3 3 3
use M3_M2  M3_M2_11193
timestamp 1745462530
transform 1 0 2548 0 1 4215
box -3 -3 3 3
use M3_M2  M3_M2_11194
timestamp 1745462530
transform 1 0 2820 0 1 4205
box -3 -3 3 3
use M3_M2  M3_M2_11195
timestamp 1745462530
transform 1 0 2652 0 1 4205
box -3 -3 3 3
use M3_M2  M3_M2_11196
timestamp 1745462530
transform 1 0 2692 0 1 4285
box -3 -3 3 3
use M3_M2  M3_M2_11197
timestamp 1745462530
transform 1 0 2588 0 1 4275
box -3 -3 3 3
use M3_M2  M3_M2_11198
timestamp 1745462530
transform 1 0 1524 0 1 4115
box -3 -3 3 3
use M3_M2  M3_M2_11199
timestamp 1745462530
transform 1 0 1244 0 1 4105
box -3 -3 3 3
use M3_M2  M3_M2_11200
timestamp 1745462530
transform 1 0 1188 0 1 4105
box -3 -3 3 3
use M3_M2  M3_M2_11201
timestamp 1745462530
transform 1 0 1124 0 1 4105
box -3 -3 3 3
use M3_M2  M3_M2_11202
timestamp 1745462530
transform 1 0 1380 0 1 4115
box -3 -3 3 3
use M3_M2  M3_M2_11203
timestamp 1745462530
transform 1 0 1212 0 1 4115
box -3 -3 3 3
use M3_M2  M3_M2_11204
timestamp 1745462530
transform 1 0 1156 0 1 4115
box -3 -3 3 3
use M3_M2  M3_M2_11205
timestamp 1745462530
transform 1 0 1060 0 1 4115
box -3 -3 3 3
use M3_M2  M3_M2_11206
timestamp 1745462530
transform 1 0 1364 0 1 4015
box -3 -3 3 3
use M3_M2  M3_M2_11207
timestamp 1745462530
transform 1 0 1308 0 1 4015
box -3 -3 3 3
use M3_M2  M3_M2_11208
timestamp 1745462530
transform 1 0 1180 0 1 4015
box -3 -3 3 3
use M3_M2  M3_M2_11209
timestamp 1745462530
transform 1 0 1140 0 1 4015
box -3 -3 3 3
use M3_M2  M3_M2_11210
timestamp 1745462530
transform 1 0 1236 0 1 3955
box -3 -3 3 3
use M3_M2  M3_M2_11211
timestamp 1745462530
transform 1 0 1180 0 1 3955
box -3 -3 3 3
use M3_M2  M3_M2_11212
timestamp 1745462530
transform 1 0 1028 0 1 3955
box -3 -3 3 3
use M3_M2  M3_M2_11213
timestamp 1745462530
transform 1 0 788 0 1 3955
box -3 -3 3 3
use M3_M2  M3_M2_11214
timestamp 1745462530
transform 1 0 1228 0 1 4025
box -3 -3 3 3
use M3_M2  M3_M2_11215
timestamp 1745462530
transform 1 0 1164 0 1 4025
box -3 -3 3 3
use M3_M2  M3_M2_11216
timestamp 1745462530
transform 1 0 1276 0 1 3995
box -3 -3 3 3
use M3_M2  M3_M2_11217
timestamp 1745462530
transform 1 0 1244 0 1 3995
box -3 -3 3 3
use M3_M2  M3_M2_11218
timestamp 1745462530
transform 1 0 660 0 1 4105
box -3 -3 3 3
use M3_M2  M3_M2_11219
timestamp 1745462530
transform 1 0 548 0 1 4105
box -3 -3 3 3
use M3_M2  M3_M2_11220
timestamp 1745462530
transform 1 0 596 0 1 4205
box -3 -3 3 3
use M3_M2  M3_M2_11221
timestamp 1745462530
transform 1 0 516 0 1 4205
box -3 -3 3 3
use M3_M2  M3_M2_11222
timestamp 1745462530
transform 1 0 980 0 1 4005
box -3 -3 3 3
use M3_M2  M3_M2_11223
timestamp 1745462530
transform 1 0 908 0 1 4005
box -3 -3 3 3
use M3_M2  M3_M2_11224
timestamp 1745462530
transform 1 0 924 0 1 4185
box -3 -3 3 3
use M3_M2  M3_M2_11225
timestamp 1745462530
transform 1 0 876 0 1 4185
box -3 -3 3 3
use M3_M2  M3_M2_11226
timestamp 1745462530
transform 1 0 804 0 1 3325
box -3 -3 3 3
use M3_M2  M3_M2_11227
timestamp 1745462530
transform 1 0 772 0 1 3325
box -3 -3 3 3
use M3_M2  M3_M2_11228
timestamp 1745462530
transform 1 0 404 0 1 3325
box -3 -3 3 3
use M3_M2  M3_M2_11229
timestamp 1745462530
transform 1 0 524 0 1 3365
box -3 -3 3 3
use M3_M2  M3_M2_11230
timestamp 1745462530
transform 1 0 276 0 1 3365
box -3 -3 3 3
use M3_M2  M3_M2_11231
timestamp 1745462530
transform 1 0 228 0 1 3355
box -3 -3 3 3
use M3_M2  M3_M2_11232
timestamp 1745462530
transform 1 0 652 0 1 3445
box -3 -3 3 3
use M3_M2  M3_M2_11233
timestamp 1745462530
transform 1 0 340 0 1 3505
box -3 -3 3 3
use M3_M2  M3_M2_11234
timestamp 1745462530
transform 1 0 340 0 1 3445
box -3 -3 3 3
use M3_M2  M3_M2_11235
timestamp 1745462530
transform 1 0 236 0 1 3505
box -3 -3 3 3
use M3_M2  M3_M2_11236
timestamp 1745462530
transform 1 0 156 0 1 3505
box -3 -3 3 3
use M3_M2  M3_M2_11237
timestamp 1745462530
transform 1 0 84 0 1 3505
box -3 -3 3 3
use M3_M2  M3_M2_11238
timestamp 1745462530
transform 1 0 524 0 1 3425
box -3 -3 3 3
use M3_M2  M3_M2_11239
timestamp 1745462530
transform 1 0 220 0 1 3415
box -3 -3 3 3
use M3_M2  M3_M2_11240
timestamp 1745462530
transform 1 0 164 0 1 3415
box -3 -3 3 3
use M3_M2  M3_M2_11241
timestamp 1745462530
transform 1 0 604 0 1 3595
box -3 -3 3 3
use M3_M2  M3_M2_11242
timestamp 1745462530
transform 1 0 220 0 1 3595
box -3 -3 3 3
use M3_M2  M3_M2_11243
timestamp 1745462530
transform 1 0 180 0 1 3585
box -3 -3 3 3
use M3_M2  M3_M2_11244
timestamp 1745462530
transform 1 0 660 0 1 3625
box -3 -3 3 3
use M3_M2  M3_M2_11245
timestamp 1745462530
transform 1 0 372 0 1 3615
box -3 -3 3 3
use M3_M2  M3_M2_11246
timestamp 1745462530
transform 1 0 340 0 1 3615
box -3 -3 3 3
use M3_M2  M3_M2_11247
timestamp 1745462530
transform 1 0 244 0 1 3625
box -3 -3 3 3
use M3_M2  M3_M2_11248
timestamp 1745462530
transform 1 0 484 0 1 3565
box -3 -3 3 3
use M3_M2  M3_M2_11249
timestamp 1745462530
transform 1 0 484 0 1 3495
box -3 -3 3 3
use M3_M2  M3_M2_11250
timestamp 1745462530
transform 1 0 404 0 1 3495
box -3 -3 3 3
use M3_M2  M3_M2_11251
timestamp 1745462530
transform 1 0 324 0 1 3565
box -3 -3 3 3
use M3_M2  M3_M2_11252
timestamp 1745462530
transform 1 0 2868 0 1 3825
box -3 -3 3 3
use M3_M2  M3_M2_11253
timestamp 1745462530
transform 1 0 2812 0 1 3825
box -3 -3 3 3
use M3_M2  M3_M2_11254
timestamp 1745462530
transform 1 0 3148 0 1 4255
box -3 -3 3 3
use M3_M2  M3_M2_11255
timestamp 1745462530
transform 1 0 3148 0 1 3845
box -3 -3 3 3
use M3_M2  M3_M2_11256
timestamp 1745462530
transform 1 0 3100 0 1 3845
box -3 -3 3 3
use M3_M2  M3_M2_11257
timestamp 1745462530
transform 1 0 3060 0 1 4255
box -3 -3 3 3
use M3_M2  M3_M2_11258
timestamp 1745462530
transform 1 0 3020 0 1 3845
box -3 -3 3 3
use M3_M2  M3_M2_11259
timestamp 1745462530
transform 1 0 3612 0 1 4215
box -3 -3 3 3
use M3_M2  M3_M2_11260
timestamp 1745462530
transform 1 0 3612 0 1 4085
box -3 -3 3 3
use M3_M2  M3_M2_11261
timestamp 1745462530
transform 1 0 3540 0 1 4215
box -3 -3 3 3
use M3_M2  M3_M2_11262
timestamp 1745462530
transform 1 0 3436 0 1 4085
box -3 -3 3 3
use M3_M2  M3_M2_11263
timestamp 1745462530
transform 1 0 3524 0 1 4265
box -3 -3 3 3
use M3_M2  M3_M2_11264
timestamp 1745462530
transform 1 0 3452 0 1 4015
box -3 -3 3 3
use M3_M2  M3_M2_11265
timestamp 1745462530
transform 1 0 3444 0 1 4265
box -3 -3 3 3
use M3_M2  M3_M2_11266
timestamp 1745462530
transform 1 0 3428 0 1 4015
box -3 -3 3 3
use M3_M2  M3_M2_11267
timestamp 1745462530
transform 1 0 3316 0 1 4015
box -3 -3 3 3
use M3_M2  M3_M2_11268
timestamp 1745462530
transform 1 0 3676 0 1 4285
box -3 -3 3 3
use M3_M2  M3_M2_11269
timestamp 1745462530
transform 1 0 3652 0 1 3845
box -3 -3 3 3
use M3_M2  M3_M2_11270
timestamp 1745462530
transform 1 0 3460 0 1 4285
box -3 -3 3 3
use M3_M2  M3_M2_11271
timestamp 1745462530
transform 1 0 3420 0 1 3845
box -3 -3 3 3
use M3_M2  M3_M2_11272
timestamp 1745462530
transform 1 0 3420 0 1 3795
box -3 -3 3 3
use M3_M2  M3_M2_11273
timestamp 1745462530
transform 1 0 3332 0 1 3795
box -3 -3 3 3
use M3_M2  M3_M2_11274
timestamp 1745462530
transform 1 0 3356 0 1 4105
box -3 -3 3 3
use M3_M2  M3_M2_11275
timestamp 1745462530
transform 1 0 3236 0 1 4105
box -3 -3 3 3
use M3_M2  M3_M2_11276
timestamp 1745462530
transform 1 0 3220 0 1 4105
box -3 -3 3 3
use M3_M2  M3_M2_11277
timestamp 1745462530
transform 1 0 2548 0 1 3975
box -3 -3 3 3
use M3_M2  M3_M2_11278
timestamp 1745462530
transform 1 0 2524 0 1 4205
box -3 -3 3 3
use M3_M2  M3_M2_11279
timestamp 1745462530
transform 1 0 2524 0 1 3975
box -3 -3 3 3
use M3_M2  M3_M2_11280
timestamp 1745462530
transform 1 0 2372 0 1 4205
box -3 -3 3 3
use M3_M2  M3_M2_11281
timestamp 1745462530
transform 1 0 2364 0 1 3975
box -3 -3 3 3
use M3_M2  M3_M2_11282
timestamp 1745462530
transform 1 0 2196 0 1 4195
box -3 -3 3 3
use M3_M2  M3_M2_11283
timestamp 1745462530
transform 1 0 2156 0 1 4105
box -3 -3 3 3
use M3_M2  M3_M2_11284
timestamp 1745462530
transform 1 0 2052 0 1 4115
box -3 -3 3 3
use M3_M2  M3_M2_11285
timestamp 1745462530
transform 1 0 2828 0 1 4045
box -3 -3 3 3
use M3_M2  M3_M2_11286
timestamp 1745462530
transform 1 0 2748 0 1 4285
box -3 -3 3 3
use M3_M2  M3_M2_11287
timestamp 1745462530
transform 1 0 2716 0 1 4045
box -3 -3 3 3
use M3_M2  M3_M2_11288
timestamp 1745462530
transform 1 0 2708 0 1 4285
box -3 -3 3 3
use M3_M2  M3_M2_11289
timestamp 1745462530
transform 1 0 3164 0 1 4295
box -3 -3 3 3
use M3_M2  M3_M2_11290
timestamp 1745462530
transform 1 0 3164 0 1 4045
box -3 -3 3 3
use M3_M2  M3_M2_11291
timestamp 1745462530
transform 1 0 3084 0 1 4295
box -3 -3 3 3
use M3_M2  M3_M2_11292
timestamp 1745462530
transform 1 0 3084 0 1 4045
box -3 -3 3 3
use M3_M2  M3_M2_11293
timestamp 1745462530
transform 1 0 3028 0 1 4295
box -3 -3 3 3
use M3_M2  M3_M2_11294
timestamp 1745462530
transform 1 0 3964 0 1 4295
box -3 -3 3 3
use M3_M2  M3_M2_11295
timestamp 1745462530
transform 1 0 3956 0 1 4125
box -3 -3 3 3
use M3_M2  M3_M2_11296
timestamp 1745462530
transform 1 0 3916 0 1 3865
box -3 -3 3 3
use M3_M2  M3_M2_11297
timestamp 1745462530
transform 1 0 3844 0 1 4125
box -3 -3 3 3
use M3_M2  M3_M2_11298
timestamp 1745462530
transform 1 0 3828 0 1 3865
box -3 -3 3 3
use M3_M2  M3_M2_11299
timestamp 1745462530
transform 1 0 3812 0 1 4295
box -3 -3 3 3
use M3_M2  M3_M2_11300
timestamp 1745462530
transform 1 0 3676 0 1 3865
box -3 -3 3 3
use M3_M2  M3_M2_11301
timestamp 1745462530
transform 1 0 3892 0 1 4165
box -3 -3 3 3
use M3_M2  M3_M2_11302
timestamp 1745462530
transform 1 0 3708 0 1 4165
box -3 -3 3 3
use M3_M2  M3_M2_11303
timestamp 1745462530
transform 1 0 3628 0 1 4165
box -3 -3 3 3
use M3_M2  M3_M2_11304
timestamp 1745462530
transform 1 0 3812 0 1 4045
box -3 -3 3 3
use M3_M2  M3_M2_11305
timestamp 1745462530
transform 1 0 3804 0 1 4125
box -3 -3 3 3
use M3_M2  M3_M2_11306
timestamp 1745462530
transform 1 0 3804 0 1 3785
box -3 -3 3 3
use M3_M2  M3_M2_11307
timestamp 1745462530
transform 1 0 3764 0 1 4125
box -3 -3 3 3
use M3_M2  M3_M2_11308
timestamp 1745462530
transform 1 0 3764 0 1 4045
box -3 -3 3 3
use M3_M2  M3_M2_11309
timestamp 1745462530
transform 1 0 3692 0 1 3785
box -3 -3 3 3
use M3_M2  M3_M2_11310
timestamp 1745462530
transform 1 0 3852 0 1 4325
box -3 -3 3 3
use M3_M2  M3_M2_11311
timestamp 1745462530
transform 1 0 3508 0 1 4325
box -3 -3 3 3
use M3_M2  M3_M2_11312
timestamp 1745462530
transform 1 0 3372 0 1 4325
box -3 -3 3 3
use M3_M2  M3_M2_11313
timestamp 1745462530
transform 1 0 3364 0 1 4215
box -3 -3 3 3
use M3_M2  M3_M2_11314
timestamp 1745462530
transform 1 0 3268 0 1 4215
box -3 -3 3 3
use M3_M2  M3_M2_11315
timestamp 1745462530
transform 1 0 2548 0 1 4095
box -3 -3 3 3
use M3_M2  M3_M2_11316
timestamp 1745462530
transform 1 0 2476 0 1 4295
box -3 -3 3 3
use M3_M2  M3_M2_11317
timestamp 1745462530
transform 1 0 2476 0 1 4095
box -3 -3 3 3
use M3_M2  M3_M2_11318
timestamp 1745462530
transform 1 0 2412 0 1 4295
box -3 -3 3 3
use M3_M2  M3_M2_11319
timestamp 1745462530
transform 1 0 2332 0 1 4295
box -3 -3 3 3
use M3_M2  M3_M2_11320
timestamp 1745462530
transform 1 0 2332 0 1 4005
box -3 -3 3 3
use M3_M2  M3_M2_11321
timestamp 1745462530
transform 1 0 2244 0 1 4295
box -3 -3 3 3
use M3_M2  M3_M2_11322
timestamp 1745462530
transform 1 0 2212 0 1 4005
box -3 -3 3 3
use M3_M2  M3_M2_11323
timestamp 1745462530
transform 1 0 2156 0 1 4295
box -3 -3 3 3
use M3_M2  M3_M2_11324
timestamp 1745462530
transform 1 0 2140 0 1 4005
box -3 -3 3 3
use M3_M2  M3_M2_11325
timestamp 1745462530
transform 1 0 2892 0 1 4145
box -3 -3 3 3
use M3_M2  M3_M2_11326
timestamp 1745462530
transform 1 0 2812 0 1 4145
box -3 -3 3 3
use M3_M2  M3_M2_11327
timestamp 1745462530
transform 1 0 2780 0 1 4145
box -3 -3 3 3
use M3_M2  M3_M2_11328
timestamp 1745462530
transform 1 0 3172 0 1 4215
box -3 -3 3 3
use M3_M2  M3_M2_11329
timestamp 1745462530
transform 1 0 3076 0 1 4215
box -3 -3 3 3
use M3_M2  M3_M2_11330
timestamp 1745462530
transform 1 0 3036 0 1 4215
box -3 -3 3 3
use M3_M2  M3_M2_11331
timestamp 1745462530
transform 1 0 3716 0 1 4035
box -3 -3 3 3
use M3_M2  M3_M2_11332
timestamp 1745462530
transform 1 0 3644 0 1 4105
box -3 -3 3 3
use M3_M2  M3_M2_11333
timestamp 1745462530
transform 1 0 3636 0 1 4035
box -3 -3 3 3
use M3_M2  M3_M2_11334
timestamp 1745462530
transform 1 0 3588 0 1 4105
box -3 -3 3 3
use M3_M2  M3_M2_11335
timestamp 1745462530
transform 1 0 2436 0 1 4305
box -3 -3 3 3
use M3_M2  M3_M2_11336
timestamp 1745462530
transform 1 0 2380 0 1 4305
box -3 -3 3 3
use M3_M2  M3_M2_11337
timestamp 1745462530
transform 1 0 2324 0 1 4305
box -3 -3 3 3
use M3_M2  M3_M2_11338
timestamp 1745462530
transform 1 0 2164 0 1 4305
box -3 -3 3 3
use M3_M2  M3_M2_11339
timestamp 1745462530
transform 1 0 2156 0 1 4145
box -3 -3 3 3
use M3_M2  M3_M2_11340
timestamp 1745462530
transform 1 0 2116 0 1 4145
box -3 -3 3 3
use M3_M2  M3_M2_11341
timestamp 1745462530
transform 1 0 2020 0 1 4145
box -3 -3 3 3
use M3_M2  M3_M2_11342
timestamp 1745462530
transform 1 0 2796 0 1 4215
box -3 -3 3 3
use M3_M2  M3_M2_11343
timestamp 1745462530
transform 1 0 2724 0 1 4215
box -3 -3 3 3
use M3_M2  M3_M2_11344
timestamp 1745462530
transform 1 0 2684 0 1 4145
box -3 -3 3 3
use M3_M2  M3_M2_11345
timestamp 1745462530
transform 1 0 2668 0 1 4145
box -3 -3 3 3
use M3_M2  M3_M2_11346
timestamp 1745462530
transform 1 0 2996 0 1 4265
box -3 -3 3 3
use M3_M2  M3_M2_11347
timestamp 1745462530
transform 1 0 2996 0 1 4195
box -3 -3 3 3
use M3_M2  M3_M2_11348
timestamp 1745462530
transform 1 0 2948 0 1 4265
box -3 -3 3 3
use M3_M2  M3_M2_11349
timestamp 1745462530
transform 1 0 2948 0 1 4195
box -3 -3 3 3
use M3_M2  M3_M2_11350
timestamp 1745462530
transform 1 0 3916 0 1 4015
box -3 -3 3 3
use M3_M2  M3_M2_11351
timestamp 1745462530
transform 1 0 3804 0 1 4015
box -3 -3 3 3
use M3_M2  M3_M2_11352
timestamp 1745462530
transform 1 0 4004 0 1 4285
box -3 -3 3 3
use M3_M2  M3_M2_11353
timestamp 1745462530
transform 1 0 3924 0 1 4285
box -3 -3 3 3
use M3_M2  M3_M2_11354
timestamp 1745462530
transform 1 0 3844 0 1 3895
box -3 -3 3 3
use M3_M2  M3_M2_11355
timestamp 1745462530
transform 1 0 3772 0 1 4105
box -3 -3 3 3
use M3_M2  M3_M2_11356
timestamp 1745462530
transform 1 0 3756 0 1 4105
box -3 -3 3 3
use M3_M2  M3_M2_11357
timestamp 1745462530
transform 1 0 3732 0 1 3895
box -3 -3 3 3
use M3_M2  M3_M2_11358
timestamp 1745462530
transform 1 0 3820 0 1 4185
box -3 -3 3 3
use M3_M2  M3_M2_11359
timestamp 1745462530
transform 1 0 3796 0 1 4185
box -3 -3 3 3
use M3_M2  M3_M2_11360
timestamp 1745462530
transform 1 0 3748 0 1 4185
box -3 -3 3 3
use M3_M2  M3_M2_11361
timestamp 1745462530
transform 1 0 2524 0 1 4275
box -3 -3 3 3
use M3_M2  M3_M2_11362
timestamp 1745462530
transform 1 0 2468 0 1 4275
box -3 -3 3 3
use M3_M2  M3_M2_11363
timestamp 1745462530
transform 1 0 2396 0 1 4275
box -3 -3 3 3
use M3_M2  M3_M2_11364
timestamp 1745462530
transform 1 0 2300 0 1 4275
box -3 -3 3 3
use M3_M2  M3_M2_11365
timestamp 1745462530
transform 1 0 2292 0 1 4285
box -3 -3 3 3
use M3_M2  M3_M2_11366
timestamp 1745462530
transform 1 0 2268 0 1 4145
box -3 -3 3 3
use M3_M2  M3_M2_11367
timestamp 1745462530
transform 1 0 2252 0 1 4285
box -3 -3 3 3
use M3_M2  M3_M2_11368
timestamp 1745462530
transform 1 0 2252 0 1 4145
box -3 -3 3 3
use M3_M2  M3_M2_11369
timestamp 1745462530
transform 1 0 2228 0 1 4285
box -3 -3 3 3
use M3_M2  M3_M2_11370
timestamp 1745462530
transform 1 0 2124 0 1 4285
box -3 -3 3 3
use M3_M2  M3_M2_11371
timestamp 1745462530
transform 1 0 2620 0 1 4045
box -3 -3 3 3
use M3_M2  M3_M2_11372
timestamp 1745462530
transform 1 0 2564 0 1 4045
box -3 -3 3 3
use M3_M2  M3_M2_11373
timestamp 1745462530
transform 1 0 2948 0 1 3985
box -3 -3 3 3
use M3_M2  M3_M2_11374
timestamp 1745462530
transform 1 0 2932 0 1 3985
box -3 -3 3 3
use M3_M2  M3_M2_11375
timestamp 1745462530
transform 1 0 2900 0 1 3985
box -3 -3 3 3
use M3_M2  M3_M2_11376
timestamp 1745462530
transform 1 0 4356 0 1 3815
box -3 -3 3 3
use M3_M2  M3_M2_11377
timestamp 1745462530
transform 1 0 4124 0 1 3825
box -3 -3 3 3
use M3_M2  M3_M2_11378
timestamp 1745462530
transform 1 0 4364 0 1 3935
box -3 -3 3 3
use M3_M2  M3_M2_11379
timestamp 1745462530
transform 1 0 4260 0 1 3935
box -3 -3 3 3
use M3_M2  M3_M2_11380
timestamp 1745462530
transform 1 0 4260 0 1 3805
box -3 -3 3 3
use M3_M2  M3_M2_11381
timestamp 1745462530
transform 1 0 4108 0 1 3935
box -3 -3 3 3
use M3_M2  M3_M2_11382
timestamp 1745462530
transform 1 0 4100 0 1 3805
box -3 -3 3 3
use M3_M2  M3_M2_11383
timestamp 1745462530
transform 1 0 4372 0 1 3775
box -3 -3 3 3
use M3_M2  M3_M2_11384
timestamp 1745462530
transform 1 0 4372 0 1 3595
box -3 -3 3 3
use M3_M2  M3_M2_11385
timestamp 1745462530
transform 1 0 4268 0 1 3595
box -3 -3 3 3
use M3_M2  M3_M2_11386
timestamp 1745462530
transform 1 0 4100 0 1 3845
box -3 -3 3 3
use M3_M2  M3_M2_11387
timestamp 1745462530
transform 1 0 4076 0 1 3785
box -3 -3 3 3
use M3_M2  M3_M2_11388
timestamp 1745462530
transform 1 0 4068 0 1 3845
box -3 -3 3 3
use M3_M2  M3_M2_11389
timestamp 1745462530
transform 1 0 4004 0 1 3615
box -3 -3 3 3
use M3_M2  M3_M2_11390
timestamp 1745462530
transform 1 0 3996 0 1 3805
box -3 -3 3 3
use M3_M2  M3_M2_11391
timestamp 1745462530
transform 1 0 3980 0 1 3805
box -3 -3 3 3
use M3_M2  M3_M2_11392
timestamp 1745462530
transform 1 0 3980 0 1 3615
box -3 -3 3 3
use M3_M2  M3_M2_11393
timestamp 1745462530
transform 1 0 3972 0 1 4095
box -3 -3 3 3
use M3_M2  M3_M2_11394
timestamp 1745462530
transform 1 0 3924 0 1 4095
box -3 -3 3 3
use M3_M2  M3_M2_11395
timestamp 1745462530
transform 1 0 3908 0 1 3615
box -3 -3 3 3
use M3_M2  M3_M2_11396
timestamp 1745462530
transform 1 0 1964 0 1 4145
box -3 -3 3 3
use M3_M2  M3_M2_11397
timestamp 1745462530
transform 1 0 1948 0 1 4145
box -3 -3 3 3
use M3_M2  M3_M2_11398
timestamp 1745462530
transform 1 0 2076 0 1 4005
box -3 -3 3 3
use M3_M2  M3_M2_11399
timestamp 1745462530
transform 1 0 2044 0 1 4005
box -3 -3 3 3
use M3_M2  M3_M2_11400
timestamp 1745462530
transform 1 0 2012 0 1 4185
box -3 -3 3 3
use M3_M2  M3_M2_11401
timestamp 1745462530
transform 1 0 2012 0 1 4005
box -3 -3 3 3
use M3_M2  M3_M2_11402
timestamp 1745462530
transform 1 0 1900 0 1 4185
box -3 -3 3 3
use M3_M2  M3_M2_11403
timestamp 1745462530
transform 1 0 2660 0 1 3935
box -3 -3 3 3
use M3_M2  M3_M2_11404
timestamp 1745462530
transform 1 0 2580 0 1 3995
box -3 -3 3 3
use M3_M2  M3_M2_11405
timestamp 1745462530
transform 1 0 2564 0 1 3995
box -3 -3 3 3
use M3_M2  M3_M2_11406
timestamp 1745462530
transform 1 0 2564 0 1 3935
box -3 -3 3 3
use M3_M2  M3_M2_11407
timestamp 1745462530
transform 1 0 2996 0 1 3825
box -3 -3 3 3
use M3_M2  M3_M2_11408
timestamp 1745462530
transform 1 0 2980 0 1 3935
box -3 -3 3 3
use M3_M2  M3_M2_11409
timestamp 1745462530
transform 1 0 2980 0 1 3825
box -3 -3 3 3
use M3_M2  M3_M2_11410
timestamp 1745462530
transform 1 0 2940 0 1 3935
box -3 -3 3 3
use M3_M2  M3_M2_11411
timestamp 1745462530
transform 1 0 2884 0 1 3825
box -3 -3 3 3
use M3_M2  M3_M2_11412
timestamp 1745462530
transform 1 0 4244 0 1 3565
box -3 -3 3 3
use M3_M2  M3_M2_11413
timestamp 1745462530
transform 1 0 4140 0 1 3715
box -3 -3 3 3
use M3_M2  M3_M2_11414
timestamp 1745462530
transform 1 0 4108 0 1 3565
box -3 -3 3 3
use M3_M2  M3_M2_11415
timestamp 1745462530
transform 1 0 4100 0 1 3715
box -3 -3 3 3
use M3_M2  M3_M2_11416
timestamp 1745462530
transform 1 0 4204 0 1 3735
box -3 -3 3 3
use M3_M2  M3_M2_11417
timestamp 1745462530
transform 1 0 4092 0 1 3735
box -3 -3 3 3
use M3_M2  M3_M2_11418
timestamp 1745462530
transform 1 0 4084 0 1 3965
box -3 -3 3 3
use M3_M2  M3_M2_11419
timestamp 1745462530
transform 1 0 4068 0 1 3735
box -3 -3 3 3
use M3_M2  M3_M2_11420
timestamp 1745462530
transform 1 0 4060 0 1 3965
box -3 -3 3 3
use M3_M2  M3_M2_11421
timestamp 1745462530
transform 1 0 4356 0 1 3675
box -3 -3 3 3
use M3_M2  M3_M2_11422
timestamp 1745462530
transform 1 0 4148 0 1 3675
box -3 -3 3 3
use M3_M2  M3_M2_11423
timestamp 1745462530
transform 1 0 4076 0 1 3935
box -3 -3 3 3
use M3_M2  M3_M2_11424
timestamp 1745462530
transform 1 0 4036 0 1 3675
box -3 -3 3 3
use M3_M2  M3_M2_11425
timestamp 1745462530
transform 1 0 4012 0 1 3935
box -3 -3 3 3
use M3_M2  M3_M2_11426
timestamp 1745462530
transform 1 0 4124 0 1 3405
box -3 -3 3 3
use M3_M2  M3_M2_11427
timestamp 1745462530
transform 1 0 4052 0 1 3695
box -3 -3 3 3
use M3_M2  M3_M2_11428
timestamp 1745462530
transform 1 0 4012 0 1 3405
box -3 -3 3 3
use M3_M2  M3_M2_11429
timestamp 1745462530
transform 1 0 3972 0 1 3695
box -3 -3 3 3
use M3_M2  M3_M2_11430
timestamp 1745462530
transform 1 0 2020 0 1 3775
box -3 -3 3 3
use M3_M2  M3_M2_11431
timestamp 1745462530
transform 1 0 1988 0 1 3775
box -3 -3 3 3
use M3_M2  M3_M2_11432
timestamp 1745462530
transform 1 0 2020 0 1 4105
box -3 -3 3 3
use M3_M2  M3_M2_11433
timestamp 1745462530
transform 1 0 1956 0 1 4285
box -3 -3 3 3
use M3_M2  M3_M2_11434
timestamp 1745462530
transform 1 0 1956 0 1 4105
box -3 -3 3 3
use M3_M2  M3_M2_11435
timestamp 1745462530
transform 1 0 1940 0 1 4285
box -3 -3 3 3
use M3_M2  M3_M2_11436
timestamp 1745462530
transform 1 0 1860 0 1 4285
box -3 -3 3 3
use M3_M2  M3_M2_11437
timestamp 1745462530
transform 1 0 1908 0 1 3965
box -3 -3 3 3
use M3_M2  M3_M2_11438
timestamp 1745462530
transform 1 0 1852 0 1 4265
box -3 -3 3 3
use M3_M2  M3_M2_11439
timestamp 1745462530
transform 1 0 1844 0 1 3995
box -3 -3 3 3
use M3_M2  M3_M2_11440
timestamp 1745462530
transform 1 0 1844 0 1 3965
box -3 -3 3 3
use M3_M2  M3_M2_11441
timestamp 1745462530
transform 1 0 1796 0 1 4265
box -3 -3 3 3
use M3_M2  M3_M2_11442
timestamp 1745462530
transform 1 0 1788 0 1 3995
box -3 -3 3 3
use M3_M2  M3_M2_11443
timestamp 1745462530
transform 1 0 1828 0 1 4115
box -3 -3 3 3
use M3_M2  M3_M2_11444
timestamp 1745462530
transform 1 0 1772 0 1 4115
box -3 -3 3 3
use M3_M2  M3_M2_11445
timestamp 1745462530
transform 1 0 4372 0 1 3345
box -3 -3 3 3
use M3_M2  M3_M2_11446
timestamp 1745462530
transform 1 0 4340 0 1 3625
box -3 -3 3 3
use M3_M2  M3_M2_11447
timestamp 1745462530
transform 1 0 4340 0 1 3345
box -3 -3 3 3
use M3_M2  M3_M2_11448
timestamp 1745462530
transform 1 0 4268 0 1 3875
box -3 -3 3 3
use M3_M2  M3_M2_11449
timestamp 1745462530
transform 1 0 4268 0 1 3345
box -3 -3 3 3
use M3_M2  M3_M2_11450
timestamp 1745462530
transform 1 0 4260 0 1 3635
box -3 -3 3 3
use M3_M2  M3_M2_11451
timestamp 1745462530
transform 1 0 4140 0 1 3875
box -3 -3 3 3
use M3_M2  M3_M2_11452
timestamp 1745462530
transform 1 0 4356 0 1 3415
box -3 -3 3 3
use M3_M2  M3_M2_11453
timestamp 1745462530
transform 1 0 4324 0 1 3685
box -3 -3 3 3
use M3_M2  M3_M2_11454
timestamp 1745462530
transform 1 0 4324 0 1 3415
box -3 -3 3 3
use M3_M2  M3_M2_11455
timestamp 1745462530
transform 1 0 4260 0 1 3415
box -3 -3 3 3
use M3_M2  M3_M2_11456
timestamp 1745462530
transform 1 0 4188 0 1 3685
box -3 -3 3 3
use M3_M2  M3_M2_11457
timestamp 1745462530
transform 1 0 4196 0 1 3525
box -3 -3 3 3
use M3_M2  M3_M2_11458
timestamp 1745462530
transform 1 0 4180 0 1 3645
box -3 -3 3 3
use M3_M2  M3_M2_11459
timestamp 1745462530
transform 1 0 4180 0 1 3225
box -3 -3 3 3
use M3_M2  M3_M2_11460
timestamp 1745462530
transform 1 0 4164 0 1 3985
box -3 -3 3 3
use M3_M2  M3_M2_11461
timestamp 1745462530
transform 1 0 4108 0 1 3775
box -3 -3 3 3
use M3_M2  M3_M2_11462
timestamp 1745462530
transform 1 0 4108 0 1 3645
box -3 -3 3 3
use M3_M2  M3_M2_11463
timestamp 1745462530
transform 1 0 4076 0 1 3225
box -3 -3 3 3
use M3_M2  M3_M2_11464
timestamp 1745462530
transform 1 0 4036 0 1 3775
box -3 -3 3 3
use M3_M2  M3_M2_11465
timestamp 1745462530
transform 1 0 4020 0 1 3985
box -3 -3 3 3
use M3_M2  M3_M2_11466
timestamp 1745462530
transform 1 0 4380 0 1 3855
box -3 -3 3 3
use M3_M2  M3_M2_11467
timestamp 1745462530
transform 1 0 4380 0 1 3645
box -3 -3 3 3
use M3_M2  M3_M2_11468
timestamp 1745462530
transform 1 0 4372 0 1 3425
box -3 -3 3 3
use M3_M2  M3_M2_11469
timestamp 1745462530
transform 1 0 4084 0 1 3865
box -3 -3 3 3
use M3_M2  M3_M2_11470
timestamp 1745462530
transform 1 0 4060 0 1 3865
box -3 -3 3 3
use M3_M2  M3_M2_11471
timestamp 1745462530
transform 1 0 4012 0 1 3385
box -3 -3 3 3
use M3_M2  M3_M2_11472
timestamp 1745462530
transform 1 0 1596 0 1 4245
box -3 -3 3 3
use M3_M2  M3_M2_11473
timestamp 1745462530
transform 1 0 1596 0 1 4205
box -3 -3 3 3
use M3_M2  M3_M2_11474
timestamp 1745462530
transform 1 0 1572 0 1 4245
box -3 -3 3 3
use M3_M2  M3_M2_11475
timestamp 1745462530
transform 1 0 1524 0 1 4205
box -3 -3 3 3
use M3_M2  M3_M2_11476
timestamp 1745462530
transform 1 0 1756 0 1 3995
box -3 -3 3 3
use M3_M2  M3_M2_11477
timestamp 1745462530
transform 1 0 1716 0 1 3995
box -3 -3 3 3
use M3_M2  M3_M2_11478
timestamp 1745462530
transform 1 0 1636 0 1 4055
box -3 -3 3 3
use M3_M2  M3_M2_11479
timestamp 1745462530
transform 1 0 1580 0 1 4055
box -3 -3 3 3
use M3_M2  M3_M2_11480
timestamp 1745462530
transform 1 0 4364 0 1 3145
box -3 -3 3 3
use M3_M2  M3_M2_11481
timestamp 1745462530
transform 1 0 4276 0 1 3495
box -3 -3 3 3
use M3_M2  M3_M2_11482
timestamp 1745462530
transform 1 0 4268 0 1 3145
box -3 -3 3 3
use M3_M2  M3_M2_11483
timestamp 1745462530
transform 1 0 4244 0 1 3145
box -3 -3 3 3
use M3_M2  M3_M2_11484
timestamp 1745462530
transform 1 0 4220 0 1 3945
box -3 -3 3 3
use M3_M2  M3_M2_11485
timestamp 1745462530
transform 1 0 4212 0 1 3495
box -3 -3 3 3
use M3_M2  M3_M2_11486
timestamp 1745462530
transform 1 0 4204 0 1 3945
box -3 -3 3 3
use M3_M2  M3_M2_11487
timestamp 1745462530
transform 1 0 4380 0 1 3535
box -3 -3 3 3
use M3_M2  M3_M2_11488
timestamp 1745462530
transform 1 0 4364 0 1 3765
box -3 -3 3 3
use M3_M2  M3_M2_11489
timestamp 1745462530
transform 1 0 4364 0 1 3605
box -3 -3 3 3
use M3_M2  M3_M2_11490
timestamp 1745462530
transform 1 0 4364 0 1 3535
box -3 -3 3 3
use M3_M2  M3_M2_11491
timestamp 1745462530
transform 1 0 4364 0 1 3195
box -3 -3 3 3
use M3_M2  M3_M2_11492
timestamp 1745462530
transform 1 0 4332 0 1 4125
box -3 -3 3 3
use M3_M2  M3_M2_11493
timestamp 1745462530
transform 1 0 4332 0 1 3815
box -3 -3 3 3
use M3_M2  M3_M2_11494
timestamp 1745462530
transform 1 0 4332 0 1 3765
box -3 -3 3 3
use M3_M2  M3_M2_11495
timestamp 1745462530
transform 1 0 4260 0 1 3195
box -3 -3 3 3
use M3_M2  M3_M2_11496
timestamp 1745462530
transform 1 0 4220 0 1 4125
box -3 -3 3 3
use M3_M2  M3_M2_11497
timestamp 1745462530
transform 1 0 4132 0 1 3815
box -3 -3 3 3
use M3_M2  M3_M2_11498
timestamp 1745462530
transform 1 0 4204 0 1 3835
box -3 -3 3 3
use M3_M2  M3_M2_11499
timestamp 1745462530
transform 1 0 4196 0 1 3345
box -3 -3 3 3
use M3_M2  M3_M2_11500
timestamp 1745462530
transform 1 0 4148 0 1 3835
box -3 -3 3 3
use M3_M2  M3_M2_11501
timestamp 1745462530
transform 1 0 4148 0 1 3545
box -3 -3 3 3
use M3_M2  M3_M2_11502
timestamp 1745462530
transform 1 0 4116 0 1 3545
box -3 -3 3 3
use M3_M2  M3_M2_11503
timestamp 1745462530
transform 1 0 4116 0 1 3345
box -3 -3 3 3
use M3_M2  M3_M2_11504
timestamp 1745462530
transform 1 0 4092 0 1 3345
box -3 -3 3 3
use M3_M2  M3_M2_11505
timestamp 1745462530
transform 1 0 4156 0 1 4015
box -3 -3 3 3
use M3_M2  M3_M2_11506
timestamp 1745462530
transform 1 0 4156 0 1 3845
box -3 -3 3 3
use M3_M2  M3_M2_11507
timestamp 1745462530
transform 1 0 4116 0 1 4015
box -3 -3 3 3
use M3_M2  M3_M2_11508
timestamp 1745462530
transform 1 0 4020 0 1 3835
box -3 -3 3 3
use M3_M2  M3_M2_11509
timestamp 1745462530
transform 1 0 4020 0 1 3775
box -3 -3 3 3
use M3_M2  M3_M2_11510
timestamp 1745462530
transform 1 0 3988 0 1 3775
box -3 -3 3 3
use M3_M2  M3_M2_11511
timestamp 1745462530
transform 1 0 3988 0 1 3745
box -3 -3 3 3
use M3_M2  M3_M2_11512
timestamp 1745462530
transform 1 0 3876 0 1 3745
box -3 -3 3 3
use M3_M2  M3_M2_11513
timestamp 1745462530
transform 1 0 1540 0 1 4055
box -3 -3 3 3
use M3_M2  M3_M2_11514
timestamp 1745462530
transform 1 0 1492 0 1 4055
box -3 -3 3 3
use M3_M2  M3_M2_11515
timestamp 1745462530
transform 1 0 1548 0 1 3825
box -3 -3 3 3
use M3_M2  M3_M2_11516
timestamp 1745462530
transform 1 0 1468 0 1 4145
box -3 -3 3 3
use M3_M2  M3_M2_11517
timestamp 1745462530
transform 1 0 1428 0 1 3825
box -3 -3 3 3
use M3_M2  M3_M2_11518
timestamp 1745462530
transform 1 0 1420 0 1 4145
box -3 -3 3 3
use M3_M2  M3_M2_11519
timestamp 1745462530
transform 1 0 692 0 1 4035
box -3 -3 3 3
use M3_M2  M3_M2_11520
timestamp 1745462530
transform 1 0 636 0 1 3805
box -3 -3 3 3
use M3_M2  M3_M2_11521
timestamp 1745462530
transform 1 0 604 0 1 4255
box -3 -3 3 3
use M3_M2  M3_M2_11522
timestamp 1745462530
transform 1 0 588 0 1 4035
box -3 -3 3 3
use M3_M2  M3_M2_11523
timestamp 1745462530
transform 1 0 564 0 1 3935
box -3 -3 3 3
use M3_M2  M3_M2_11524
timestamp 1745462530
transform 1 0 564 0 1 3805
box -3 -3 3 3
use M3_M2  M3_M2_11525
timestamp 1745462530
transform 1 0 556 0 1 4255
box -3 -3 3 3
use M3_M2  M3_M2_11526
timestamp 1745462530
transform 1 0 556 0 1 4035
box -3 -3 3 3
use M3_M2  M3_M2_11527
timestamp 1745462530
transform 1 0 540 0 1 3935
box -3 -3 3 3
use M3_M2  M3_M2_11528
timestamp 1745462530
transform 1 0 700 0 1 4025
box -3 -3 3 3
use M3_M2  M3_M2_11529
timestamp 1745462530
transform 1 0 636 0 1 4285
box -3 -3 3 3
use M3_M2  M3_M2_11530
timestamp 1745462530
transform 1 0 596 0 1 4025
box -3 -3 3 3
use M3_M2  M3_M2_11531
timestamp 1745462530
transform 1 0 532 0 1 4285
box -3 -3 3 3
use M3_M2  M3_M2_11532
timestamp 1745462530
transform 1 0 516 0 1 4025
box -3 -3 3 3
use M3_M2  M3_M2_11533
timestamp 1745462530
transform 1 0 1236 0 1 3785
box -3 -3 3 3
use M3_M2  M3_M2_11534
timestamp 1745462530
transform 1 0 1212 0 1 3785
box -3 -3 3 3
use M3_M2  M3_M2_11535
timestamp 1745462530
transform 1 0 1164 0 1 3785
box -3 -3 3 3
use M3_M2  M3_M2_11536
timestamp 1745462530
transform 1 0 708 0 1 4245
box -3 -3 3 3
use M3_M2  M3_M2_11537
timestamp 1745462530
transform 1 0 460 0 1 3845
box -3 -3 3 3
use M3_M2  M3_M2_11538
timestamp 1745462530
transform 1 0 460 0 1 3785
box -3 -3 3 3
use M3_M2  M3_M2_11539
timestamp 1745462530
transform 1 0 108 0 1 4245
box -3 -3 3 3
use M3_M2  M3_M2_11540
timestamp 1745462530
transform 1 0 108 0 1 3845
box -3 -3 3 3
use M3_M2  M3_M2_11541
timestamp 1745462530
transform 1 0 68 0 1 3845
box -3 -3 3 3
use M3_M2  M3_M2_11542
timestamp 1745462530
transform 1 0 1300 0 1 3795
box -3 -3 3 3
use M3_M2  M3_M2_11543
timestamp 1745462530
transform 1 0 1196 0 1 3865
box -3 -3 3 3
use M3_M2  M3_M2_11544
timestamp 1745462530
transform 1 0 1196 0 1 3795
box -3 -3 3 3
use M3_M2  M3_M2_11545
timestamp 1745462530
transform 1 0 724 0 1 4235
box -3 -3 3 3
use M3_M2  M3_M2_11546
timestamp 1745462530
transform 1 0 476 0 1 3865
box -3 -3 3 3
use M3_M2  M3_M2_11547
timestamp 1745462530
transform 1 0 428 0 1 3975
box -3 -3 3 3
use M3_M2  M3_M2_11548
timestamp 1745462530
transform 1 0 404 0 1 3975
box -3 -3 3 3
use M3_M2  M3_M2_11549
timestamp 1745462530
transform 1 0 396 0 1 4235
box -3 -3 3 3
use M3_M2  M3_M2_11550
timestamp 1745462530
transform 1 0 212 0 1 3975
box -3 -3 3 3
use M3_M2  M3_M2_11551
timestamp 1745462530
transform 1 0 484 0 1 4155
box -3 -3 3 3
use M3_M2  M3_M2_11552
timestamp 1745462530
transform 1 0 340 0 1 4155
box -3 -3 3 3
use M3_M2  M3_M2_11553
timestamp 1745462530
transform 1 0 964 0 1 3935
box -3 -3 3 3
use M3_M2  M3_M2_11554
timestamp 1745462530
transform 1 0 852 0 1 3935
box -3 -3 3 3
use M3_M2  M3_M2_11555
timestamp 1745462530
transform 1 0 596 0 1 3935
box -3 -3 3 3
use M3_M2  M3_M2_11556
timestamp 1745462530
transform 1 0 1076 0 1 3975
box -3 -3 3 3
use M3_M2  M3_M2_11557
timestamp 1745462530
transform 1 0 812 0 1 3975
box -3 -3 3 3
use M3_M2  M3_M2_11558
timestamp 1745462530
transform 1 0 804 0 1 4245
box -3 -3 3 3
use M3_M2  M3_M2_11559
timestamp 1745462530
transform 1 0 748 0 1 4245
box -3 -3 3 3
use M3_M2  M3_M2_11560
timestamp 1745462530
transform 1 0 460 0 1 3985
box -3 -3 3 3
use M3_M2  M3_M2_11561
timestamp 1745462530
transform 1 0 340 0 1 3985
box -3 -3 3 3
use M3_M2  M3_M2_11562
timestamp 1745462530
transform 1 0 828 0 1 3995
box -3 -3 3 3
use M3_M2  M3_M2_11563
timestamp 1745462530
transform 1 0 796 0 1 3995
box -3 -3 3 3
use M3_M2  M3_M2_11564
timestamp 1745462530
transform 1 0 4380 0 1 4095
box -3 -3 3 3
use M3_M2  M3_M2_11565
timestamp 1745462530
transform 1 0 4356 0 1 4215
box -3 -3 3 3
use M3_M2  M3_M2_11566
timestamp 1745462530
transform 1 0 4356 0 1 4015
box -3 -3 3 3
use M3_M2  M3_M2_11567
timestamp 1745462530
transform 1 0 260 0 1 4155
box -3 -3 3 3
use M3_M2  M3_M2_11568
timestamp 1745462530
transform 1 0 252 0 1 3995
box -3 -3 3 3
use M3_M2  M3_M2_11569
timestamp 1745462530
transform 1 0 196 0 1 4155
box -3 -3 3 3
use M3_M2  M3_M2_11570
timestamp 1745462530
transform 1 0 108 0 1 4005
box -3 -3 3 3
use M3_M2  M3_M2_11571
timestamp 1745462530
transform 1 0 156 0 1 4095
box -3 -3 3 3
use M3_M2  M3_M2_11572
timestamp 1745462530
transform 1 0 84 0 1 4095
box -3 -3 3 3
use M3_M2  M3_M2_11573
timestamp 1745462530
transform 1 0 164 0 1 4135
box -3 -3 3 3
use M3_M2  M3_M2_11574
timestamp 1745462530
transform 1 0 84 0 1 4135
box -3 -3 3 3
use M3_M2  M3_M2_11575
timestamp 1745462530
transform 1 0 140 0 1 4195
box -3 -3 3 3
use M3_M2  M3_M2_11576
timestamp 1745462530
transform 1 0 132 0 1 4115
box -3 -3 3 3
use M3_M2  M3_M2_11577
timestamp 1745462530
transform 1 0 84 0 1 4125
box -3 -3 3 3
use M3_M2  M3_M2_11578
timestamp 1745462530
transform 1 0 76 0 1 4195
box -3 -3 3 3
use M3_M2  M3_M2_11579
timestamp 1745462530
transform 1 0 540 0 1 3705
box -3 -3 3 3
use M3_M2  M3_M2_11580
timestamp 1745462530
transform 1 0 524 0 1 3825
box -3 -3 3 3
use M3_M2  M3_M2_11581
timestamp 1745462530
transform 1 0 452 0 1 3825
box -3 -3 3 3
use M3_M2  M3_M2_11582
timestamp 1745462530
transform 1 0 452 0 1 3705
box -3 -3 3 3
use M3_M2  M3_M2_11583
timestamp 1745462530
transform 1 0 292 0 1 3825
box -3 -3 3 3
use M3_M2  M3_M2_11584
timestamp 1745462530
transform 1 0 188 0 1 3825
box -3 -3 3 3
use M3_M2  M3_M2_11585
timestamp 1745462530
transform 1 0 2108 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_11586
timestamp 1745462530
transform 1 0 2036 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_11587
timestamp 1745462530
transform 1 0 2012 0 1 1675
box -3 -3 3 3
use M3_M2  M3_M2_11588
timestamp 1745462530
transform 1 0 1844 0 1 3135
box -3 -3 3 3
use M3_M2  M3_M2_11589
timestamp 1745462530
transform 1 0 892 0 1 3135
box -3 -3 3 3
use M3_M2  M3_M2_11590
timestamp 1745462530
transform 1 0 292 0 1 2125
box -3 -3 3 3
use M3_M2  M3_M2_11591
timestamp 1745462530
transform 1 0 292 0 1 1675
box -3 -3 3 3
use M3_M2  M3_M2_11592
timestamp 1745462530
transform 1 0 212 0 1 3135
box -3 -3 3 3
use M3_M2  M3_M2_11593
timestamp 1745462530
transform 1 0 212 0 1 2865
box -3 -3 3 3
use M3_M2  M3_M2_11594
timestamp 1745462530
transform 1 0 116 0 1 2865
box -3 -3 3 3
use M3_M2  M3_M2_11595
timestamp 1745462530
transform 1 0 116 0 1 2365
box -3 -3 3 3
use M3_M2  M3_M2_11596
timestamp 1745462530
transform 1 0 76 0 1 2365
box -3 -3 3 3
use M3_M2  M3_M2_11597
timestamp 1745462530
transform 1 0 76 0 1 2245
box -3 -3 3 3
use M3_M2  M3_M2_11598
timestamp 1745462530
transform 1 0 76 0 1 2125
box -3 -3 3 3
use M3_M2  M3_M2_11599
timestamp 1745462530
transform 1 0 652 0 1 3845
box -3 -3 3 3
use M3_M2  M3_M2_11600
timestamp 1745462530
transform 1 0 588 0 1 4225
box -3 -3 3 3
use M3_M2  M3_M2_11601
timestamp 1745462530
transform 1 0 556 0 1 3845
box -3 -3 3 3
use M3_M2  M3_M2_11602
timestamp 1745462530
transform 1 0 540 0 1 4225
box -3 -3 3 3
use M3_M2  M3_M2_11603
timestamp 1745462530
transform 1 0 468 0 1 4225
box -3 -3 3 3
use NAND2X1  NAND2X1_0
timestamp 1745462530
transform 1 0 2176 0 1 2570
box -8 -3 32 105
use NAND2X1  NAND2X1_1
timestamp 1745462530
transform 1 0 2312 0 1 2570
box -8 -3 32 105
use NAND2X1  NAND2X1_2
timestamp 1745462530
transform 1 0 264 0 -1 3570
box -8 -3 32 105
use NAND2X1  NAND2X1_3
timestamp 1745462530
transform 1 0 352 0 -1 3570
box -8 -3 32 105
use NAND2X1  NAND2X1_4
timestamp 1745462530
transform 1 0 1104 0 1 3770
box -8 -3 32 105
use NAND2X1  NAND2X1_5
timestamp 1745462530
transform 1 0 776 0 1 3170
box -8 -3 32 105
use NAND2X1  NAND2X1_6
timestamp 1745462530
transform 1 0 2432 0 -1 2370
box -8 -3 32 105
use NAND2X1  NAND2X1_7
timestamp 1745462530
transform 1 0 2440 0 1 2570
box -8 -3 32 105
use NAND2X1  NAND2X1_8
timestamp 1745462530
transform 1 0 2392 0 -1 2370
box -8 -3 32 105
use NAND2X1  NAND2X1_9
timestamp 1745462530
transform 1 0 2416 0 1 2170
box -8 -3 32 105
use NAND2X1  NAND2X1_10
timestamp 1745462530
transform 1 0 2384 0 1 2170
box -8 -3 32 105
use NAND2X1  NAND2X1_11
timestamp 1745462530
transform 1 0 2344 0 1 2170
box -8 -3 32 105
use NAND2X1  NAND2X1_12
timestamp 1745462530
transform 1 0 2088 0 -1 3770
box -8 -3 32 105
use NAND2X1  NAND2X1_13
timestamp 1745462530
transform 1 0 2296 0 -1 3970
box -8 -3 32 105
use NAND2X1  NAND2X1_14
timestamp 1745462530
transform 1 0 2064 0 1 3770
box -8 -3 32 105
use NAND2X1  NAND2X1_15
timestamp 1745462530
transform 1 0 2104 0 1 3970
box -8 -3 32 105
use NAND2X1  NAND2X1_16
timestamp 1745462530
transform 1 0 2504 0 1 3770
box -8 -3 32 105
use NAND2X1  NAND2X1_17
timestamp 1745462530
transform 1 0 2728 0 -1 3970
box -8 -3 32 105
use NAND2X1  NAND2X1_18
timestamp 1745462530
transform 1 0 2584 0 1 3770
box -8 -3 32 105
use NAND2X1  NAND2X1_19
timestamp 1745462530
transform 1 0 1920 0 -1 3770
box -8 -3 32 105
use NAND2X1  NAND2X1_20
timestamp 1745462530
transform 1 0 1832 0 -1 3770
box -8 -3 32 105
use NAND2X1  NAND2X1_21
timestamp 1745462530
transform 1 0 2992 0 -1 3970
box -8 -3 32 105
use NAND2X1  NAND2X1_22
timestamp 1745462530
transform 1 0 1824 0 1 2170
box -8 -3 32 105
use NAND2X1  NAND2X1_23
timestamp 1745462530
transform 1 0 1656 0 1 1570
box -8 -3 32 105
use NAND2X1  NAND2X1_24
timestamp 1745462530
transform 1 0 1752 0 -1 1770
box -8 -3 32 105
use NAND2X1  NAND2X1_25
timestamp 1745462530
transform 1 0 1832 0 -1 1770
box -8 -3 32 105
use NAND2X1  NAND2X1_26
timestamp 1745462530
transform 1 0 1248 0 -1 2170
box -8 -3 32 105
use NAND2X1  NAND2X1_27
timestamp 1745462530
transform 1 0 1448 0 -1 2170
box -8 -3 32 105
use NAND2X1  NAND2X1_28
timestamp 1745462530
transform 1 0 3272 0 1 570
box -8 -3 32 105
use NAND2X1  NAND2X1_29
timestamp 1745462530
transform 1 0 3304 0 1 570
box -8 -3 32 105
use NAND2X1  NAND2X1_30
timestamp 1745462530
transform 1 0 3232 0 1 570
box -8 -3 32 105
use NAND2X1  NAND2X1_31
timestamp 1745462530
transform 1 0 3200 0 1 570
box -8 -3 32 105
use NAND2X1  NAND2X1_32
timestamp 1745462530
transform 1 0 2616 0 1 570
box -8 -3 32 105
use NAND2X1  NAND2X1_33
timestamp 1745462530
transform 1 0 2576 0 1 570
box -8 -3 32 105
use NAND2X1  NAND2X1_34
timestamp 1745462530
transform 1 0 2656 0 -1 770
box -8 -3 32 105
use NAND2X1  NAND2X1_35
timestamp 1745462530
transform 1 0 2656 0 1 570
box -8 -3 32 105
use NAND2X1  NAND2X1_36
timestamp 1745462530
transform 1 0 2640 0 -1 2370
box -8 -3 32 105
use NAND2X1  NAND2X1_37
timestamp 1745462530
transform 1 0 2584 0 -1 2370
box -8 -3 32 105
use NAND2X1  NAND2X1_38
timestamp 1745462530
transform 1 0 3304 0 1 1370
box -8 -3 32 105
use NAND2X1  NAND2X1_39
timestamp 1745462530
transform 1 0 3344 0 1 1370
box -8 -3 32 105
use NAND2X1  NAND2X1_40
timestamp 1745462530
transform 1 0 3256 0 1 1370
box -8 -3 32 105
use NAND2X1  NAND2X1_41
timestamp 1745462530
transform 1 0 3280 0 -1 1370
box -8 -3 32 105
use NAND2X1  NAND2X1_42
timestamp 1745462530
transform 1 0 912 0 1 2370
box -8 -3 32 105
use NAND2X1  NAND2X1_43
timestamp 1745462530
transform 1 0 840 0 1 2370
box -8 -3 32 105
use NAND2X1  NAND2X1_44
timestamp 1745462530
transform 1 0 912 0 -1 2570
box -8 -3 32 105
use NAND2X1  NAND2X1_45
timestamp 1745462530
transform 1 0 864 0 1 2370
box -8 -3 32 105
use NAND2X1  NAND2X1_46
timestamp 1745462530
transform 1 0 1024 0 1 2370
box -8 -3 32 105
use NAND2X1  NAND2X1_47
timestamp 1745462530
transform 1 0 2128 0 -1 2370
box -8 -3 32 105
use NAND2X1  NAND2X1_48
timestamp 1745462530
transform 1 0 2088 0 -1 2370
box -8 -3 32 105
use NAND2X1  NAND2X1_49
timestamp 1745462530
transform 1 0 1576 0 1 570
box -8 -3 32 105
use NAND2X1  NAND2X1_50
timestamp 1745462530
transform 1 0 1512 0 1 570
box -8 -3 32 105
use NAND2X1  NAND2X1_51
timestamp 1745462530
transform 1 0 1544 0 1 570
box -8 -3 32 105
use NAND2X1  NAND2X1_52
timestamp 1745462530
transform 1 0 1576 0 -1 770
box -8 -3 32 105
use NAND2X1  NAND2X1_53
timestamp 1745462530
transform 1 0 928 0 -1 770
box -8 -3 32 105
use NAND2X1  NAND2X1_54
timestamp 1745462530
transform 1 0 816 0 1 570
box -8 -3 32 105
use NAND2X1  NAND2X1_55
timestamp 1745462530
transform 1 0 888 0 -1 770
box -8 -3 32 105
use NAND2X1  NAND2X1_56
timestamp 1745462530
transform 1 0 848 0 -1 770
box -8 -3 32 105
use NAND2X1  NAND2X1_57
timestamp 1745462530
transform 1 0 2232 0 -1 3170
box -8 -3 32 105
use NAND2X1  NAND2X1_58
timestamp 1745462530
transform 1 0 984 0 1 3170
box -8 -3 32 105
use NAND2X1  NAND2X1_59
timestamp 1745462530
transform 1 0 1272 0 -1 3170
box -8 -3 32 105
use NAND2X1  NAND2X1_60
timestamp 1745462530
transform 1 0 1096 0 -1 3370
box -8 -3 32 105
use NAND2X1  NAND2X1_61
timestamp 1745462530
transform 1 0 1304 0 1 2370
box -8 -3 32 105
use NAND2X1  NAND2X1_62
timestamp 1745462530
transform 1 0 1624 0 -1 3770
box -8 -3 32 105
use NAND2X1  NAND2X1_63
timestamp 1745462530
transform 1 0 1656 0 1 3570
box -8 -3 32 105
use NAND2X1  NAND2X1_64
timestamp 1745462530
transform 1 0 1624 0 1 3570
box -8 -3 32 105
use NAND2X1  NAND2X1_65
timestamp 1745462530
transform 1 0 1568 0 -1 3570
box -8 -3 32 105
use NAND2X1  NAND2X1_66
timestamp 1745462530
transform 1 0 1608 0 1 3170
box -8 -3 32 105
use NAND2X1  NAND2X1_67
timestamp 1745462530
transform 1 0 1656 0 -1 3170
box -8 -3 32 105
use NAND2X1  NAND2X1_68
timestamp 1745462530
transform 1 0 1584 0 1 3170
box -8 -3 32 105
use NAND2X1  NAND2X1_69
timestamp 1745462530
transform 1 0 1296 0 1 3770
box -8 -3 32 105
use NAND2X1  NAND2X1_70
timestamp 1745462530
transform 1 0 1176 0 1 3770
box -8 -3 32 105
use NAND2X1  NAND2X1_71
timestamp 1745462530
transform 1 0 1208 0 1 3770
box -8 -3 32 105
use NAND2X1  NAND2X1_72
timestamp 1745462530
transform 1 0 1272 0 1 3770
box -8 -3 32 105
use NAND2X1  NAND2X1_73
timestamp 1745462530
transform 1 0 1000 0 -1 4170
box -8 -3 32 105
use NAND2X1  NAND2X1_74
timestamp 1745462530
transform 1 0 848 0 1 3970
box -8 -3 32 105
use NAND2X1  NAND2X1_75
timestamp 1745462530
transform 1 0 152 0 -1 3970
box -8 -3 32 105
use NAND2X1  NAND2X1_76
timestamp 1745462530
transform 1 0 96 0 -1 4170
box -8 -3 32 105
use NAND2X1  NAND2X1_77
timestamp 1745462530
transform 1 0 120 0 1 4170
box -8 -3 32 105
use NAND2X1  NAND2X1_78
timestamp 1745462530
transform 1 0 784 0 -1 4170
box -8 -3 32 105
use NAND2X1  NAND2X1_79
timestamp 1745462530
transform 1 0 1040 0 -1 3970
box -8 -3 32 105
use NAND2X1  NAND2X1_80
timestamp 1745462530
transform 1 0 1160 0 1 3970
box -8 -3 32 105
use NAND2X1  NAND2X1_81
timestamp 1745462530
transform 1 0 1288 0 1 3970
box -8 -3 32 105
use NAND2X1  NAND2X1_82
timestamp 1745462530
transform 1 0 1144 0 -1 4170
box -8 -3 32 105
use NAND2X1  NAND2X1_83
timestamp 1745462530
transform 1 0 1200 0 -1 4170
box -8 -3 32 105
use NAND2X1  NAND2X1_84
timestamp 1745462530
transform 1 0 1168 0 -1 4170
box -8 -3 32 105
use NAND2X1  NAND2X1_85
timestamp 1745462530
transform 1 0 1224 0 -1 4170
box -8 -3 32 105
use NAND2X1  NAND2X1_86
timestamp 1745462530
transform 1 0 464 0 -1 3970
box -8 -3 32 105
use NAND3X1  NAND3X1_0
timestamp 1745462530
transform 1 0 2256 0 -1 2770
box -8 -3 40 105
use NAND3X1  NAND3X1_1
timestamp 1745462530
transform 1 0 384 0 -1 3570
box -8 -3 40 105
use NAND3X1  NAND3X1_2
timestamp 1745462530
transform 1 0 1176 0 1 2970
box -8 -3 40 105
use NAND3X1  NAND3X1_3
timestamp 1745462530
transform 1 0 1696 0 1 2970
box -8 -3 40 105
use NAND3X1  NAND3X1_4
timestamp 1745462530
transform 1 0 1848 0 -1 3570
box -8 -3 40 105
use NAND3X1  NAND3X1_5
timestamp 1745462530
transform 1 0 2472 0 1 2970
box -8 -3 40 105
use NAND3X1  NAND3X1_6
timestamp 1745462530
transform 1 0 2264 0 1 3370
box -8 -3 40 105
use NAND3X1  NAND3X1_7
timestamp 1745462530
transform 1 0 1816 0 1 3570
box -8 -3 40 105
use NAND3X1  NAND3X1_8
timestamp 1745462530
transform 1 0 2360 0 1 2970
box -8 -3 40 105
use NAND3X1  NAND3X1_9
timestamp 1745462530
transform 1 0 2216 0 1 3370
box -8 -3 40 105
use NAND3X1  NAND3X1_10
timestamp 1745462530
transform 1 0 1728 0 1 3570
box -8 -3 40 105
use NAND3X1  NAND3X1_11
timestamp 1745462530
transform 1 0 2672 0 -1 3170
box -8 -3 40 105
use NAND3X1  NAND3X1_12
timestamp 1745462530
transform 1 0 2120 0 -1 3570
box -8 -3 40 105
use NAND3X1  NAND3X1_13
timestamp 1745462530
transform 1 0 1768 0 -1 3570
box -8 -3 40 105
use NAND3X1  NAND3X1_14
timestamp 1745462530
transform 1 0 2568 0 1 2970
box -8 -3 40 105
use NAND3X1  NAND3X1_15
timestamp 1745462530
transform 1 0 2144 0 1 3370
box -8 -3 40 105
use NAND3X1  NAND3X1_16
timestamp 1745462530
transform 1 0 1832 0 1 3370
box -8 -3 40 105
use NAND3X1  NAND3X1_17
timestamp 1745462530
transform 1 0 2720 0 1 2970
box -8 -3 40 105
use NAND3X1  NAND3X1_18
timestamp 1745462530
transform 1 0 2064 0 -1 3370
box -8 -3 40 105
use NAND3X1  NAND3X1_19
timestamp 1745462530
transform 1 0 1792 0 1 3370
box -8 -3 40 105
use NAND3X1  NAND3X1_20
timestamp 1745462530
transform 1 0 2752 0 1 2970
box -8 -3 40 105
use NAND3X1  NAND3X1_21
timestamp 1745462530
transform 1 0 2224 0 -1 3370
box -8 -3 40 105
use NAND3X1  NAND3X1_22
timestamp 1745462530
transform 1 0 1664 0 -1 3370
box -8 -3 40 105
use NAND3X1  NAND3X1_23
timestamp 1745462530
transform 1 0 2976 0 -1 3170
box -8 -3 40 105
use NAND3X1  NAND3X1_24
timestamp 1745462530
transform 1 0 3016 0 -1 3370
box -8 -3 40 105
use NAND3X1  NAND3X1_25
timestamp 1745462530
transform 1 0 1768 0 1 3170
box -8 -3 40 105
use NAND3X1  NAND3X1_26
timestamp 1745462530
transform 1 0 3032 0 1 2970
box -8 -3 40 105
use NAND3X1  NAND3X1_27
timestamp 1745462530
transform 1 0 3152 0 1 3170
box -8 -3 40 105
use NAND3X1  NAND3X1_28
timestamp 1745462530
transform 1 0 1704 0 -1 3370
box -8 -3 40 105
use NAND3X1  NAND3X1_29
timestamp 1745462530
transform 1 0 3064 0 -1 3170
box -8 -3 40 105
use NAND3X1  NAND3X1_30
timestamp 1745462530
transform 1 0 3128 0 -1 3370
box -8 -3 40 105
use NAND3X1  NAND3X1_31
timestamp 1745462530
transform 1 0 1688 0 1 3170
box -8 -3 40 105
use NAND3X1  NAND3X1_32
timestamp 1745462530
transform 1 0 3000 0 1 2970
box -8 -3 40 105
use NAND3X1  NAND3X1_33
timestamp 1745462530
transform 1 0 3096 0 1 3170
box -8 -3 40 105
use NAND3X1  NAND3X1_34
timestamp 1745462530
transform 1 0 1624 0 -1 3370
box -8 -3 40 105
use NAND3X1  NAND3X1_35
timestamp 1745462530
transform 1 0 3024 0 -1 3170
box -8 -3 40 105
use NAND3X1  NAND3X1_36
timestamp 1745462530
transform 1 0 3064 0 1 3170
box -8 -3 40 105
use NAND3X1  NAND3X1_37
timestamp 1745462530
transform 1 0 1648 0 1 3170
box -8 -3 40 105
use NAND3X1  NAND3X1_38
timestamp 1745462530
transform 1 0 2832 0 1 2970
box -8 -3 40 105
use NAND3X1  NAND3X1_39
timestamp 1745462530
transform 1 0 2928 0 1 3170
box -8 -3 40 105
use NAND3X1  NAND3X1_40
timestamp 1745462530
transform 1 0 1728 0 1 3170
box -8 -3 40 105
use NAND3X1  NAND3X1_41
timestamp 1745462530
transform 1 0 1696 0 -1 3570
box -8 -3 40 105
use NAND3X1  NAND3X1_42
timestamp 1745462530
transform 1 0 2608 0 1 2970
box -8 -3 40 105
use NAND3X1  NAND3X1_43
timestamp 1745462530
transform 1 0 2888 0 1 2970
box -8 -3 40 105
use NAND3X1  NAND3X1_44
timestamp 1745462530
transform 1 0 2992 0 1 3170
box -8 -3 40 105
use NAND3X1  NAND3X1_45
timestamp 1745462530
transform 1 0 2328 0 -1 3370
box -8 -3 40 105
use NAND3X1  NAND3X1_46
timestamp 1745462530
transform 1 0 1728 0 1 3370
box -8 -3 40 105
use NAND3X1  NAND3X1_47
timestamp 1745462530
transform 1 0 1656 0 1 3370
box -8 -3 40 105
use NAND3X1  NAND3X1_48
timestamp 1745462530
transform 1 0 2904 0 -1 3170
box -8 -3 40 105
use NAND3X1  NAND3X1_49
timestamp 1745462530
transform 1 0 2600 0 -1 3170
box -8 -3 40 105
use NAND3X1  NAND3X1_50
timestamp 1745462530
transform 1 0 2272 0 -1 3370
box -8 -3 40 105
use NAND3X1  NAND3X1_51
timestamp 1745462530
transform 1 0 2312 0 1 3170
box -8 -3 40 105
use NAND3X1  NAND3X1_52
timestamp 1745462530
transform 1 0 2192 0 1 3770
box -8 -3 40 105
use NAND3X1  NAND3X1_53
timestamp 1745462530
transform 1 0 2312 0 1 3770
box -8 -3 40 105
use NAND3X1  NAND3X1_54
timestamp 1745462530
transform 1 0 3432 0 1 3770
box -8 -3 40 105
use NAND3X1  NAND3X1_55
timestamp 1745462530
transform 1 0 3552 0 -1 3770
box -8 -3 40 105
use NAND3X1  NAND3X1_56
timestamp 1745462530
transform 1 0 1680 0 -1 3170
box -8 -3 40 105
use NAND3X1  NAND3X1_57
timestamp 1745462530
transform 1 0 2704 0 1 3770
box -8 -3 40 105
use NAND3X1  NAND3X1_58
timestamp 1745462530
transform 1 0 3504 0 -1 3970
box -8 -3 40 105
use NAND3X1  NAND3X1_59
timestamp 1745462530
transform 1 0 3568 0 1 3770
box -8 -3 40 105
use NAND3X1  NAND3X1_60
timestamp 1745462530
transform 1 0 1656 0 -1 3770
box -8 -3 40 105
use NAND3X1  NAND3X1_61
timestamp 1745462530
transform 1 0 1688 0 1 3570
box -8 -3 40 105
use NAND3X1  NAND3X1_62
timestamp 1745462530
transform 1 0 1776 0 1 2170
box -8 -3 40 105
use NAND3X1  NAND3X1_63
timestamp 1745462530
transform 1 0 3856 0 1 970
box -8 -3 40 105
use NAND3X1  NAND3X1_64
timestamp 1745462530
transform 1 0 2976 0 1 970
box -8 -3 40 105
use NAND3X1  NAND3X1_65
timestamp 1745462530
transform 1 0 3984 0 -1 2770
box -8 -3 40 105
use NAND3X1  NAND3X1_66
timestamp 1745462530
transform 1 0 3864 0 -1 2170
box -8 -3 40 105
use NAND3X1  NAND3X1_67
timestamp 1745462530
transform 1 0 656 0 1 2170
box -8 -3 40 105
use NAND3X1  NAND3X1_68
timestamp 1745462530
transform 1 0 1944 0 -1 2370
box -8 -3 40 105
use NAND3X1  NAND3X1_69
timestamp 1745462530
transform 1 0 1648 0 1 970
box -8 -3 40 105
use NAND3X1  NAND3X1_70
timestamp 1745462530
transform 1 0 664 0 1 970
box -8 -3 40 105
use NAND3X1  NAND3X1_71
timestamp 1745462530
transform 1 0 1488 0 1 1570
box -8 -3 40 105
use NAND3X1  NAND3X1_72
timestamp 1745462530
transform 1 0 3272 0 1 770
box -8 -3 40 105
use NAND3X1  NAND3X1_73
timestamp 1745462530
transform 1 0 3000 0 1 770
box -8 -3 40 105
use NAND3X1  NAND3X1_74
timestamp 1745462530
transform 1 0 3136 0 1 2570
box -8 -3 40 105
use NAND3X1  NAND3X1_75
timestamp 1745462530
transform 1 0 3072 0 -1 1770
box -8 -3 40 105
use NAND3X1  NAND3X1_76
timestamp 1745462530
transform 1 0 728 0 -1 2170
box -8 -3 40 105
use NAND3X1  NAND3X1_77
timestamp 1745462530
transform 1 0 1416 0 1 2370
box -8 -3 40 105
use NAND3X1  NAND3X1_78
timestamp 1745462530
transform 1 0 1472 0 -1 970
box -8 -3 40 105
use NAND3X1  NAND3X1_79
timestamp 1745462530
transform 1 0 680 0 1 770
box -8 -3 40 105
use NAND3X1  NAND3X1_80
timestamp 1745462530
transform 1 0 1712 0 1 1570
box -8 -3 40 105
use NAND3X1  NAND3X1_81
timestamp 1745462530
transform 1 0 3856 0 -1 970
box -8 -3 40 105
use NAND3X1  NAND3X1_82
timestamp 1745462530
transform 1 0 2416 0 -1 970
box -8 -3 40 105
use NAND3X1  NAND3X1_83
timestamp 1745462530
transform 1 0 4032 0 1 2570
box -8 -3 40 105
use NAND3X1  NAND3X1_84
timestamp 1745462530
transform 1 0 3408 0 -1 1770
box -8 -3 40 105
use NAND3X1  NAND3X1_85
timestamp 1745462530
transform 1 0 680 0 -1 2170
box -8 -3 40 105
use NAND3X1  NAND3X1_86
timestamp 1745462530
transform 1 0 1592 0 1 2370
box -8 -3 40 105
use NAND3X1  NAND3X1_87
timestamp 1745462530
transform 1 0 1840 0 -1 970
box -8 -3 40 105
use NAND3X1  NAND3X1_88
timestamp 1745462530
transform 1 0 728 0 1 770
box -8 -3 40 105
use NAND3X1  NAND3X1_89
timestamp 1745462530
transform 1 0 1896 0 -1 1770
box -8 -3 40 105
use NAND3X1  NAND3X1_90
timestamp 1745462530
transform 1 0 3744 0 1 770
box -8 -3 40 105
use NAND3X1  NAND3X1_91
timestamp 1745462530
transform 1 0 2552 0 1 770
box -8 -3 40 105
use NAND3X1  NAND3X1_92
timestamp 1745462530
transform 1 0 3784 0 1 2570
box -8 -3 40 105
use NAND3X1  NAND3X1_93
timestamp 1745462530
transform 1 0 3752 0 1 1570
box -8 -3 40 105
use NAND3X1  NAND3X1_94
timestamp 1745462530
transform 1 0 832 0 -1 2170
box -8 -3 40 105
use NAND3X1  NAND3X1_95
timestamp 1745462530
transform 1 0 1848 0 1 2370
box -8 -3 40 105
use NAND3X1  NAND3X1_96
timestamp 1745462530
transform 1 0 1992 0 1 770
box -8 -3 40 105
use NAND3X1  NAND3X1_97
timestamp 1745462530
transform 1 0 848 0 1 770
box -8 -3 40 105
use NAND3X1  NAND3X1_98
timestamp 1745462530
transform 1 0 1104 0 1 2170
box -8 -3 40 105
use NAND3X1  NAND3X1_99
timestamp 1745462530
transform 1 0 3432 0 1 770
box -8 -3 40 105
use NAND3X1  NAND3X1_100
timestamp 1745462530
transform 1 0 2584 0 1 770
box -8 -3 40 105
use NAND3X1  NAND3X1_101
timestamp 1745462530
transform 1 0 3320 0 -1 2770
box -8 -3 40 105
use NAND3X1  NAND3X1_102
timestamp 1745462530
transform 1 0 3296 0 1 1970
box -8 -3 40 105
use NAND3X1  NAND3X1_103
timestamp 1745462530
transform 1 0 856 0 1 2170
box -8 -3 40 105
use NAND3X1  NAND3X1_104
timestamp 1745462530
transform 1 0 1088 0 1 2370
box -8 -3 40 105
use NAND3X1  NAND3X1_105
timestamp 1745462530
transform 1 0 1224 0 -1 1170
box -8 -3 40 105
use NAND3X1  NAND3X1_106
timestamp 1745462530
transform 1 0 808 0 1 970
box -8 -3 40 105
use NAND3X1  NAND3X1_107
timestamp 1745462530
transform 1 0 1488 0 -1 2170
box -8 -3 40 105
use NAND3X1  NAND3X1_108
timestamp 1745462530
transform 1 0 3576 0 1 770
box -8 -3 40 105
use NAND3X1  NAND3X1_109
timestamp 1745462530
transform 1 0 2840 0 -1 970
box -8 -3 40 105
use NAND3X1  NAND3X1_110
timestamp 1745462530
transform 1 0 2232 0 -1 2170
box -8 -3 40 105
use NAND3X1  NAND3X1_111
timestamp 1745462530
transform 1 0 3520 0 1 2570
box -8 -3 40 105
use NAND3X1  NAND3X1_112
timestamp 1745462530
transform 1 0 3504 0 1 1970
box -8 -3 40 105
use NAND3X1  NAND3X1_113
timestamp 1745462530
transform 1 0 2256 0 -1 2370
box -8 -3 40 105
use NAND3X1  NAND3X1_114
timestamp 1745462530
transform 1 0 2280 0 -1 2170
box -8 -3 40 105
use NAND3X1  NAND3X1_115
timestamp 1745462530
transform 1 0 752 0 1 2170
box -8 -3 40 105
use NAND3X1  NAND3X1_116
timestamp 1745462530
transform 1 0 1472 0 1 2370
box -8 -3 40 105
use NAND3X1  NAND3X1_117
timestamp 1745462530
transform 1 0 2152 0 1 2170
box -8 -3 40 105
use NAND3X1  NAND3X1_118
timestamp 1745462530
transform 1 0 1160 0 -1 970
box -8 -3 40 105
use NAND3X1  NAND3X1_119
timestamp 1745462530
transform 1 0 2184 0 -1 2170
box -8 -3 40 105
use NAND3X1  NAND3X1_120
timestamp 1745462530
transform 1 0 736 0 -1 970
box -8 -3 40 105
use NAND3X1  NAND3X1_121
timestamp 1745462530
transform 1 0 2360 0 1 2370
box -8 -3 40 105
use NAND3X1  NAND3X1_122
timestamp 1745462530
transform 1 0 2304 0 1 2370
box -8 -3 40 105
use NAND3X1  NAND3X1_123
timestamp 1745462530
transform 1 0 2256 0 -1 2570
box -8 -3 40 105
use NAND3X1  NAND3X1_124
timestamp 1745462530
transform 1 0 2272 0 1 2170
box -8 -3 40 105
use NAND3X1  NAND3X1_125
timestamp 1745462530
transform 1 0 2296 0 -1 2370
box -8 -3 40 105
use NAND3X1  NAND3X1_126
timestamp 1745462530
transform 1 0 2088 0 -1 2170
box -8 -3 40 105
use NAND3X1  NAND3X1_127
timestamp 1745462530
transform 1 0 2352 0 -1 2370
box -8 -3 40 105
use NAND3X1  NAND3X1_128
timestamp 1745462530
transform 1 0 2136 0 -1 2170
box -8 -3 40 105
use NAND3X1  NAND3X1_129
timestamp 1745462530
transform 1 0 2304 0 -1 2570
box -8 -3 40 105
use NAND3X1  NAND3X1_130
timestamp 1745462530
transform 1 0 1088 0 1 3170
box -8 -3 40 105
use NAND3X1  NAND3X1_131
timestamp 1745462530
transform 1 0 2160 0 -1 2370
box -8 -3 40 105
use NAND3X1  NAND3X1_132
timestamp 1745462530
transform 1 0 2256 0 1 2370
box -8 -3 40 105
use NAND3X1  NAND3X1_133
timestamp 1745462530
transform 1 0 1584 0 1 2970
box -8 -3 40 105
use NAND3X1  NAND3X1_134
timestamp 1745462530
transform 1 0 1056 0 1 3370
box -8 -3 40 105
use NAND3X1  NAND3X1_135
timestamp 1745462530
transform 1 0 1032 0 -1 3570
box -8 -3 40 105
use NAND3X1  NAND3X1_136
timestamp 1745462530
transform 1 0 1544 0 1 3570
box -8 -3 40 105
use NAND3X1  NAND3X1_137
timestamp 1745462530
transform 1 0 1584 0 1 3570
box -8 -3 40 105
use NAND3X1  NAND3X1_138
timestamp 1745462530
transform 1 0 1496 0 -1 3370
box -8 -3 40 105
use NAND3X1  NAND3X1_139
timestamp 1745462530
transform 1 0 1424 0 1 3370
box -8 -3 40 105
use NAND3X1  NAND3X1_140
timestamp 1745462530
transform 1 0 1536 0 -1 3370
box -8 -3 40 105
use NAND3X1  NAND3X1_141
timestamp 1745462530
transform 1 0 1520 0 1 3170
box -8 -3 40 105
use NAND3X1  NAND3X1_142
timestamp 1745462530
transform 1 0 712 0 -1 4170
box -8 -3 40 105
use NAND3X1  NAND3X1_143
timestamp 1745462530
transform 1 0 928 0 -1 4170
box -8 -3 40 105
use NAND3X1  NAND3X1_144
timestamp 1745462530
transform 1 0 304 0 1 3970
box -8 -3 40 105
use NAND3X1  NAND3X1_145
timestamp 1745462530
transform 1 0 688 0 1 3970
box -8 -3 40 105
use NAND3X1  NAND3X1_146
timestamp 1745462530
transform 1 0 608 0 -1 4170
box -8 -3 40 105
use NAND3X1  NAND3X1_147
timestamp 1745462530
transform 1 0 216 0 1 3970
box -8 -3 40 105
use NAND3X1  NAND3X1_148
timestamp 1745462530
transform 1 0 120 0 -1 4170
box -8 -3 40 105
use NAND3X1  NAND3X1_149
timestamp 1745462530
transform 1 0 80 0 1 3970
box -8 -3 40 105
use NAND3X1  NAND3X1_150
timestamp 1745462530
transform 1 0 184 0 1 4170
box -8 -3 40 105
use NAND3X1  NAND3X1_151
timestamp 1745462530
transform 1 0 1072 0 1 3970
box -8 -3 40 105
use NAND3X1  NAND3X1_152
timestamp 1745462530
transform 1 0 1072 0 -1 4170
box -8 -3 40 105
use NOR2X1  NOR2X1_0
timestamp 1745462530
transform 1 0 2184 0 -1 2570
box -8 -3 32 105
use NOR2X1  NOR2X1_1
timestamp 1745462530
transform 1 0 2272 0 1 2570
box -8 -3 32 105
use NOR2X1  NOR2X1_2
timestamp 1745462530
transform 1 0 2224 0 -1 2770
box -8 -3 32 105
use NOR2X1  NOR2X1_3
timestamp 1745462530
transform 1 0 2296 0 -1 2770
box -8 -3 32 105
use NOR2X1  NOR2X1_4
timestamp 1745462530
transform 1 0 1792 0 1 2970
box -8 -3 32 105
use NOR2X1  NOR2X1_5
timestamp 1745462530
transform 1 0 872 0 1 3170
box -8 -3 32 105
use NOR2X1  NOR2X1_6
timestamp 1745462530
transform 1 0 3080 0 1 3570
box -8 -3 32 105
use NOR2X1  NOR2X1_7
timestamp 1745462530
transform 1 0 3384 0 -1 3770
box -8 -3 32 105
use NOR2X1  NOR2X1_8
timestamp 1745462530
transform 1 0 3264 0 -1 3770
box -8 -3 32 105
use NOR2X1  NOR2X1_9
timestamp 1745462530
transform 1 0 3320 0 1 3570
box -8 -3 32 105
use NOR2X1  NOR2X1_10
timestamp 1745462530
transform 1 0 3152 0 1 3570
box -8 -3 32 105
use NOR2X1  NOR2X1_11
timestamp 1745462530
transform 1 0 2376 0 1 3570
box -8 -3 32 105
use NOR2X1  NOR2X1_12
timestamp 1745462530
transform 1 0 2096 0 1 3570
box -8 -3 32 105
use NOR2X1  NOR2X1_13
timestamp 1745462530
transform 1 0 2856 0 1 3570
box -8 -3 32 105
use NOR2X1  NOR2X1_14
timestamp 1745462530
transform 1 0 3088 0 -1 3770
box -8 -3 32 105
use NOR2X1  NOR2X1_15
timestamp 1745462530
transform 1 0 3624 0 1 3570
box -8 -3 32 105
use NOR2X1  NOR2X1_16
timestamp 1745462530
transform 1 0 3456 0 1 3570
box -8 -3 32 105
use NOR2X1  NOR2X1_17
timestamp 1745462530
transform 1 0 3488 0 1 3570
box -8 -3 32 105
use NOR2X1  NOR2X1_18
timestamp 1745462530
transform 1 0 3184 0 1 3770
box -8 -3 32 105
use NOR2X1  NOR2X1_19
timestamp 1745462530
transform 1 0 2432 0 1 3770
box -8 -3 32 105
use NOR2X1  NOR2X1_20
timestamp 1745462530
transform 1 0 2320 0 -1 3770
box -8 -3 32 105
use NOR2X1  NOR2X1_21
timestamp 1745462530
transform 1 0 2448 0 1 2970
box -8 -3 32 105
use NOR2X1  NOR2X1_22
timestamp 1745462530
transform 1 0 2744 0 1 3570
box -8 -3 32 105
use NOR2X1  NOR2X1_23
timestamp 1745462530
transform 1 0 3016 0 -1 3770
box -8 -3 32 105
use NOR2X1  NOR2X1_24
timestamp 1745462530
transform 1 0 3320 0 -1 3770
box -8 -3 32 105
use NOR2X1  NOR2X1_25
timestamp 1745462530
transform 1 0 3288 0 -1 3770
box -8 -3 32 105
use NOR2X1  NOR2X1_26
timestamp 1745462530
transform 1 0 3208 0 1 3570
box -8 -3 32 105
use NOR2X1  NOR2X1_27
timestamp 1745462530
transform 1 0 3208 0 1 3770
box -8 -3 32 105
use NOR2X1  NOR2X1_28
timestamp 1745462530
transform 1 0 2400 0 1 3770
box -8 -3 32 105
use NOR2X1  NOR2X1_29
timestamp 1745462530
transform 1 0 2184 0 -1 3770
box -8 -3 32 105
use NOR2X1  NOR2X1_30
timestamp 1745462530
transform 1 0 2408 0 1 2970
box -8 -3 32 105
use NOR2X1  NOR2X1_31
timestamp 1745462530
transform 1 0 2184 0 1 3370
box -8 -3 32 105
use NOR2X1  NOR2X1_32
timestamp 1745462530
transform 1 0 2704 0 -1 3770
box -8 -3 32 105
use NOR2X1  NOR2X1_33
timestamp 1745462530
transform 1 0 2952 0 -1 3770
box -8 -3 32 105
use NOR2X1  NOR2X1_34
timestamp 1745462530
transform 1 0 3696 0 1 3570
box -8 -3 32 105
use NOR2X1  NOR2X1_35
timestamp 1745462530
transform 1 0 3760 0 -1 3770
box -8 -3 32 105
use NOR2X1  NOR2X1_36
timestamp 1745462530
transform 1 0 3712 0 -1 3570
box -8 -3 32 105
use NOR2X1  NOR2X1_37
timestamp 1745462530
transform 1 0 3688 0 -1 3770
box -8 -3 32 105
use NOR2X1  NOR2X1_38
timestamp 1745462530
transform 1 0 2504 0 -1 3770
box -8 -3 32 105
use NOR2X1  NOR2X1_39
timestamp 1745462530
transform 1 0 2288 0 1 3570
box -8 -3 32 105
use NOR2X1  NOR2X1_40
timestamp 1745462530
transform 1 0 2080 0 -1 3570
box -8 -3 32 105
use NOR2X1  NOR2X1_41
timestamp 1745462530
transform 1 0 2672 0 1 3570
box -8 -3 32 105
use NOR2X1  NOR2X1_42
timestamp 1745462530
transform 1 0 2928 0 1 3570
box -8 -3 32 105
use NOR2X1  NOR2X1_43
timestamp 1745462530
transform 1 0 3848 0 1 3570
box -8 -3 32 105
use NOR2X1  NOR2X1_44
timestamp 1745462530
transform 1 0 3872 0 1 3570
box -8 -3 32 105
use NOR2X1  NOR2X1_45
timestamp 1745462530
transform 1 0 3888 0 -1 3570
box -8 -3 32 105
use NOR2X1  NOR2X1_46
timestamp 1745462530
transform 1 0 3816 0 -1 3570
box -8 -3 32 105
use NOR2X1  NOR2X1_47
timestamp 1745462530
transform 1 0 1952 0 -1 3570
box -8 -3 32 105
use NOR2X1  NOR2X1_48
timestamp 1745462530
transform 1 0 2048 0 -1 3570
box -8 -3 32 105
use NOR2X1  NOR2X1_49
timestamp 1745462530
transform 1 0 1744 0 -1 3570
box -8 -3 32 105
use NOR2X1  NOR2X1_50
timestamp 1745462530
transform 1 0 2152 0 -1 3370
box -8 -3 32 105
use NOR2X1  NOR2X1_51
timestamp 1745462530
transform 1 0 2664 0 -1 3370
box -8 -3 32 105
use NOR2X1  NOR2X1_52
timestamp 1745462530
transform 1 0 2968 0 1 3370
box -8 -3 32 105
use NOR2X1  NOR2X1_53
timestamp 1745462530
transform 1 0 3872 0 -1 3370
box -8 -3 32 105
use NOR2X1  NOR2X1_54
timestamp 1745462530
transform 1 0 3896 0 1 3370
box -8 -3 32 105
use NOR2X1  NOR2X1_55
timestamp 1745462530
transform 1 0 3920 0 1 3370
box -8 -3 32 105
use NOR2X1  NOR2X1_56
timestamp 1745462530
transform 1 0 3768 0 1 3370
box -8 -3 32 105
use NOR2X1  NOR2X1_57
timestamp 1745462530
transform 1 0 2024 0 1 3370
box -8 -3 32 105
use NOR2X1  NOR2X1_58
timestamp 1745462530
transform 1 0 1928 0 1 3370
box -8 -3 32 105
use NOR2X1  NOR2X1_59
timestamp 1745462530
transform 1 0 1816 0 -1 3570
box -8 -3 32 105
use NOR2X1  NOR2X1_60
timestamp 1745462530
transform 1 0 2800 0 1 2970
box -8 -3 32 105
use NOR2X1  NOR2X1_61
timestamp 1745462530
transform 1 0 2024 0 -1 3370
box -8 -3 32 105
use NOR2X1  NOR2X1_62
timestamp 1745462530
transform 1 0 2016 0 1 3170
box -8 -3 32 105
use NOR2X1  NOR2X1_63
timestamp 1745462530
transform 1 0 1928 0 -1 3370
box -8 -3 32 105
use NOR2X1  NOR2X1_64
timestamp 1745462530
transform 1 0 3872 0 1 3170
box -8 -3 32 105
use NOR2X1  NOR2X1_65
timestamp 1745462530
transform 1 0 3848 0 -1 3370
box -8 -3 32 105
use NOR2X1  NOR2X1_66
timestamp 1745462530
transform 1 0 3896 0 1 3170
box -8 -3 32 105
use NOR2X1  NOR2X1_67
timestamp 1745462530
transform 1 0 3688 0 1 3170
box -8 -3 32 105
use NOR2X1  NOR2X1_68
timestamp 1745462530
transform 1 0 1864 0 1 3170
box -8 -3 32 105
use NOR2X1  NOR2X1_69
timestamp 1745462530
transform 1 0 1816 0 -1 3170
box -8 -3 32 105
use NOR2X1  NOR2X1_70
timestamp 1745462530
transform 1 0 2680 0 1 2970
box -8 -3 32 105
use NOR2X1  NOR2X1_71
timestamp 1745462530
transform 1 0 1752 0 -1 3370
box -8 -3 32 105
use NOR2X1  NOR2X1_72
timestamp 1745462530
transform 1 0 1896 0 -1 3370
box -8 -3 32 105
use NOR2X1  NOR2X1_73
timestamp 1745462530
transform 1 0 3760 0 -1 3170
box -8 -3 32 105
use NOR2X1  NOR2X1_74
timestamp 1745462530
transform 1 0 3712 0 1 3170
box -8 -3 32 105
use NOR2X1  NOR2X1_75
timestamp 1745462530
transform 1 0 3608 0 1 3170
box -8 -3 32 105
use NOR2X1  NOR2X1_76
timestamp 1745462530
transform 1 0 3248 0 1 3170
box -8 -3 32 105
use NOR2X1  NOR2X1_77
timestamp 1745462530
transform 1 0 2088 0 1 3170
box -8 -3 32 105
use NOR2X1  NOR2X1_78
timestamp 1745462530
transform 1 0 2816 0 1 3370
box -8 -3 32 105
use NOR2X1  NOR2X1_79
timestamp 1745462530
transform 1 0 1672 0 -1 3570
box -8 -3 32 105
use NOR2X1  NOR2X1_80
timestamp 1745462530
transform 1 0 2656 0 1 2970
box -8 -3 32 105
use NOR2X1  NOR2X1_81
timestamp 1745462530
transform 1 0 2120 0 -1 3370
box -8 -3 32 105
use NOR2X1  NOR2X1_82
timestamp 1745462530
transform 1 0 2232 0 1 3170
box -8 -3 32 105
use NOR2X1  NOR2X1_83
timestamp 1745462530
transform 1 0 1696 0 1 3370
box -8 -3 32 105
use NOR2X1  NOR2X1_84
timestamp 1745462530
transform 1 0 2528 0 -1 1770
box -8 -3 32 105
use NOR2X1  NOR2X1_85
timestamp 1745462530
transform 1 0 2080 0 1 970
box -8 -3 32 105
use NOR2X1  NOR2X1_86
timestamp 1745462530
transform 1 0 2096 0 1 1370
box -8 -3 32 105
use NOR2X1  NOR2X1_87
timestamp 1745462530
transform 1 0 816 0 -1 2370
box -8 -3 32 105
use NOR2X1  NOR2X1_88
timestamp 1745462530
transform 1 0 960 0 1 1770
box -8 -3 32 105
use NOR2X1  NOR2X1_89
timestamp 1745462530
transform 1 0 3720 0 -1 2570
box -8 -3 32 105
use NOR2X1  NOR2X1_90
timestamp 1745462530
transform 1 0 3768 0 -1 2370
box -8 -3 32 105
use NOR2X1  NOR2X1_91
timestamp 1745462530
transform 1 0 3704 0 -1 970
box -8 -3 32 105
use NOR2X1  NOR2X1_92
timestamp 1745462530
transform 1 0 3712 0 1 1170
box -8 -3 32 105
use NOR2X1  NOR2X1_93
timestamp 1745462530
transform 1 0 784 0 1 970
box -8 -3 32 105
use NOR2X1  NOR2X1_94
timestamp 1745462530
transform 1 0 1104 0 -1 1570
box -8 -3 32 105
use NOR2X1  NOR2X1_95
timestamp 1745462530
transform 1 0 1904 0 -1 2570
box -8 -3 32 105
use NOR2X1  NOR2X1_96
timestamp 1745462530
transform 1 0 1864 0 1 1770
box -8 -3 32 105
use NOR2X1  NOR2X1_97
timestamp 1745462530
transform 1 0 3136 0 1 1370
box -8 -3 32 105
use NOR2X1  NOR2X1_98
timestamp 1745462530
transform 1 0 2648 0 1 1570
box -8 -3 32 105
use NOR2X1  NOR2X1_99
timestamp 1745462530
transform 1 0 2480 0 -1 1170
box -8 -3 32 105
use NOR2X1  NOR2X1_100
timestamp 1745462530
transform 1 0 2464 0 -1 1370
box -8 -3 32 105
use NOR2X1  NOR2X1_101
timestamp 1745462530
transform 1 0 2560 0 -1 1770
box -8 -3 32 105
use NOR2X1  NOR2X1_102
timestamp 1745462530
transform 1 0 1064 0 1 970
box -8 -3 32 105
use NOR2X1  NOR2X1_103
timestamp 1745462530
transform 1 0 1152 0 -1 1570
box -8 -3 32 105
use NOR2X1  NOR2X1_104
timestamp 1745462530
transform 1 0 792 0 1 2370
box -8 -3 32 105
use NOR2X1  NOR2X1_105
timestamp 1745462530
transform 1 0 936 0 -1 1770
box -8 -3 32 105
use NOR2X1  NOR2X1_106
timestamp 1745462530
transform 1 0 3560 0 -1 2570
box -8 -3 32 105
use NOR2X1  NOR2X1_107
timestamp 1745462530
transform 1 0 3504 0 -1 2370
box -8 -3 32 105
use NOR2X1  NOR2X1_108
timestamp 1745462530
transform 1 0 3536 0 -1 970
box -8 -3 32 105
use NOR2X1  NOR2X1_109
timestamp 1745462530
transform 1 0 3504 0 1 1170
box -8 -3 32 105
use NOR2X1  NOR2X1_110
timestamp 1745462530
transform 1 0 928 0 1 1170
box -8 -3 32 105
use NOR2X1  NOR2X1_111
timestamp 1745462530
transform 1 0 1152 0 1 1370
box -8 -3 32 105
use NOR2X1  NOR2X1_112
timestamp 1745462530
transform 1 0 1416 0 1 2570
box -8 -3 32 105
use NOR2X1  NOR2X1_113
timestamp 1745462530
transform 1 0 1400 0 1 1570
box -8 -3 32 105
use NOR2X1  NOR2X1_114
timestamp 1745462530
transform 1 0 3248 0 -1 1970
box -8 -3 32 105
use NOR2X1  NOR2X1_115
timestamp 1745462530
transform 1 0 2776 0 1 1970
box -8 -3 32 105
use NOR2X1  NOR2X1_116
timestamp 1745462530
transform 1 0 2784 0 -1 1170
box -8 -3 32 105
use NOR2X1  NOR2X1_117
timestamp 1745462530
transform 1 0 2776 0 1 1370
box -8 -3 32 105
use NOR2X1  NOR2X1_118
timestamp 1745462530
transform 1 0 2440 0 -1 1970
box -8 -3 32 105
use NOR2X1  NOR2X1_119
timestamp 1745462530
transform 1 0 1144 0 -1 1170
box -8 -3 32 105
use NOR2X1  NOR2X1_120
timestamp 1745462530
transform 1 0 1192 0 1 1370
box -8 -3 32 105
use NOR2X1  NOR2X1_121
timestamp 1745462530
transform 1 0 888 0 1 1970
box -8 -3 32 105
use NOR2X1  NOR2X1_122
timestamp 1745462530
transform 1 0 1040 0 -1 1770
box -8 -3 32 105
use NOR2X1  NOR2X1_123
timestamp 1745462530
transform 1 0 3376 0 1 2570
box -8 -3 32 105
use NOR2X1  NOR2X1_124
timestamp 1745462530
transform 1 0 3296 0 1 2170
box -8 -3 32 105
use NOR2X1  NOR2X1_125
timestamp 1745462530
transform 1 0 3344 0 -1 1170
box -8 -3 32 105
use NOR2X1  NOR2X1_126
timestamp 1745462530
transform 1 0 3384 0 -1 1370
box -8 -3 32 105
use NOR2X1  NOR2X1_127
timestamp 1745462530
transform 1 0 936 0 -1 1170
box -8 -3 32 105
use NOR2X1  NOR2X1_128
timestamp 1745462530
transform 1 0 1200 0 -1 1370
box -8 -3 32 105
use NOR2X1  NOR2X1_129
timestamp 1745462530
transform 1 0 1112 0 1 2570
box -8 -3 32 105
use NOR2X1  NOR2X1_130
timestamp 1745462530
transform 1 0 1104 0 1 1770
box -8 -3 32 105
use NOR2X1  NOR2X1_131
timestamp 1745462530
transform 1 0 3080 0 -1 1970
box -8 -3 32 105
use NOR2X1  NOR2X1_132
timestamp 1745462530
transform 1 0 2512 0 1 1970
box -8 -3 32 105
use NOR2X1  NOR2X1_133
timestamp 1745462530
transform 1 0 2440 0 -1 1170
box -8 -3 32 105
use NOR2X1  NOR2X1_134
timestamp 1745462530
transform 1 0 2512 0 -1 1570
box -8 -3 32 105
use NOR2X1  NOR2X1_135
timestamp 1745462530
transform 1 0 2520 0 1 2970
box -8 -3 32 105
use NOR2X1  NOR2X1_136
timestamp 1745462530
transform 1 0 2344 0 -1 1970
box -8 -3 32 105
use NOR2X1  NOR2X1_137
timestamp 1745462530
transform 1 0 1656 0 -1 1170
box -8 -3 32 105
use NOR2X1  NOR2X1_138
timestamp 1745462530
transform 1 0 1720 0 -1 1570
box -8 -3 32 105
use NOR2X1  NOR2X1_139
timestamp 1745462530
transform 1 0 560 0 1 2170
box -8 -3 32 105
use NOR2X1  NOR2X1_140
timestamp 1745462530
transform 1 0 1032 0 -1 1970
box -8 -3 32 105
use NOR2X1  NOR2X1_141
timestamp 1745462530
transform 1 0 4080 0 -1 2570
box -8 -3 32 105
use NOR2X1  NOR2X1_142
timestamp 1745462530
transform 1 0 4072 0 -1 2370
box -8 -3 32 105
use NOR2X1  NOR2X1_143
timestamp 1745462530
transform 1 0 4040 0 -1 1170
box -8 -3 32 105
use NOR2X1  NOR2X1_144
timestamp 1745462530
transform 1 0 3976 0 -1 1370
box -8 -3 32 105
use NOR2X1  NOR2X1_145
timestamp 1745462530
transform 1 0 568 0 1 1170
box -8 -3 32 105
use NOR2X1  NOR2X1_146
timestamp 1745462530
transform 1 0 968 0 1 1370
box -8 -3 32 105
use NOR2X1  NOR2X1_147
timestamp 1745462530
transform 1 0 2080 0 1 2370
box -8 -3 32 105
use NOR2X1  NOR2X1_148
timestamp 1745462530
transform 1 0 2056 0 -1 1970
box -8 -3 32 105
use NOR2X1  NOR2X1_149
timestamp 1745462530
transform 1 0 3960 0 -1 2170
box -8 -3 32 105
use NOR2X1  NOR2X1_150
timestamp 1745462530
transform 1 0 3112 0 1 1970
box -8 -3 32 105
use NOR2X1  NOR2X1_151
timestamp 1745462530
transform 1 0 3168 0 -1 1170
box -8 -3 32 105
use NOR2X1  NOR2X1_152
timestamp 1745462530
transform 1 0 3152 0 -1 1370
box -8 -3 32 105
use NOR2X1  NOR2X1_153
timestamp 1745462530
transform 1 0 2256 0 -1 1770
box -8 -3 32 105
use NOR2X1  NOR2X1_154
timestamp 1745462530
transform 1 0 1776 0 -1 1170
box -8 -3 32 105
use NOR2X1  NOR2X1_155
timestamp 1745462530
transform 1 0 1840 0 -1 1570
box -8 -3 32 105
use NOR2X1  NOR2X1_156
timestamp 1745462530
transform 1 0 664 0 1 1970
box -8 -3 32 105
use NOR2X1  NOR2X1_157
timestamp 1745462530
transform 1 0 976 0 1 1570
box -8 -3 32 105
use NOR2X1  NOR2X1_158
timestamp 1745462530
transform 1 0 4048 0 1 2370
box -8 -3 32 105
use NOR2X1  NOR2X1_159
timestamp 1745462530
transform 1 0 4056 0 1 2170
box -8 -3 32 105
use NOR2X1  NOR2X1_160
timestamp 1745462530
transform 1 0 4064 0 -1 1170
box -8 -3 32 105
use NOR2X1  NOR2X1_161
timestamp 1745462530
transform 1 0 4016 0 -1 1370
box -8 -3 32 105
use NOR2X1  NOR2X1_162
timestamp 1745462530
transform 1 0 624 0 -1 1170
box -8 -3 32 105
use NOR2X1  NOR2X1_163
timestamp 1745462530
transform 1 0 1000 0 -1 1570
box -8 -3 32 105
use NOR2X1  NOR2X1_164
timestamp 1745462530
transform 1 0 1592 0 1 2570
box -8 -3 32 105
use NOR2X1  NOR2X1_165
timestamp 1745462530
transform 1 0 1576 0 -1 1770
box -8 -3 32 105
use NOR2X1  NOR2X1_166
timestamp 1745462530
transform 1 0 2944 0 -1 1570
box -8 -3 32 105
use NOR2X1  NOR2X1_167
timestamp 1745462530
transform 1 0 2600 0 1 1570
box -8 -3 32 105
use NOR2X1  NOR2X1_168
timestamp 1745462530
transform 1 0 2256 0 1 970
box -8 -3 32 105
use NOR2X1  NOR2X1_169
timestamp 1745462530
transform 1 0 2264 0 1 1370
box -8 -3 32 105
use NOR2X1  NOR2X1_170
timestamp 1745462530
transform 1 0 2392 0 -1 1770
box -8 -3 32 105
use NOR2X1  NOR2X1_171
timestamp 1745462530
transform 1 0 1504 0 -1 1170
box -8 -3 32 105
use NOR2X1  NOR2X1_172
timestamp 1745462530
transform 1 0 1448 0 -1 1570
box -8 -3 32 105
use NOR2X1  NOR2X1_173
timestamp 1745462530
transform 1 0 680 0 -1 2370
box -8 -3 32 105
use NOR2X1  NOR2X1_174
timestamp 1745462530
transform 1 0 1064 0 1 1770
box -8 -3 32 105
use NOR2X1  NOR2X1_175
timestamp 1745462530
transform 1 0 3128 0 -1 2570
box -8 -3 32 105
use NOR2X1  NOR2X1_176
timestamp 1745462530
transform 1 0 3144 0 1 1970
box -8 -3 32 105
use NOR2X1  NOR2X1_177
timestamp 1745462530
transform 1 0 3200 0 1 970
box -8 -3 32 105
use NOR2X1  NOR2X1_178
timestamp 1745462530
transform 1 0 3144 0 1 1170
box -8 -3 32 105
use NOR2X1  NOR2X1_179
timestamp 1745462530
transform 1 0 632 0 1 970
box -8 -3 32 105
use NOR2X1  NOR2X1_180
timestamp 1745462530
transform 1 0 1056 0 1 1370
box -8 -3 32 105
use NOR2X1  NOR2X1_181
timestamp 1745462530
transform 1 0 2160 0 1 1770
box -8 -3 32 105
use NOR2X1  NOR2X1_182
timestamp 1745462530
transform 1 0 1312 0 1 2570
box -8 -3 32 105
use NOR2X1  NOR2X1_183
timestamp 1745462530
transform 1 0 1256 0 1 1570
box -8 -3 32 105
use NOR2X1  NOR2X1_184
timestamp 1745462530
transform 1 0 2128 0 1 1770
box -8 -3 32 105
use NOR2X1  NOR2X1_185
timestamp 1745462530
transform 1 0 3104 0 1 1370
box -8 -3 32 105
use NOR2X1  NOR2X1_186
timestamp 1745462530
transform 1 0 2960 0 1 1570
box -8 -3 32 105
use NOR2X1  NOR2X1_187
timestamp 1745462530
transform 1 0 2184 0 -1 1970
box -8 -3 32 105
use NOR2X1  NOR2X1_188
timestamp 1745462530
transform 1 0 3040 0 -1 1170
box -8 -3 32 105
use NOR2X1  NOR2X1_189
timestamp 1745462530
transform 1 0 2400 0 1 2570
box -8 -3 32 105
use NOR2X1  NOR2X1_190
timestamp 1745462530
transform 1 0 3048 0 -1 1370
box -8 -3 32 105
use NOR2X1  NOR2X1_191
timestamp 1745462530
transform 1 0 2192 0 -1 1770
box -8 -3 32 105
use NOR2X1  NOR2X1_192
timestamp 1745462530
transform 1 0 2456 0 -1 2570
box -8 -3 32 105
use NOR2X1  NOR2X1_193
timestamp 1745462530
transform 1 0 2416 0 -1 2570
box -8 -3 32 105
use NOR2X1  NOR2X1_194
timestamp 1745462530
transform 1 0 2360 0 -1 2570
box -8 -3 32 105
use NOR2X1  NOR2X1_195
timestamp 1745462530
transform 1 0 2096 0 1 3370
box -8 -3 32 105
use NOR2X1  NOR2X1_196
timestamp 1745462530
transform 1 0 3936 0 1 3770
box -8 -3 32 105
use NOR2X1  NOR2X1_197
timestamp 1745462530
transform 1 0 1888 0 -1 3170
box -8 -3 32 105
use NOR2X1  NOR2X1_198
timestamp 1745462530
transform 1 0 4008 0 -1 3770
box -8 -3 32 105
use NOR2X1  NOR2X1_199
timestamp 1745462530
transform 1 0 1952 0 -1 3170
box -8 -3 32 105
use NOR2X1  NOR2X1_200
timestamp 1745462530
transform 1 0 4112 0 1 3770
box -8 -3 32 105
use NOR2X1  NOR2X1_201
timestamp 1745462530
transform 1 0 4192 0 -1 3770
box -8 -3 32 105
use NOR2X1  NOR2X1_202
timestamp 1745462530
transform 1 0 1976 0 -1 3170
box -8 -3 32 105
use NOR2X1  NOR2X1_203
timestamp 1745462530
transform 1 0 1912 0 -1 3170
box -8 -3 32 105
use NOR2X1  NOR2X1_204
timestamp 1745462530
transform 1 0 1880 0 -1 3770
box -8 -3 32 105
use NOR2X1  NOR2X1_205
timestamp 1745462530
transform 1 0 1784 0 -1 3770
box -8 -3 32 105
use NOR2X1  NOR2X1_206
timestamp 1745462530
transform 1 0 3728 0 1 970
box -8 -3 32 105
use NOR2X1  NOR2X1_207
timestamp 1745462530
transform 1 0 3856 0 -1 370
box -8 -3 32 105
use NOR2X1  NOR2X1_208
timestamp 1745462530
transform 1 0 2920 0 1 570
box -8 -3 32 105
use NOR2X1  NOR2X1_209
timestamp 1745462530
transform 1 0 3904 0 1 2170
box -8 -3 32 105
use NOR2X1  NOR2X1_210
timestamp 1745462530
transform 1 0 3872 0 -1 1970
box -8 -3 32 105
use NOR2X1  NOR2X1_211
timestamp 1745462530
transform 1 0 1752 0 1 2170
box -8 -3 32 105
use NOR2X1  NOR2X1_212
timestamp 1745462530
transform 1 0 648 0 1 2370
box -8 -3 32 105
use NOR2X1  NOR2X1_213
timestamp 1745462530
transform 1 0 1920 0 -1 2370
box -8 -3 32 105
use NOR2X1  NOR2X1_214
timestamp 1745462530
transform 1 0 1616 0 1 970
box -8 -3 32 105
use NOR2X1  NOR2X1_215
timestamp 1745462530
transform 1 0 1648 0 -1 770
box -8 -3 32 105
use NOR2X1  NOR2X1_216
timestamp 1745462530
transform 1 0 416 0 -1 970
box -8 -3 32 105
use NOR2X1  NOR2X1_217
timestamp 1745462530
transform 1 0 3144 0 1 770
box -8 -3 32 105
use NOR2X1  NOR2X1_218
timestamp 1745462530
transform 1 0 3312 0 -1 570
box -8 -3 32 105
use NOR2X1  NOR2X1_219
timestamp 1745462530
transform 1 0 2976 0 -1 770
box -8 -3 32 105
use NOR2X1  NOR2X1_220
timestamp 1745462530
transform 1 0 3040 0 -1 1770
box -8 -3 32 105
use NOR2X1  NOR2X1_221
timestamp 1745462530
transform 1 0 3368 0 1 1570
box -8 -3 32 105
use NOR2X1  NOR2X1_222
timestamp 1745462530
transform 1 0 1408 0 -1 2170
box -8 -3 32 105
use NOR2X1  NOR2X1_223
timestamp 1745462530
transform 1 0 696 0 1 2770
box -8 -3 32 105
use NOR2X1  NOR2X1_224
timestamp 1745462530
transform 1 0 1304 0 -1 2370
box -8 -3 32 105
use NOR2X1  NOR2X1_225
timestamp 1745462530
transform 1 0 1520 0 -1 970
box -8 -3 32 105
use NOR2X1  NOR2X1_226
timestamp 1745462530
transform 1 0 1472 0 1 570
box -8 -3 32 105
use NOR2X1  NOR2X1_227
timestamp 1745462530
transform 1 0 520 0 1 770
box -8 -3 32 105
use NOR2X1  NOR2X1_228
timestamp 1745462530
transform 1 0 3168 0 -1 970
box -8 -3 32 105
use NOR2X1  NOR2X1_229
timestamp 1745462530
transform 1 0 3856 0 1 370
box -8 -3 32 105
use NOR2X1  NOR2X1_230
timestamp 1745462530
transform 1 0 2432 0 1 570
box -8 -3 32 105
use NOR2X1  NOR2X1_231
timestamp 1745462530
transform 1 0 3448 0 -1 1770
box -8 -3 32 105
use NOR2X1  NOR2X1_232
timestamp 1745462530
transform 1 0 3544 0 -1 1570
box -8 -3 32 105
use NOR2X1  NOR2X1_233
timestamp 1745462530
transform 1 0 1608 0 1 2170
box -8 -3 32 105
use NOR2X1  NOR2X1_234
timestamp 1745462530
transform 1 0 680 0 1 2570
box -8 -3 32 105
use NOR2X1  NOR2X1_235
timestamp 1745462530
transform 1 0 1608 0 -1 2370
box -8 -3 32 105
use NOR2X1  NOR2X1_236
timestamp 1745462530
transform 1 0 1704 0 -1 970
box -8 -3 32 105
use NOR2X1  NOR2X1_237
timestamp 1745462530
transform 1 0 1856 0 1 570
box -8 -3 32 105
use NOR2X1  NOR2X1_238
timestamp 1745462530
transform 1 0 456 0 -1 770
box -8 -3 32 105
use NOR2X1  NOR2X1_239
timestamp 1745462530
transform 1 0 3544 0 1 770
box -8 -3 32 105
use NOR2X1  NOR2X1_240
timestamp 1745462530
transform 1 0 3672 0 1 570
box -8 -3 32 105
use NOR2X1  NOR2X1_241
timestamp 1745462530
transform 1 0 2568 0 -1 770
box -8 -3 32 105
use NOR2X1  NOR2X1_242
timestamp 1745462530
transform 1 0 3768 0 -1 1770
box -8 -3 32 105
use NOR2X1  NOR2X1_243
timestamp 1745462530
transform 1 0 3816 0 -1 1570
box -8 -3 32 105
use NOR2X1  NOR2X1_244
timestamp 1745462530
transform 1 0 1864 0 -1 2170
box -8 -3 32 105
use NOR2X1  NOR2X1_245
timestamp 1745462530
transform 1 0 824 0 1 2770
box -8 -3 32 105
use NOR2X1  NOR2X1_246
timestamp 1745462530
transform 1 0 1824 0 -1 2370
box -8 -3 32 105
use NOR2X1  NOR2X1_247
timestamp 1745462530
transform 1 0 1904 0 1 770
box -8 -3 32 105
use NOR2X1  NOR2X1_248
timestamp 1745462530
transform 1 0 2032 0 -1 570
box -8 -3 32 105
use NOR2X1  NOR2X1_249
timestamp 1745462530
transform 1 0 352 0 -1 770
box -8 -3 32 105
use NOR2X1  NOR2X1_250
timestamp 1745462530
transform 1 0 3240 0 1 770
box -8 -3 32 105
use NOR2X1  NOR2X1_251
timestamp 1745462530
transform 1 0 3464 0 1 570
box -8 -3 32 105
use NOR2X1  NOR2X1_252
timestamp 1745462530
transform 1 0 2464 0 1 570
box -8 -3 32 105
use NOR2X1  NOR2X1_253
timestamp 1745462530
transform 1 0 3248 0 -1 2170
box -8 -3 32 105
use NOR2X1  NOR2X1_254
timestamp 1745462530
transform 1 0 3464 0 -1 1970
box -8 -3 32 105
use NOR2X1  NOR2X1_255
timestamp 1745462530
transform 1 0 1072 0 1 2170
box -8 -3 32 105
use NOR2X1  NOR2X1_256
timestamp 1745462530
transform 1 0 888 0 1 2570
box -8 -3 32 105
use NOR2X1  NOR2X1_257
timestamp 1745462530
transform 1 0 1136 0 1 2370
box -8 -3 32 105
use NOR2X1  NOR2X1_258
timestamp 1745462530
transform 1 0 1176 0 -1 1170
box -8 -3 32 105
use NOR2X1  NOR2X1_259
timestamp 1745462530
transform 1 0 1200 0 1 570
box -8 -3 32 105
use NOR2X1  NOR2X1_260
timestamp 1745462530
transform 1 0 320 0 1 970
box -8 -3 32 105
use NOR2X1  NOR2X1_261
timestamp 1745462530
transform 1 0 3200 0 -1 970
box -8 -3 32 105
use NOR2X1  NOR2X1_262
timestamp 1745462530
transform 1 0 3616 0 1 370
box -8 -3 32 105
use NOR2X1  NOR2X1_263
timestamp 1745462530
transform 1 0 3208 0 -1 1170
box -8 -3 32 105
use NOR2X1  NOR2X1_264
timestamp 1745462530
transform 1 0 3240 0 -1 1170
box -8 -3 32 105
use NOR2X1  NOR2X1_265
timestamp 1745462530
transform 1 0 3208 0 -1 1370
box -8 -3 32 105
use NOR2X1  NOR2X1_266
timestamp 1745462530
transform 1 0 3184 0 1 1170
box -8 -3 32 105
use NOR2X1  NOR2X1_267
timestamp 1745462530
transform 1 0 2816 0 1 570
box -8 -3 32 105
use NOR2X1  NOR2X1_268
timestamp 1745462530
transform 1 0 2728 0 1 970
box -8 -3 32 105
use NOR2X1  NOR2X1_269
timestamp 1745462530
transform 1 0 2680 0 1 970
box -8 -3 32 105
use NOR2X1  NOR2X1_270
timestamp 1745462530
transform 1 0 2664 0 -1 1370
box -8 -3 32 105
use NOR2X1  NOR2X1_271
timestamp 1745462530
transform 1 0 2424 0 -1 1370
box -8 -3 32 105
use NOR2X1  NOR2X1_272
timestamp 1745462530
transform 1 0 3496 0 -1 2170
box -8 -3 32 105
use NOR2X1  NOR2X1_273
timestamp 1745462530
transform 1 0 2880 0 -1 2370
box -8 -3 32 105
use NOR2X1  NOR2X1_274
timestamp 1745462530
transform 1 0 2672 0 -1 2570
box -8 -3 32 105
use NOR2X1  NOR2X1_275
timestamp 1745462530
transform 1 0 2704 0 -1 2570
box -8 -3 32 105
use NOR2X1  NOR2X1_276
timestamp 1745462530
transform 1 0 2672 0 1 2370
box -8 -3 32 105
use NOR2X1  NOR2X1_277
timestamp 1745462530
transform 1 0 2624 0 1 2370
box -8 -3 32 105
use NOR2X1  NOR2X1_278
timestamp 1745462530
transform 1 0 3704 0 -1 1970
box -8 -3 32 105
use NOR2X1  NOR2X1_279
timestamp 1745462530
transform 1 0 3168 0 1 1770
box -8 -3 32 105
use NOR2X1  NOR2X1_280
timestamp 1745462530
transform 1 0 3208 0 1 1770
box -8 -3 32 105
use NOR2X1  NOR2X1_281
timestamp 1745462530
transform 1 0 2904 0 1 2370
box -8 -3 32 105
use NOR2X1  NOR2X1_282
timestamp 1745462530
transform 1 0 2952 0 -1 1970
box -8 -3 32 105
use NOR2X1  NOR2X1_283
timestamp 1745462530
transform 1 0 1488 0 1 2170
box -8 -3 32 105
use NOR2X1  NOR2X1_284
timestamp 1745462530
transform 1 0 672 0 -1 2770
box -8 -3 32 105
use NOR2X1  NOR2X1_285
timestamp 1745462530
transform 1 0 976 0 1 2170
box -8 -3 32 105
use NOR2X1  NOR2X1_286
timestamp 1745462530
transform 1 0 952 0 1 2170
box -8 -3 32 105
use NOR2X1  NOR2X1_287
timestamp 1745462530
transform 1 0 1088 0 -1 1970
box -8 -3 32 105
use NOR2X1  NOR2X1_288
timestamp 1745462530
transform 1 0 936 0 -1 2170
box -8 -3 32 105
use NOR2X1  NOR2X1_289
timestamp 1745462530
transform 1 0 1408 0 -1 2370
box -8 -3 32 105
use NOR2X1  NOR2X1_290
timestamp 1745462530
transform 1 0 2080 0 -1 2570
box -8 -3 32 105
use NOR2X1  NOR2X1_291
timestamp 1745462530
transform 1 0 2184 0 1 2370
box -8 -3 32 105
use NOR2X1  NOR2X1_292
timestamp 1745462530
transform 1 0 2136 0 1 2370
box -8 -3 32 105
use NOR2X1  NOR2X1_293
timestamp 1745462530
transform 1 0 1120 0 -1 970
box -8 -3 32 105
use NOR2X1  NOR2X1_294
timestamp 1745462530
transform 1 0 1168 0 1 570
box -8 -3 32 105
use NOR2X1  NOR2X1_295
timestamp 1745462530
transform 1 0 1392 0 -1 1170
box -8 -3 32 105
use NOR2X1  NOR2X1_296
timestamp 1745462530
transform 1 0 1584 0 1 970
box -8 -3 32 105
use NOR2X1  NOR2X1_297
timestamp 1745462530
transform 1 0 2280 0 1 1170
box -8 -3 32 105
use NOR2X1  NOR2X1_298
timestamp 1745462530
transform 1 0 1216 0 1 1170
box -8 -3 32 105
use NOR2X1  NOR2X1_299
timestamp 1745462530
transform 1 0 512 0 -1 970
box -8 -3 32 105
use NOR2X1  NOR2X1_300
timestamp 1745462530
transform 1 0 1024 0 -1 1170
box -8 -3 32 105
use NOR2X1  NOR2X1_301
timestamp 1745462530
transform 1 0 960 0 1 970
box -8 -3 32 105
use NOR2X1  NOR2X1_302
timestamp 1745462530
transform 1 0 1160 0 1 1170
box -8 -3 32 105
use NOR2X1  NOR2X1_303
timestamp 1745462530
transform 1 0 1112 0 1 1170
box -8 -3 32 105
use NOR2X1  NOR2X1_304
timestamp 1745462530
transform 1 0 2208 0 -1 2570
box -8 -3 32 105
use NOR2X1  NOR2X1_305
timestamp 1745462530
transform 1 0 1136 0 -1 3170
box -8 -3 32 105
use NOR2X1  NOR2X1_306
timestamp 1745462530
transform 1 0 2168 0 -1 3170
box -8 -3 32 105
use NOR2X1  NOR2X1_307
timestamp 1745462530
transform 1 0 504 0 1 3170
box -8 -3 32 105
use NOR2X1  NOR2X1_308
timestamp 1745462530
transform 1 0 1088 0 -1 3570
box -8 -3 32 105
use NOR2X1  NOR2X1_309
timestamp 1745462530
transform 1 0 1520 0 1 2970
box -8 -3 32 105
use NOR2X1  NOR2X1_310
timestamp 1745462530
transform 1 0 1472 0 -1 3770
box -8 -3 32 105
use NOR2X1  NOR2X1_311
timestamp 1745462530
transform 1 0 1536 0 -1 3570
box -8 -3 32 105
use NOR2X1  NOR2X1_312
timestamp 1745462530
transform 1 0 1336 0 1 3570
box -8 -3 32 105
use NOR2X1  NOR2X1_313
timestamp 1745462530
transform 1 0 624 0 1 4170
box -8 -3 32 105
use NOR2X1  NOR2X1_314
timestamp 1745462530
transform 1 0 688 0 -1 4170
box -8 -3 32 105
use NOR2X1  NOR2X1_315
timestamp 1745462530
transform 1 0 464 0 -1 4170
box -8 -3 32 105
use NOR2X1  NOR2X1_316
timestamp 1745462530
transform 1 0 544 0 -1 3970
box -8 -3 32 105
use NOR2X1  NOR2X1_317
timestamp 1745462530
transform 1 0 136 0 1 3970
box -8 -3 32 105
use NOR2X1  NOR2X1_318
timestamp 1745462530
transform 1 0 192 0 -1 4170
box -8 -3 32 105
use NOR2X1  NOR2X1_319
timestamp 1745462530
transform 1 0 152 0 -1 4170
box -8 -3 32 105
use NOR2X1  NOR2X1_320
timestamp 1745462530
transform 1 0 72 0 -1 4170
box -8 -3 32 105
use NOR2X1  NOR2X1_321
timestamp 1745462530
transform 1 0 1400 0 -1 4170
box -8 -3 32 105
use NOR2X1  NOR2X1_322
timestamp 1745462530
transform 1 0 1896 0 -1 4170
box -8 -3 32 105
use NOR2X1  NOR2X1_323
timestamp 1745462530
transform 1 0 1856 0 1 4170
box -8 -3 32 105
use NOR2X1  NOR2X1_324
timestamp 1745462530
transform 1 0 1488 0 1 4170
box -8 -3 32 105
use NOR2X1  NOR2X1_325
timestamp 1745462530
transform 1 0 1944 0 1 4170
box -8 -3 32 105
use NOR2X1  NOR2X1_326
timestamp 1745462530
transform 1 0 1968 0 1 4170
box -8 -3 32 105
use NOR2X1  NOR2X1_327
timestamp 1745462530
transform 1 0 4144 0 -1 4170
box -8 -3 32 105
use NOR2X1  NOR2X1_328
timestamp 1745462530
transform 1 0 3920 0 -1 4170
box -8 -3 32 105
use NOR2X1  NOR2X1_329
timestamp 1745462530
transform 1 0 3984 0 -1 4170
box -8 -3 32 105
use NOR2X1  NOR2X1_330
timestamp 1745462530
transform 1 0 4232 0 -1 3970
box -8 -3 32 105
use NOR2X1  NOR2X1_331
timestamp 1745462530
transform 1 0 4096 0 -1 3970
box -8 -3 32 105
use NOR2X1  NOR2X1_332
timestamp 1745462530
transform 1 0 4072 0 -1 3970
box -8 -3 32 105
use NOR2X1  NOR2X1_333
timestamp 1745462530
transform 1 0 4248 0 -1 4170
box -8 -3 32 105
use NOR2X1  NOR2X1_334
timestamp 1745462530
transform 1 0 4104 0 1 4170
box -8 -3 32 105
use NOR2X1  NOR2X1_335
timestamp 1745462530
transform 1 0 4096 0 1 3970
box -8 -3 32 105
use NOR2X1  NOR2X1_336
timestamp 1745462530
transform 1 0 4232 0 1 3970
box -8 -3 32 105
use NOR2X1  NOR2X1_337
timestamp 1745462530
transform 1 0 4120 0 1 3970
box -8 -3 32 105
use NOR2X1  NOR2X1_338
timestamp 1745462530
transform 1 0 4128 0 -1 3970
box -8 -3 32 105
use NOR2X1  NOR2X1_339
timestamp 1745462530
transform 1 0 1576 0 -1 4170
box -8 -3 32 105
use NOR2X1  NOR2X1_340
timestamp 1745462530
transform 1 0 2912 0 1 4170
box -8 -3 32 105
use NOR2X1  NOR2X1_341
timestamp 1745462530
transform 1 0 2936 0 1 4170
box -8 -3 32 105
use NOR2X1  NOR2X1_342
timestamp 1745462530
transform 1 0 1736 0 1 4170
box -8 -3 32 105
use NOR2X1  NOR2X1_343
timestamp 1745462530
transform 1 0 2616 0 1 4170
box -8 -3 32 105
use NOR2X1  NOR2X1_344
timestamp 1745462530
transform 1 0 2560 0 1 4170
box -8 -3 32 105
use NOR2X1  NOR2X1_345
timestamp 1745462530
transform 1 0 1128 0 1 3970
box -8 -3 32 105
use NOR2X1  NOR2X1_346
timestamp 1745462530
transform 1 0 1048 0 -1 4170
box -8 -3 32 105
use NOR2X1  NOR2X1_347
timestamp 1745462530
transform 1 0 1112 0 -1 4170
box -8 -3 32 105
use NOR2X1  NOR2X1_348
timestamp 1745462530
transform 1 0 768 0 -1 3970
box -8 -3 32 105
use NOR2X1  NOR2X1_349
timestamp 1745462530
transform 1 0 480 0 1 3970
box -8 -3 32 105
use NOR2X1  NOR2X1_350
timestamp 1745462530
transform 1 0 744 0 -1 3970
box -8 -3 32 105
use OAI21X1  OAI21X1_0
timestamp 1745462530
transform 1 0 2200 0 1 2570
box -8 -3 34 105
use OAI21X1  OAI21X1_1
timestamp 1745462530
transform 1 0 2240 0 1 2570
box -8 -3 34 105
use OAI21X1  OAI21X1_2
timestamp 1745462530
transform 1 0 320 0 -1 3570
box -8 -3 34 105
use OAI21X1  OAI21X1_3
timestamp 1745462530
transform 1 0 280 0 1 3570
box -8 -3 34 105
use OAI21X1  OAI21X1_4
timestamp 1745462530
transform 1 0 184 0 1 3570
box -8 -3 34 105
use OAI21X1  OAI21X1_5
timestamp 1745462530
transform 1 0 184 0 1 3370
box -8 -3 34 105
use OAI21X1  OAI21X1_6
timestamp 1745462530
transform 1 0 240 0 1 3370
box -8 -3 34 105
use OAI21X1  OAI21X1_7
timestamp 1745462530
transform 1 0 968 0 -1 3770
box -8 -3 34 105
use OAI21X1  OAI21X1_8
timestamp 1745462530
transform 1 0 1128 0 1 3770
box -8 -3 34 105
use OAI21X1  OAI21X1_9
timestamp 1745462530
transform 1 0 1208 0 1 2970
box -8 -3 34 105
use OAI21X1  OAI21X1_10
timestamp 1745462530
transform 1 0 800 0 1 3170
box -8 -3 34 105
use OAI21X1  OAI21X1_11
timestamp 1745462530
transform 1 0 2968 0 1 3570
box -8 -3 34 105
use OAI21X1  OAI21X1_12
timestamp 1745462530
transform 1 0 3072 0 1 3370
box -8 -3 34 105
use OAI21X1  OAI21X1_13
timestamp 1745462530
transform 1 0 3408 0 -1 3770
box -8 -3 34 105
use OAI21X1  OAI21X1_14
timestamp 1745462530
transform 1 0 3304 0 -1 3370
box -8 -3 34 105
use OAI21X1  OAI21X1_15
timestamp 1745462530
transform 1 0 3344 0 -1 3770
box -8 -3 34 105
use OAI21X1  OAI21X1_16
timestamp 1745462530
transform 1 0 3232 0 1 3370
box -8 -3 34 105
use OAI21X1  OAI21X1_17
timestamp 1745462530
transform 1 0 3344 0 1 3570
box -8 -3 34 105
use OAI21X1  OAI21X1_18
timestamp 1745462530
transform 1 0 3264 0 -1 3370
box -8 -3 34 105
use OAI21X1  OAI21X1_19
timestamp 1745462530
transform 1 0 3120 0 1 3570
box -8 -3 34 105
use OAI21X1  OAI21X1_20
timestamp 1745462530
transform 1 0 3152 0 1 3370
box -8 -3 34 105
use OAI21X1  OAI21X1_21
timestamp 1745462530
transform 1 0 2328 0 1 3570
box -8 -3 34 105
use OAI21X1  OAI21X1_22
timestamp 1745462530
transform 1 0 2392 0 1 3370
box -8 -3 34 105
use OAI21X1  OAI21X1_23
timestamp 1745462530
transform 1 0 2136 0 1 3570
box -8 -3 34 105
use OAI21X1  OAI21X1_24
timestamp 1745462530
transform 1 0 2352 0 1 3370
box -8 -3 34 105
use OAI21X1  OAI21X1_25
timestamp 1745462530
transform 1 0 2824 0 1 3570
box -8 -3 34 105
use OAI21X1  OAI21X1_26
timestamp 1745462530
transform 1 0 2832 0 -1 3570
box -8 -3 34 105
use OAI21X1  OAI21X1_27
timestamp 1745462530
transform 1 0 3056 0 -1 3770
box -8 -3 34 105
use OAI21X1  OAI21X1_28
timestamp 1745462530
transform 1 0 3048 0 1 3570
box -8 -3 34 105
use OAI21X1  OAI21X1_29
timestamp 1745462530
transform 1 0 3592 0 1 3570
box -8 -3 34 105
use OAI21X1  OAI21X1_30
timestamp 1745462530
transform 1 0 3416 0 -1 3570
box -8 -3 34 105
use OAI21X1  OAI21X1_31
timestamp 1745462530
transform 1 0 3424 0 1 3570
box -8 -3 34 105
use OAI21X1  OAI21X1_32
timestamp 1745462530
transform 1 0 3392 0 1 3570
box -8 -3 34 105
use OAI21X1  OAI21X1_33
timestamp 1745462530
transform 1 0 3512 0 1 3570
box -8 -3 34 105
use OAI21X1  OAI21X1_34
timestamp 1745462530
transform 1 0 3392 0 1 3370
box -8 -3 34 105
use OAI21X1  OAI21X1_35
timestamp 1745462530
transform 1 0 3120 0 -1 3770
box -8 -3 34 105
use OAI21X1  OAI21X1_36
timestamp 1745462530
transform 1 0 3136 0 -1 3570
box -8 -3 34 105
use OAI21X1  OAI21X1_37
timestamp 1745462530
transform 1 0 2408 0 -1 3770
box -8 -3 34 105
use OAI21X1  OAI21X1_38
timestamp 1745462530
transform 1 0 2504 0 1 3570
box -8 -3 34 105
use OAI21X1  OAI21X1_39
timestamp 1745462530
transform 1 0 2272 0 -1 3770
box -8 -3 34 105
use OAI21X1  OAI21X1_40
timestamp 1745462530
transform 1 0 2328 0 -1 3570
box -8 -3 34 105
use OAI21X1  OAI21X1_41
timestamp 1745462530
transform 1 0 2768 0 1 3570
box -8 -3 34 105
use OAI21X1  OAI21X1_42
timestamp 1745462530
transform 1 0 2744 0 -1 3570
box -8 -3 34 105
use OAI21X1  OAI21X1_43
timestamp 1745462530
transform 1 0 2984 0 -1 3770
box -8 -3 34 105
use OAI21X1  OAI21X1_44
timestamp 1745462530
transform 1 0 3000 0 1 3570
box -8 -3 34 105
use OAI21X1  OAI21X1_45
timestamp 1745462530
transform 1 0 3224 0 -1 3770
box -8 -3 34 105
use OAI21X1  OAI21X1_46
timestamp 1745462530
transform 1 0 3296 0 -1 3570
box -8 -3 34 105
use OAI21X1  OAI21X1_47
timestamp 1745462530
transform 1 0 3192 0 -1 3770
box -8 -3 34 105
use OAI21X1  OAI21X1_48
timestamp 1745462530
transform 1 0 3288 0 1 3570
box -8 -3 34 105
use OAI21X1  OAI21X1_49
timestamp 1745462530
transform 1 0 3176 0 1 3570
box -8 -3 34 105
use OAI21X1  OAI21X1_50
timestamp 1745462530
transform 1 0 3312 0 1 3370
box -8 -3 34 105
use OAI21X1  OAI21X1_51
timestamp 1745462530
transform 1 0 3152 0 -1 3770
box -8 -3 34 105
use OAI21X1  OAI21X1_52
timestamp 1745462530
transform 1 0 3216 0 -1 3570
box -8 -3 34 105
use OAI21X1  OAI21X1_53
timestamp 1745462530
transform 1 0 2352 0 -1 3770
box -8 -3 34 105
use OAI21X1  OAI21X1_54
timestamp 1745462530
transform 1 0 2408 0 1 3570
box -8 -3 34 105
use OAI21X1  OAI21X1_55
timestamp 1745462530
transform 1 0 2216 0 -1 3770
box -8 -3 34 105
use OAI21X1  OAI21X1_56
timestamp 1745462530
transform 1 0 2232 0 -1 3570
box -8 -3 34 105
use OAI21X1  OAI21X1_57
timestamp 1745462530
transform 1 0 2736 0 -1 3770
box -8 -3 34 105
use OAI21X1  OAI21X1_58
timestamp 1745462530
transform 1 0 2648 0 -1 3570
box -8 -3 34 105
use OAI21X1  OAI21X1_59
timestamp 1745462530
transform 1 0 2920 0 -1 3770
box -8 -3 34 105
use OAI21X1  OAI21X1_60
timestamp 1745462530
transform 1 0 2928 0 -1 3570
box -8 -3 34 105
use OAI21X1  OAI21X1_61
timestamp 1745462530
transform 1 0 3720 0 1 3570
box -8 -3 34 105
use OAI21X1  OAI21X1_62
timestamp 1745462530
transform 1 0 3672 0 -1 3570
box -8 -3 34 105
use OAI21X1  OAI21X1_63
timestamp 1745462530
transform 1 0 3728 0 -1 3770
box -8 -3 34 105
use OAI21X1  OAI21X1_64
timestamp 1745462530
transform 1 0 3656 0 1 3570
box -8 -3 34 105
use OAI21X1  OAI21X1_65
timestamp 1745462530
transform 1 0 3736 0 -1 3570
box -8 -3 34 105
use OAI21X1  OAI21X1_66
timestamp 1745462530
transform 1 0 3592 0 -1 3570
box -8 -3 34 105
use OAI21X1  OAI21X1_67
timestamp 1745462530
transform 1 0 3656 0 -1 3770
box -8 -3 34 105
use OAI21X1  OAI21X1_68
timestamp 1745462530
transform 1 0 3632 0 -1 3570
box -8 -3 34 105
use OAI21X1  OAI21X1_69
timestamp 1745462530
transform 1 0 2456 0 -1 3770
box -8 -3 34 105
use OAI21X1  OAI21X1_70
timestamp 1745462530
transform 1 0 2584 0 1 3570
box -8 -3 34 105
use OAI21X1  OAI21X1_71
timestamp 1745462530
transform 1 0 2248 0 1 3570
box -8 -3 34 105
use OAI21X1  OAI21X1_72
timestamp 1745462530
transform 1 0 2288 0 -1 3570
box -8 -3 34 105
use OAI21X1  OAI21X1_73
timestamp 1745462530
transform 1 0 2704 0 1 3570
box -8 -3 34 105
use OAI21X1  OAI21X1_74
timestamp 1745462530
transform 1 0 2680 0 1 3370
box -8 -3 34 105
use OAI21X1  OAI21X1_75
timestamp 1745462530
transform 1 0 2896 0 1 3570
box -8 -3 34 105
use OAI21X1  OAI21X1_76
timestamp 1745462530
transform 1 0 2928 0 1 3370
box -8 -3 34 105
use OAI21X1  OAI21X1_77
timestamp 1745462530
transform 1 0 3800 0 1 3570
box -8 -3 34 105
use OAI21X1  OAI21X1_78
timestamp 1745462530
transform 1 0 3664 0 1 3370
box -8 -3 34 105
use OAI21X1  OAI21X1_79
timestamp 1745462530
transform 1 0 3768 0 1 3570
box -8 -3 34 105
use OAI21X1  OAI21X1_80
timestamp 1745462530
transform 1 0 3696 0 1 3370
box -8 -3 34 105
use OAI21X1  OAI21X1_81
timestamp 1745462530
transform 1 0 3856 0 -1 3570
box -8 -3 34 105
use OAI21X1  OAI21X1_82
timestamp 1745462530
transform 1 0 3592 0 1 3370
box -8 -3 34 105
use OAI21X1  OAI21X1_83
timestamp 1745462530
transform 1 0 3784 0 -1 3570
box -8 -3 34 105
use OAI21X1  OAI21X1_84
timestamp 1745462530
transform 1 0 3624 0 1 3370
box -8 -3 34 105
use OAI21X1  OAI21X1_85
timestamp 1745462530
transform 1 0 1904 0 -1 3570
box -8 -3 34 105
use OAI21X1  OAI21X1_86
timestamp 1745462530
transform 1 0 2432 0 1 3370
box -8 -3 34 105
use OAI21X1  OAI21X1_87
timestamp 1745462530
transform 1 0 1992 0 -1 3570
box -8 -3 34 105
use OAI21X1  OAI21X1_88
timestamp 1745462530
transform 1 0 2312 0 1 3370
box -8 -3 34 105
use OAI21X1  OAI21X1_89
timestamp 1745462530
transform 1 0 2624 0 -1 3370
box -8 -3 34 105
use OAI21X1  OAI21X1_90
timestamp 1745462530
transform 1 0 2704 0 -1 3370
box -8 -3 34 105
use OAI21X1  OAI21X1_91
timestamp 1745462530
transform 1 0 2992 0 1 3370
box -8 -3 34 105
use OAI21X1  OAI21X1_92
timestamp 1745462530
transform 1 0 2968 0 -1 3370
box -8 -3 34 105
use OAI21X1  OAI21X1_93
timestamp 1745462530
transform 1 0 3768 0 -1 3370
box -8 -3 34 105
use OAI21X1  OAI21X1_94
timestamp 1745462530
transform 1 0 3616 0 -1 3370
box -8 -3 34 105
use OAI21X1  OAI21X1_95
timestamp 1745462530
transform 1 0 3808 0 1 3370
box -8 -3 34 105
use OAI21X1  OAI21X1_96
timestamp 1745462530
transform 1 0 3648 0 -1 3370
box -8 -3 34 105
use OAI21X1  OAI21X1_97
timestamp 1745462530
transform 1 0 3840 0 1 3370
box -8 -3 34 105
use OAI21X1  OAI21X1_98
timestamp 1745462530
transform 1 0 3536 0 -1 3370
box -8 -3 34 105
use OAI21X1  OAI21X1_99
timestamp 1745462530
transform 1 0 3736 0 1 3370
box -8 -3 34 105
use OAI21X1  OAI21X1_100
timestamp 1745462530
transform 1 0 3576 0 -1 3370
box -8 -3 34 105
use OAI21X1  OAI21X1_101
timestamp 1745462530
transform 1 0 1976 0 1 3370
box -8 -3 34 105
use OAI21X1  OAI21X1_102
timestamp 1745462530
transform 1 0 2440 0 -1 3370
box -8 -3 34 105
use OAI21X1  OAI21X1_103
timestamp 1745462530
transform 1 0 1888 0 1 3370
box -8 -3 34 105
use OAI21X1  OAI21X1_104
timestamp 1745462530
transform 1 0 2384 0 -1 3370
box -8 -3 34 105
use OAI21X1  OAI21X1_105
timestamp 1745462530
transform 1 0 1960 0 1 3170
box -8 -3 34 105
use OAI21X1  OAI21X1_106
timestamp 1745462530
transform 1 0 2656 0 1 3170
box -8 -3 34 105
use OAI21X1  OAI21X1_107
timestamp 1745462530
transform 1 0 1976 0 -1 3370
box -8 -3 34 105
use OAI21X1  OAI21X1_108
timestamp 1745462530
transform 1 0 2824 0 1 3170
box -8 -3 34 105
use OAI21X1  OAI21X1_109
timestamp 1745462530
transform 1 0 3784 0 1 3170
box -8 -3 34 105
use OAI21X1  OAI21X1_110
timestamp 1745462530
transform 1 0 3584 0 -1 3170
box -8 -3 34 105
use OAI21X1  OAI21X1_111
timestamp 1745462530
transform 1 0 3808 0 -1 3370
box -8 -3 34 105
use OAI21X1  OAI21X1_112
timestamp 1745462530
transform 1 0 3568 0 1 3170
box -8 -3 34 105
use OAI21X1  OAI21X1_113
timestamp 1745462530
transform 1 0 3824 0 1 3170
box -8 -3 34 105
use OAI21X1  OAI21X1_114
timestamp 1745462530
transform 1 0 3536 0 -1 3170
box -8 -3 34 105
use OAI21X1  OAI21X1_115
timestamp 1745462530
transform 1 0 3696 0 -1 3370
box -8 -3 34 105
use OAI21X1  OAI21X1_116
timestamp 1745462530
transform 1 0 3528 0 1 3170
box -8 -3 34 105
use OAI21X1  OAI21X1_117
timestamp 1745462530
transform 1 0 1912 0 1 3170
box -8 -3 34 105
use OAI21X1  OAI21X1_118
timestamp 1745462530
transform 1 0 2480 0 1 3170
box -8 -3 34 105
use OAI21X1  OAI21X1_119
timestamp 1745462530
transform 1 0 1816 0 1 3170
box -8 -3 34 105
use OAI21X1  OAI21X1_120
timestamp 1745462530
transform 1 0 2336 0 -1 3170
box -8 -3 34 105
use OAI21X1  OAI21X1_121
timestamp 1745462530
transform 1 0 1792 0 -1 3370
box -8 -3 34 105
use OAI21X1  OAI21X1_122
timestamp 1745462530
transform 1 0 2600 0 1 3170
box -8 -3 34 105
use OAI21X1  OAI21X1_123
timestamp 1745462530
transform 1 0 1848 0 -1 3370
box -8 -3 34 105
use OAI21X1  OAI21X1_124
timestamp 1745462530
transform 1 0 2816 0 -1 3370
box -8 -3 34 105
use OAI21X1  OAI21X1_125
timestamp 1745462530
transform 1 0 3744 0 1 3170
box -8 -3 34 105
use OAI21X1  OAI21X1_126
timestamp 1745462530
transform 1 0 3320 0 -1 3170
box -8 -3 34 105
use OAI21X1  OAI21X1_127
timestamp 1745462530
transform 1 0 3728 0 -1 3370
box -8 -3 34 105
use OAI21X1  OAI21X1_128
timestamp 1745462530
transform 1 0 3432 0 1 3170
box -8 -3 34 105
use OAI21X1  OAI21X1_129
timestamp 1745462530
transform 1 0 3640 0 1 3170
box -8 -3 34 105
use OAI21X1  OAI21X1_130
timestamp 1745462530
transform 1 0 3392 0 1 3170
box -8 -3 34 105
use OAI21X1  OAI21X1_131
timestamp 1745462530
transform 1 0 3080 0 -1 3370
box -8 -3 34 105
use OAI21X1  OAI21X1_132
timestamp 1745462530
transform 1 0 3216 0 1 3170
box -8 -3 34 105
use OAI21X1  OAI21X1_133
timestamp 1745462530
transform 1 0 2128 0 1 3170
box -8 -3 34 105
use OAI21X1  OAI21X1_134
timestamp 1745462530
transform 1 0 2360 0 1 3170
box -8 -3 34 105
use OAI21X1  OAI21X1_135
timestamp 1745462530
transform 1 0 2776 0 1 3370
box -8 -3 34 105
use OAI21X1  OAI21X1_136
timestamp 1745462530
transform 1 0 2840 0 1 3370
box -8 -3 34 105
use OAI21X1  OAI21X1_137
timestamp 1745462530
transform 1 0 2184 0 1 3170
box -8 -3 34 105
use OAI21X1  OAI21X1_138
timestamp 1745462530
transform 1 0 2272 0 -1 3170
box -8 -3 34 105
use OAI21X1  OAI21X1_139
timestamp 1745462530
transform 1 0 2040 0 1 770
box -8 -3 34 105
use OAI21X1  OAI21X1_140
timestamp 1745462530
transform 1 0 2080 0 -1 1370
box -8 -3 34 105
use OAI21X1  OAI21X1_141
timestamp 1745462530
transform 1 0 776 0 -1 2370
box -8 -3 34 105
use OAI21X1  OAI21X1_142
timestamp 1745462530
transform 1 0 912 0 1 1770
box -8 -3 34 105
use OAI21X1  OAI21X1_143
timestamp 1745462530
transform 1 0 3760 0 -1 2570
box -8 -3 34 105
use OAI21X1  OAI21X1_144
timestamp 1745462530
transform 1 0 3072 0 -1 2370
box -8 -3 34 105
use OAI21X1  OAI21X1_145
timestamp 1745462530
transform 1 0 3744 0 -1 770
box -8 -3 34 105
use OAI21X1  OAI21X1_146
timestamp 1745462530
transform 1 0 3664 0 1 1170
box -8 -3 34 105
use OAI21X1  OAI21X1_147
timestamp 1745462530
transform 1 0 800 0 -1 770
box -8 -3 34 105
use OAI21X1  OAI21X1_148
timestamp 1745462530
transform 1 0 1048 0 -1 1570
box -8 -3 34 105
use OAI21X1  OAI21X1_149
timestamp 1745462530
transform 1 0 1856 0 -1 2570
box -8 -3 34 105
use OAI21X1  OAI21X1_150
timestamp 1745462530
transform 1 0 1920 0 1 1770
box -8 -3 34 105
use OAI21X1  OAI21X1_151
timestamp 1745462530
transform 1 0 3704 0 -1 1570
box -8 -3 34 105
use OAI21X1  OAI21X1_152
timestamp 1745462530
transform 1 0 2656 0 -1 1770
box -8 -3 34 105
use OAI21X1  OAI21X1_153
timestamp 1745462530
transform 1 0 2520 0 -1 770
box -8 -3 34 105
use OAI21X1  OAI21X1_154
timestamp 1745462530
transform 1 0 2512 0 -1 1370
box -8 -3 34 105
use OAI21X1  OAI21X1_155
timestamp 1745462530
transform 1 0 1056 0 1 770
box -8 -3 34 105
use OAI21X1  OAI21X1_156
timestamp 1745462530
transform 1 0 1216 0 -1 1570
box -8 -3 34 105
use OAI21X1  OAI21X1_157
timestamp 1745462530
transform 1 0 760 0 -1 2570
box -8 -3 34 105
use OAI21X1  OAI21X1_158
timestamp 1745462530
transform 1 0 872 0 -1 1770
box -8 -3 34 105
use OAI21X1  OAI21X1_159
timestamp 1745462530
transform 1 0 3608 0 -1 2570
box -8 -3 34 105
use OAI21X1  OAI21X1_160
timestamp 1745462530
transform 1 0 3024 0 -1 2370
box -8 -3 34 105
use OAI21X1  OAI21X1_161
timestamp 1745462530
transform 1 0 3608 0 -1 770
box -8 -3 34 105
use OAI21X1  OAI21X1_162
timestamp 1745462530
transform 1 0 3536 0 1 1170
box -8 -3 34 105
use OAI21X1  OAI21X1_163
timestamp 1745462530
transform 1 0 784 0 -1 970
box -8 -3 34 105
use OAI21X1  OAI21X1_164
timestamp 1745462530
transform 1 0 1104 0 1 1370
box -8 -3 34 105
use OAI21X1  OAI21X1_165
timestamp 1745462530
transform 1 0 1472 0 -1 2770
box -8 -3 34 105
use OAI21X1  OAI21X1_166
timestamp 1745462530
transform 1 0 1336 0 1 1570
box -8 -3 34 105
use OAI21X1  OAI21X1_167
timestamp 1745462530
transform 1 0 3392 0 -1 1970
box -8 -3 34 105
use OAI21X1  OAI21X1_168
timestamp 1745462530
transform 1 0 2736 0 -1 2170
box -8 -3 34 105
use OAI21X1  OAI21X1_169
timestamp 1745462530
transform 1 0 2776 0 1 770
box -8 -3 34 105
use OAI21X1  OAI21X1_170
timestamp 1745462530
transform 1 0 2728 0 1 1370
box -8 -3 34 105
use OAI21X1  OAI21X1_171
timestamp 1745462530
transform 1 0 1072 0 -1 970
box -8 -3 34 105
use OAI21X1  OAI21X1_172
timestamp 1745462530
transform 1 0 1248 0 1 1370
box -8 -3 34 105
use OAI21X1  OAI21X1_173
timestamp 1745462530
transform 1 0 848 0 -1 2370
box -8 -3 34 105
use OAI21X1  OAI21X1_174
timestamp 1745462530
transform 1 0 984 0 -1 1770
box -8 -3 34 105
use OAI21X1  OAI21X1_175
timestamp 1745462530
transform 1 0 3424 0 1 2570
box -8 -3 34 105
use OAI21X1  OAI21X1_176
timestamp 1745462530
transform 1 0 2864 0 1 2170
box -8 -3 34 105
use OAI21X1  OAI21X1_177
timestamp 1745462530
transform 1 0 3376 0 1 770
box -8 -3 34 105
use OAI21X1  OAI21X1_178
timestamp 1745462530
transform 1 0 3336 0 -1 1370
box -8 -3 34 105
use OAI21X1  OAI21X1_179
timestamp 1745462530
transform 1 0 832 0 -1 970
box -8 -3 34 105
use OAI21X1  OAI21X1_180
timestamp 1745462530
transform 1 0 1152 0 -1 1370
box -8 -3 34 105
use OAI21X1  OAI21X1_181
timestamp 1745462530
transform 1 0 1168 0 -1 2770
box -8 -3 34 105
use OAI21X1  OAI21X1_182
timestamp 1745462530
transform 1 0 1152 0 1 1770
box -8 -3 34 105
use OAI21X1  OAI21X1_183
timestamp 1745462530
transform 1 0 3440 0 1 1970
box -8 -3 34 105
use OAI21X1  OAI21X1_184
timestamp 1745462530
transform 1 0 2536 0 -1 2170
box -8 -3 34 105
use OAI21X1  OAI21X1_185
timestamp 1745462530
transform 1 0 2448 0 1 770
box -8 -3 34 105
use OAI21X1  OAI21X1_186
timestamp 1745462530
transform 1 0 2448 0 -1 1570
box -8 -3 34 105
use OAI21X1  OAI21X1_187
timestamp 1745462530
transform 1 0 1624 0 1 770
box -8 -3 34 105
use OAI21X1  OAI21X1_188
timestamp 1745462530
transform 1 0 1712 0 1 1370
box -8 -3 34 105
use OAI21X1  OAI21X1_189
timestamp 1745462530
transform 1 0 536 0 -1 2370
box -8 -3 34 105
use OAI21X1  OAI21X1_190
timestamp 1745462530
transform 1 0 976 0 -1 1970
box -8 -3 34 105
use OAI21X1  OAI21X1_191
timestamp 1745462530
transform 1 0 4112 0 -1 2570
box -8 -3 34 105
use OAI21X1  OAI21X1_192
timestamp 1745462530
transform 1 0 2968 0 -1 2370
box -8 -3 34 105
use OAI21X1  OAI21X1_193
timestamp 1745462530
transform 1 0 3976 0 -1 970
box -8 -3 34 105
use OAI21X1  OAI21X1_194
timestamp 1745462530
transform 1 0 3864 0 -1 1370
box -8 -3 34 105
use OAI21X1  OAI21X1_195
timestamp 1745462530
transform 1 0 624 0 1 770
box -8 -3 34 105
use OAI21X1  OAI21X1_196
timestamp 1745462530
transform 1 0 920 0 1 1370
box -8 -3 34 105
use OAI21X1  OAI21X1_197
timestamp 1745462530
transform 1 0 2024 0 -1 2570
box -8 -3 34 105
use OAI21X1  OAI21X1_198
timestamp 1745462530
transform 1 0 2008 0 1 1770
box -8 -3 34 105
use OAI21X1  OAI21X1_199
timestamp 1745462530
transform 1 0 3992 0 -1 2170
box -8 -3 34 105
use OAI21X1  OAI21X1_200
timestamp 1745462530
transform 1 0 3056 0 1 1970
box -8 -3 34 105
use OAI21X1  OAI21X1_201
timestamp 1745462530
transform 1 0 3112 0 -1 970
box -8 -3 34 105
use OAI21X1  OAI21X1_202
timestamp 1745462530
transform 1 0 3096 0 -1 1370
box -8 -3 34 105
use OAI21X1  OAI21X1_203
timestamp 1745462530
transform 1 0 1768 0 1 770
box -8 -3 34 105
use OAI21X1  OAI21X1_204
timestamp 1745462530
transform 1 0 1888 0 -1 1570
box -8 -3 34 105
use OAI21X1  OAI21X1_205
timestamp 1745462530
transform 1 0 576 0 -1 2370
box -8 -3 34 105
use OAI21X1  OAI21X1_206
timestamp 1745462530
transform 1 0 912 0 1 1570
box -8 -3 34 105
use OAI21X1  OAI21X1_207
timestamp 1745462530
transform 1 0 4080 0 1 2370
box -8 -3 34 105
use OAI21X1  OAI21X1_208
timestamp 1745462530
transform 1 0 2920 0 -1 2370
box -8 -3 34 105
use OAI21X1  OAI21X1_209
timestamp 1745462530
transform 1 0 4032 0 -1 970
box -8 -3 34 105
use OAI21X1  OAI21X1_210
timestamp 1745462530
transform 1 0 3920 0 -1 1370
box -8 -3 34 105
use OAI21X1  OAI21X1_211
timestamp 1745462530
transform 1 0 568 0 -1 770
box -8 -3 34 105
use OAI21X1  OAI21X1_212
timestamp 1745462530
transform 1 0 944 0 -1 1570
box -8 -3 34 105
use OAI21X1  OAI21X1_213
timestamp 1745462530
transform 1 0 1616 0 -1 2770
box -8 -3 34 105
use OAI21X1  OAI21X1_214
timestamp 1745462530
transform 1 0 1512 0 -1 1770
box -8 -3 34 105
use OAI21X1  OAI21X1_215
timestamp 1745462530
transform 1 0 3232 0 -1 1570
box -8 -3 34 105
use OAI21X1  OAI21X1_216
timestamp 1745462530
transform 1 0 2600 0 -1 1770
box -8 -3 34 105
use OAI21X1  OAI21X1_217
timestamp 1745462530
transform 1 0 2248 0 1 770
box -8 -3 34 105
use OAI21X1  OAI21X1_218
timestamp 1745462530
transform 1 0 2320 0 1 1370
box -8 -3 34 105
use OAI21X1  OAI21X1_219
timestamp 1745462530
transform 1 0 1496 0 -1 770
box -8 -3 34 105
use OAI21X1  OAI21X1_220
timestamp 1745462530
transform 1 0 1504 0 -1 1570
box -8 -3 34 105
use OAI21X1  OAI21X1_221
timestamp 1745462530
transform 1 0 608 0 1 2370
box -8 -3 34 105
use OAI21X1  OAI21X1_222
timestamp 1745462530
transform 1 0 1016 0 1 1770
box -8 -3 34 105
use OAI21X1  OAI21X1_223
timestamp 1745462530
transform 1 0 3208 0 -1 2570
box -8 -3 34 105
use OAI21X1  OAI21X1_224
timestamp 1745462530
transform 1 0 2720 0 1 1970
box -8 -3 34 105
use OAI21X1  OAI21X1_225
timestamp 1745462530
transform 1 0 3280 0 -1 770
box -8 -3 34 105
use OAI21X1  OAI21X1_226
timestamp 1745462530
transform 1 0 3096 0 1 1170
box -8 -3 34 105
use OAI21X1  OAI21X1_227
timestamp 1745462530
transform 1 0 616 0 -1 770
box -8 -3 34 105
use OAI21X1  OAI21X1_228
timestamp 1745462530
transform 1 0 1016 0 1 1370
box -8 -3 34 105
use OAI21X1  OAI21X1_229
timestamp 1745462530
transform 1 0 1328 0 -1 2770
box -8 -3 34 105
use OAI21X1  OAI21X1_230
timestamp 1745462530
transform 1 0 1240 0 -1 1770
box -8 -3 34 105
use OAI21X1  OAI21X1_231
timestamp 1745462530
transform 1 0 3160 0 -1 1570
box -8 -3 34 105
use OAI21X1  OAI21X1_232
timestamp 1745462530
transform 1 0 2896 0 1 1570
box -8 -3 34 105
use OAI21X1  OAI21X1_233
timestamp 1745462530
transform 1 0 3008 0 -1 770
box -8 -3 34 105
use OAI21X1  OAI21X1_234
timestamp 1745462530
transform 1 0 3000 0 -1 1370
box -8 -3 34 105
use OAI21X1  OAI21X1_235
timestamp 1745462530
transform 1 0 2352 0 1 3770
box -8 -3 34 105
use OAI21X1  OAI21X1_236
timestamp 1745462530
transform 1 0 2264 0 1 3770
box -8 -3 34 105
use OAI21X1  OAI21X1_237
timestamp 1745462530
transform 1 0 2096 0 1 3770
box -8 -3 34 105
use OAI21X1  OAI21X1_238
timestamp 1745462530
transform 1 0 2664 0 1 3770
box -8 -3 34 105
use OAI21X1  OAI21X1_239
timestamp 1745462530
transform 1 0 2736 0 1 3770
box -8 -3 34 105
use OAI21X1  OAI21X1_240
timestamp 1745462530
transform 1 0 808 0 -1 3570
box -8 -3 34 105
use OAI21X1  OAI21X1_241
timestamp 1745462530
transform 1 0 848 0 -1 3570
box -8 -3 34 105
use OAI21X1  OAI21X1_242
timestamp 1745462530
transform 1 0 992 0 1 3570
box -8 -3 34 105
use OAI21X1  OAI21X1_243
timestamp 1745462530
transform 1 0 832 0 1 3370
box -8 -3 34 105
use OAI21X1  OAI21X1_244
timestamp 1745462530
transform 1 0 1248 0 1 3170
box -8 -3 34 105
use OAI21X1  OAI21X1_245
timestamp 1745462530
transform 1 0 1416 0 -1 3170
box -8 -3 34 105
use OAI21X1  OAI21X1_246
timestamp 1745462530
transform 1 0 1352 0 1 3170
box -8 -3 34 105
use OAI21X1  OAI21X1_247
timestamp 1745462530
transform 1 0 1024 0 1 3170
box -8 -3 34 105
use OAI21X1  OAI21X1_248
timestamp 1745462530
transform 1 0 1384 0 1 2170
box -8 -3 34 105
use OAI21X1  OAI21X1_249
timestamp 1745462530
transform 1 0 1376 0 -1 2570
box -8 -3 34 105
use OAI21X1  OAI21X1_250
timestamp 1745462530
transform 1 0 1440 0 1 2170
box -8 -3 34 105
use OAI21X1  OAI21X1_251
timestamp 1745462530
transform 1 0 992 0 -1 2570
box -8 -3 34 105
use OAI21X1  OAI21X1_252
timestamp 1745462530
transform 1 0 712 0 -1 2570
box -8 -3 34 105
use OAI21X1  OAI21X1_253
timestamp 1745462530
transform 1 0 512 0 -1 2570
box -8 -3 34 105
use OAI21X1  OAI21X1_254
timestamp 1745462530
transform 1 0 944 0 -1 2570
box -8 -3 34 105
use OAI21X1  OAI21X1_255
timestamp 1745462530
transform 1 0 448 0 1 2370
box -8 -3 34 105
use OAI21X1  OAI21X1_256
timestamp 1745462530
transform 1 0 432 0 1 770
box -8 -3 34 105
use OAI21X1  OAI21X1_257
timestamp 1745462530
transform 1 0 416 0 1 570
box -8 -3 34 105
use OAI21X1  OAI21X1_258
timestamp 1745462530
transform 1 0 408 0 -1 570
box -8 -3 34 105
use OAI21X1  OAI21X1_259
timestamp 1745462530
transform 1 0 512 0 -1 570
box -8 -3 34 105
use OAI21X1  OAI21X1_260
timestamp 1745462530
transform 1 0 1232 0 -1 570
box -8 -3 34 105
use OAI21X1  OAI21X1_261
timestamp 1745462530
transform 1 0 1288 0 -1 570
box -8 -3 34 105
use OAI21X1  OAI21X1_262
timestamp 1745462530
transform 1 0 1888 0 1 570
box -8 -3 34 105
use OAI21X1  OAI21X1_263
timestamp 1745462530
transform 1 0 1976 0 -1 570
box -8 -3 34 105
use OAI21X1  OAI21X1_264
timestamp 1745462530
transform 1 0 2600 0 -1 770
box -8 -3 34 105
use OAI21X1  OAI21X1_265
timestamp 1745462530
transform 1 0 2568 0 -1 570
box -8 -3 34 105
use OAI21X1  OAI21X1_266
timestamp 1745462530
transform 1 0 2608 0 -1 570
box -8 -3 34 105
use OAI21X1  OAI21X1_267
timestamp 1745462530
transform 1 0 2648 0 -1 570
box -8 -3 34 105
use OAI21X1  OAI21X1_268
timestamp 1745462530
transform 1 0 3504 0 -1 570
box -8 -3 34 105
use OAI21X1  OAI21X1_269
timestamp 1745462530
transform 1 0 3576 0 1 370
box -8 -3 34 105
use OAI21X1  OAI21X1_270
timestamp 1745462530
transform 1 0 3544 0 -1 570
box -8 -3 34 105
use OAI21X1  OAI21X1_271
timestamp 1745462530
transform 1 0 3792 0 -1 570
box -8 -3 34 105
use OAI21X1  OAI21X1_272
timestamp 1745462530
transform 1 0 3768 0 -1 1570
box -8 -3 34 105
use OAI21X1  OAI21X1_273
timestamp 1745462530
transform 1 0 4000 0 -1 1970
box -8 -3 34 105
use OAI21X1  OAI21X1_274
timestamp 1745462530
transform 1 0 3824 0 -1 1970
box -8 -3 34 105
use OAI21X1  OAI21X1_275
timestamp 1745462530
transform 1 0 3960 0 -1 1970
box -8 -3 34 105
use OAI21X1  OAI21X1_276
timestamp 1745462530
transform 1 0 3856 0 -1 2370
box -8 -3 34 105
use OAI21X1  OAI21X1_277
timestamp 1745462530
transform 1 0 3824 0 1 2370
box -8 -3 34 105
use OAI21X1  OAI21X1_278
timestamp 1745462530
transform 1 0 2304 0 1 2770
box -8 -3 34 105
use OAI21X1  OAI21X1_279
timestamp 1745462530
transform 1 0 2224 0 -1 2970
box -8 -3 34 105
use OAI21X1  OAI21X1_280
timestamp 1745462530
transform 1 0 2144 0 1 2770
box -8 -3 34 105
use OAI21X1  OAI21X1_281
timestamp 1745462530
transform 1 0 2048 0 1 2770
box -8 -3 34 105
use OAI21X1  OAI21X1_282
timestamp 1745462530
transform 1 0 2216 0 1 2970
box -8 -3 34 105
use OAI21X1  OAI21X1_283
timestamp 1745462530
transform 1 0 2096 0 1 2770
box -8 -3 34 105
use OAI21X1  OAI21X1_284
timestamp 1745462530
transform 1 0 696 0 1 3170
box -8 -3 34 105
use OAI21X1  OAI21X1_285
timestamp 1745462530
transform 1 0 648 0 1 3170
box -8 -3 34 105
use OAI21X1  OAI21X1_286
timestamp 1745462530
transform 1 0 912 0 1 3170
box -8 -3 34 105
use OAI21X1  OAI21X1_287
timestamp 1745462530
transform 1 0 1272 0 1 2970
box -8 -3 34 105
use OAI21X1  OAI21X1_288
timestamp 1745462530
transform 1 0 1424 0 -1 3770
box -8 -3 34 105
use OAI21X1  OAI21X1_289
timestamp 1745462530
transform 1 0 1376 0 1 3570
box -8 -3 34 105
use OAI21X1  OAI21X1_290
timestamp 1745462530
transform 1 0 1416 0 1 3570
box -8 -3 34 105
use OAI21X1  OAI21X1_291
timestamp 1745462530
transform 1 0 1328 0 -1 3770
box -8 -3 34 105
use OAI21X1  OAI21X1_292
timestamp 1745462530
transform 1 0 1368 0 -1 3570
box -8 -3 34 105
use OAI21X1  OAI21X1_293
timestamp 1745462530
transform 1 0 1408 0 -1 3370
box -8 -3 34 105
use OAI21X1  OAI21X1_294
timestamp 1745462530
transform 1 0 1384 0 1 3370
box -8 -3 34 105
use OAI21X1  OAI21X1_295
timestamp 1745462530
transform 1 0 576 0 1 4170
box -8 -3 34 105
use OAI21X1  OAI21X1_296
timestamp 1745462530
transform 1 0 752 0 -1 4170
box -8 -3 34 105
use OAI21X1  OAI21X1_297
timestamp 1745462530
transform 1 0 968 0 -1 4170
box -8 -3 34 105
use OAI21X1  OAI21X1_298
timestamp 1745462530
transform 1 0 1344 0 -1 4170
box -8 -3 34 105
use OAI21X1  OAI21X1_299
timestamp 1745462530
transform 1 0 896 0 -1 4170
box -8 -3 34 105
use OAI21X1  OAI21X1_300
timestamp 1745462530
transform 1 0 848 0 -1 4170
box -8 -3 34 105
use OAI21X1  OAI21X1_301
timestamp 1745462530
transform 1 0 424 0 1 3970
box -8 -3 34 105
use OAI21X1  OAI21X1_302
timestamp 1745462530
transform 1 0 336 0 1 3970
box -8 -3 34 105
use OAI21X1  OAI21X1_303
timestamp 1745462530
transform 1 0 264 0 1 3970
box -8 -3 34 105
use OAI21X1  OAI21X1_304
timestamp 1745462530
transform 1 0 504 0 1 3970
box -8 -3 34 105
use OAI21X1  OAI21X1_305
timestamp 1745462530
transform 1 0 560 0 1 3970
box -8 -3 34 105
use OAI21X1  OAI21X1_306
timestamp 1745462530
transform 1 0 648 0 1 3970
box -8 -3 34 105
use OAI21X1  OAI21X1_307
timestamp 1745462530
transform 1 0 584 0 -1 3970
box -8 -3 34 105
use OAI21X1  OAI21X1_308
timestamp 1745462530
transform 1 0 192 0 1 3770
box -8 -3 34 105
use OAI21X1  OAI21X1_309
timestamp 1745462530
transform 1 0 80 0 1 4170
box -8 -3 34 105
use OAI21X1  OAI21X1_310
timestamp 1745462530
transform 1 0 80 0 -1 3970
box -8 -3 34 105
use OAI21X1  OAI21X1_311
timestamp 1745462530
transform 1 0 1424 0 -1 4170
box -8 -3 34 105
use OAI21X1  OAI21X1_312
timestamp 1745462530
transform 1 0 1456 0 -1 4170
box -8 -3 34 105
use OAI21X1  OAI21X1_313
timestamp 1745462530
transform 1 0 1864 0 -1 4170
box -8 -3 34 105
use OAI21X1  OAI21X1_314
timestamp 1745462530
transform 1 0 1824 0 1 4170
box -8 -3 34 105
use OAI21X1  OAI21X1_315
timestamp 1745462530
transform 1 0 1488 0 -1 4170
box -8 -3 34 105
use OAI21X1  OAI21X1_316
timestamp 1745462530
transform 1 0 1512 0 1 4170
box -8 -3 34 105
use OAI21X1  OAI21X1_317
timestamp 1745462530
transform 1 0 1912 0 1 4170
box -8 -3 34 105
use OAI21X1  OAI21X1_318
timestamp 1745462530
transform 1 0 1992 0 1 4170
box -8 -3 34 105
use OAI21X1  OAI21X1_319
timestamp 1745462530
transform 1 0 4112 0 -1 4170
box -8 -3 34 105
use OAI21X1  OAI21X1_320
timestamp 1745462530
transform 1 0 4072 0 -1 4170
box -8 -3 34 105
use OAI21X1  OAI21X1_321
timestamp 1745462530
transform 1 0 3944 0 -1 4170
box -8 -3 34 105
use OAI21X1  OAI21X1_322
timestamp 1745462530
transform 1 0 4008 0 1 4170
box -8 -3 34 105
use OAI21X1  OAI21X1_323
timestamp 1745462530
transform 1 0 4200 0 -1 3970
box -8 -3 34 105
use OAI21X1  OAI21X1_324
timestamp 1745462530
transform 1 0 4160 0 -1 3970
box -8 -3 34 105
use OAI21X1  OAI21X1_325
timestamp 1745462530
transform 1 0 3952 0 1 3970
box -8 -3 34 105
use OAI21X1  OAI21X1_326
timestamp 1745462530
transform 1 0 3992 0 -1 3970
box -8 -3 34 105
use OAI21X1  OAI21X1_327
timestamp 1745462530
transform 1 0 4216 0 -1 4170
box -8 -3 34 105
use OAI21X1  OAI21X1_328
timestamp 1745462530
transform 1 0 4176 0 -1 4170
box -8 -3 34 105
use OAI21X1  OAI21X1_329
timestamp 1745462530
transform 1 0 4072 0 1 4170
box -8 -3 34 105
use OAI21X1  OAI21X1_330
timestamp 1745462530
transform 1 0 4040 0 1 4170
box -8 -3 34 105
use OAI21X1  OAI21X1_331
timestamp 1745462530
transform 1 0 4200 0 1 3970
box -8 -3 34 105
use OAI21X1  OAI21X1_332
timestamp 1745462530
transform 1 0 4160 0 1 3970
box -8 -3 34 105
use OAI21X1  OAI21X1_333
timestamp 1745462530
transform 1 0 4040 0 -1 4170
box -8 -3 34 105
use OAI21X1  OAI21X1_334
timestamp 1745462530
transform 1 0 4008 0 1 3970
box -8 -3 34 105
use OAI21X1  OAI21X1_335
timestamp 1745462530
transform 1 0 1544 0 -1 4170
box -8 -3 34 105
use OAI21X1  OAI21X1_336
timestamp 1745462530
transform 1 0 1760 0 1 4170
box -8 -3 34 105
use OAI21X1  OAI21X1_337
timestamp 1745462530
transform 1 0 2880 0 1 4170
box -8 -3 34 105
use OAI21X1  OAI21X1_338
timestamp 1745462530
transform 1 0 2960 0 1 4170
box -8 -3 34 105
use OAI21X1  OAI21X1_339
timestamp 1745462530
transform 1 0 1704 0 -1 4170
box -8 -3 34 105
use OAI21X1  OAI21X1_340
timestamp 1745462530
transform 1 0 1792 0 1 4170
box -8 -3 34 105
use OAI21X1  OAI21X1_341
timestamp 1745462530
transform 1 0 2640 0 1 4170
box -8 -3 34 105
use OAI21X1  OAI21X1_342
timestamp 1745462530
transform 1 0 2584 0 1 4170
box -8 -3 34 105
use OAI22X1  OAI22X1_0
timestamp 1745462530
transform 1 0 104 0 -1 3570
box -8 -3 46 105
use OAI22X1  OAI22X1_1
timestamp 1745462530
transform 1 0 3112 0 1 3770
box -8 -3 46 105
use OAI22X1  OAI22X1_2
timestamp 1745462530
transform 1 0 3360 0 -1 3970
box -8 -3 46 105
use OAI22X1  OAI22X1_3
timestamp 1745462530
transform 1 0 3288 0 -1 3970
box -8 -3 46 105
use OAI22X1  OAI22X1_4
timestamp 1745462530
transform 1 0 3344 0 1 3770
box -8 -3 46 105
use OAI22X1  OAI22X1_5
timestamp 1745462530
transform 1 0 3152 0 -1 3970
box -8 -3 46 105
use OAI22X1  OAI22X1_6
timestamp 1745462530
transform 1 0 2376 0 -1 3970
box -8 -3 46 105
use OAI22X1  OAI22X1_7
timestamp 1745462530
transform 1 0 2064 0 -1 3970
box -8 -3 46 105
use OAI22X1  OAI22X1_8
timestamp 1745462530
transform 1 0 2832 0 -1 3970
box -8 -3 46 105
use OAI22X1  OAI22X1_9
timestamp 1745462530
transform 1 0 3080 0 -1 3970
box -8 -3 46 105
use OAI22X1  OAI22X1_10
timestamp 1745462530
transform 1 0 3624 0 1 3770
box -8 -3 46 105
use OAI22X1  OAI22X1_11
timestamp 1745462530
transform 1 0 3592 0 -1 3970
box -8 -3 46 105
use OAI22X1  OAI22X1_12
timestamp 1745462530
transform 1 0 3584 0 -1 3770
box -8 -3 46 105
use OAI22X1  OAI22X1_13
timestamp 1745462530
transform 1 0 3224 0 -1 4170
box -8 -3 46 105
use OAI22X1  OAI22X1_14
timestamp 1745462530
transform 1 0 2368 0 1 3970
box -8 -3 46 105
use OAI22X1  OAI22X1_15
timestamp 1745462530
transform 1 0 2208 0 -1 3970
box -8 -3 46 105
use OAI22X1  OAI22X1_16
timestamp 1745462530
transform 1 0 2736 0 -1 4170
box -8 -3 46 105
use OAI22X1  OAI22X1_17
timestamp 1745462530
transform 1 0 3008 0 -1 4170
box -8 -3 46 105
use OAI22X1  OAI22X1_18
timestamp 1745462530
transform 1 0 3480 0 -1 4170
box -8 -3 46 105
use OAI22X1  OAI22X1_19
timestamp 1745462530
transform 1 0 3376 0 -1 4170
box -8 -3 46 105
use OAI22X1  OAI22X1_20
timestamp 1745462530
transform 1 0 3496 0 1 3970
box -8 -3 46 105
use OAI22X1  OAI22X1_21
timestamp 1745462530
transform 1 0 3168 0 -1 4170
box -8 -3 46 105
use OAI22X1  OAI22X1_22
timestamp 1745462530
transform 1 0 2400 0 -1 4170
box -8 -3 46 105
use OAI22X1  OAI22X1_23
timestamp 1745462530
transform 1 0 2168 0 -1 4170
box -8 -3 46 105
use OAI22X1  OAI22X1_24
timestamp 1745462530
transform 1 0 2640 0 -1 4170
box -8 -3 46 105
use OAI22X1  OAI22X1_25
timestamp 1745462530
transform 1 0 2976 0 1 3970
box -8 -3 46 105
use OAI22X1  OAI22X1_26
timestamp 1745462530
transform 1 0 3752 0 1 3970
box -8 -3 46 105
use OAI22X1  OAI22X1_27
timestamp 1745462530
transform 1 0 3848 0 -1 4170
box -8 -3 46 105
use OAI22X1  OAI22X1_28
timestamp 1745462530
transform 1 0 3680 0 -1 3970
box -8 -3 46 105
use OAI22X1  OAI22X1_29
timestamp 1745462530
transform 1 0 3704 0 -1 4170
box -8 -3 46 105
use OAI22X1  OAI22X1_30
timestamp 1745462530
transform 1 0 2480 0 -1 4170
box -8 -3 46 105
use OAI22X1  OAI22X1_31
timestamp 1745462530
transform 1 0 2280 0 -1 4170
box -8 -3 46 105
use OAI22X1  OAI22X1_32
timestamp 1745462530
transform 1 0 2584 0 1 3970
box -8 -3 46 105
use OAI22X1  OAI22X1_33
timestamp 1745462530
transform 1 0 2912 0 -1 3970
box -8 -3 46 105
use OAI22X1  OAI22X1_34
timestamp 1745462530
transform 1 0 4296 0 -1 3770
box -8 -3 46 105
use OAI22X1  OAI22X1_35
timestamp 1745462530
transform 1 0 4208 0 1 3770
box -8 -3 46 105
use OAI22X1  OAI22X1_36
timestamp 1745462530
transform 1 0 4224 0 1 3570
box -8 -3 46 105
use OAI22X1  OAI22X1_37
timestamp 1745462530
transform 1 0 3952 0 -1 3570
box -8 -3 46 105
use OAI22X1  OAI22X1_38
timestamp 1745462530
transform 1 0 1976 0 -1 3770
box -8 -3 46 105
use OAI22X1  OAI22X1_39
timestamp 1745462530
transform 1 0 2008 0 -1 3970
box -8 -3 46 105
use OAI22X1  OAI22X1_40
timestamp 1745462530
transform 1 0 2672 0 -1 3970
box -8 -3 46 105
use OAI22X1  OAI22X1_41
timestamp 1745462530
transform 1 0 2848 0 -1 3770
box -8 -3 46 105
use OAI22X1  OAI22X1_42
timestamp 1745462530
transform 1 0 4064 0 -1 3570
box -8 -3 46 105
use OAI22X1  OAI22X1_43
timestamp 1745462530
transform 1 0 4040 0 1 3570
box -8 -3 46 105
use OAI22X1  OAI22X1_44
timestamp 1745462530
transform 1 0 4128 0 1 3370
box -8 -3 46 105
use OAI22X1  OAI22X1_45
timestamp 1745462530
transform 1 0 3960 0 1 3370
box -8 -3 46 105
use OAI22X1  OAI22X1_46
timestamp 1745462530
transform 1 0 2008 0 1 3570
box -8 -3 46 105
use OAI22X1  OAI22X1_47
timestamp 1745462530
transform 1 0 1920 0 -1 3970
box -8 -3 46 105
use OAI22X1  OAI22X1_48
timestamp 1745462530
transform 1 0 1856 0 -1 3970
box -8 -3 46 105
use OAI22X1  OAI22X1_49
timestamp 1745462530
transform 1 0 1776 0 -1 3970
box -8 -3 46 105
use OAI22X1  OAI22X1_50
timestamp 1745462530
transform 1 0 4216 0 -1 3370
box -8 -3 46 105
use OAI22X1  OAI22X1_51
timestamp 1745462530
transform 1 0 4208 0 1 3370
box -8 -3 46 105
use OAI22X1  OAI22X1_52
timestamp 1745462530
transform 1 0 4024 0 1 3170
box -8 -3 46 105
use OAI22X1  OAI22X1_53
timestamp 1745462530
transform 1 0 3944 0 1 3170
box -8 -3 46 105
use OAI22X1  OAI22X1_54
timestamp 1745462530
transform 1 0 1656 0 1 3770
box -8 -3 46 105
use OAI22X1  OAI22X1_55
timestamp 1745462530
transform 1 0 1640 0 -1 3970
box -8 -3 46 105
use OAI22X1  OAI22X1_56
timestamp 1745462530
transform 1 0 1704 0 -1 3970
box -8 -3 46 105
use OAI22X1  OAI22X1_57
timestamp 1745462530
transform 1 0 1680 0 1 3970
box -8 -3 46 105
use OAI22X1  OAI22X1_58
timestamp 1745462530
transform 1 0 4200 0 -1 3170
box -8 -3 46 105
use OAI22X1  OAI22X1_59
timestamp 1745462530
transform 1 0 4208 0 1 3170
box -8 -3 46 105
use OAI22X1  OAI22X1_60
timestamp 1745462530
transform 1 0 4024 0 -1 3370
box -8 -3 46 105
use OAI22X1  OAI22X1_61
timestamp 1745462530
transform 1 0 3816 0 -1 3770
box -8 -3 46 105
use OAI22X1  OAI22X1_62
timestamp 1745462530
transform 1 0 1552 0 -1 3770
box -8 -3 46 105
use OAI22X1  OAI22X1_63
timestamp 1745462530
transform 1 0 2776 0 -1 3770
box -8 -3 46 105
use OAI22X1  OAI22X1_64
timestamp 1745462530
transform 1 0 1584 0 1 3770
box -8 -3 46 105
use OAI22X1  OAI22X1_65
timestamp 1745462530
transform 1 0 2120 0 1 970
box -8 -3 46 105
use OAI22X1  OAI22X1_66
timestamp 1745462530
transform 1 0 2088 0 1 770
box -8 -3 46 105
use OAI22X1  OAI22X1_67
timestamp 1745462530
transform 1 0 712 0 -1 2370
box -8 -3 46 105
use OAI22X1  OAI22X1_68
timestamp 1745462530
transform 1 0 928 0 1 1970
box -8 -3 46 105
use OAI22X1  OAI22X1_69
timestamp 1745462530
transform 1 0 3664 0 -1 2570
box -8 -3 46 105
use OAI22X1  OAI22X1_70
timestamp 1745462530
transform 1 0 3800 0 -1 2370
box -8 -3 46 105
use OAI22X1  OAI22X1_71
timestamp 1745462530
transform 1 0 3640 0 -1 970
box -8 -3 46 105
use OAI22X1  OAI22X1_72
timestamp 1745462530
transform 1 0 3800 0 1 770
box -8 -3 46 105
use OAI22X1  OAI22X1_73
timestamp 1745462530
transform 1 0 712 0 1 970
box -8 -3 46 105
use OAI22X1  OAI22X1_74
timestamp 1745462530
transform 1 0 1000 0 1 770
box -8 -3 46 105
use OAI22X1  OAI22X1_75
timestamp 1745462530
transform 1 0 1944 0 -1 2570
box -8 -3 46 105
use OAI22X1  OAI22X1_76
timestamp 1745462530
transform 1 0 1912 0 1 1970
box -8 -3 46 105
use OAI22X1  OAI22X1_77
timestamp 1745462530
transform 1 0 3192 0 1 1370
box -8 -3 46 105
use OAI22X1  OAI22X1_78
timestamp 1745462530
transform 1 0 3704 0 1 1570
box -8 -3 46 105
use OAI22X1  OAI22X1_79
timestamp 1745462530
transform 1 0 2496 0 1 970
box -8 -3 46 105
use OAI22X1  OAI22X1_80
timestamp 1745462530
transform 1 0 2384 0 1 770
box -8 -3 46 105
use OAI22X1  OAI22X1_81
timestamp 1745462530
transform 1 0 1008 0 1 970
box -8 -3 46 105
use OAI22X1  OAI22X1_82
timestamp 1745462530
transform 1 0 1112 0 1 770
box -8 -3 46 105
use OAI22X1  OAI22X1_83
timestamp 1745462530
transform 1 0 744 0 1 2370
box -8 -3 46 105
use OAI22X1  OAI22X1_84
timestamp 1745462530
transform 1 0 976 0 1 1970
box -8 -3 46 105
use OAI22X1  OAI22X1_85
timestamp 1745462530
transform 1 0 3496 0 -1 2570
box -8 -3 46 105
use OAI22X1  OAI22X1_86
timestamp 1745462530
transform 1 0 3544 0 -1 2370
box -8 -3 46 105
use OAI22X1  OAI22X1_87
timestamp 1745462530
transform 1 0 3576 0 -1 970
box -8 -3 46 105
use OAI22X1  OAI22X1_88
timestamp 1745462530
transform 1 0 3688 0 1 770
box -8 -3 46 105
use OAI22X1  OAI22X1_89
timestamp 1745462530
transform 1 0 872 0 1 1170
box -8 -3 46 105
use OAI22X1  OAI22X1_90
timestamp 1745462530
transform 1 0 1008 0 -1 970
box -8 -3 46 105
use OAI22X1  OAI22X1_91
timestamp 1745462530
transform 1 0 1464 0 1 2570
box -8 -3 46 105
use OAI22X1  OAI22X1_92
timestamp 1745462530
transform 1 0 1448 0 1 1770
box -8 -3 46 105
use OAI22X1  OAI22X1_93
timestamp 1745462530
transform 1 0 3192 0 -1 1970
box -8 -3 46 105
use OAI22X1  OAI22X1_94
timestamp 1745462530
transform 1 0 3360 0 -1 2170
box -8 -3 46 105
use OAI22X1  OAI22X1_95
timestamp 1745462530
transform 1 0 2736 0 -1 1170
box -8 -3 46 105
use OAI22X1  OAI22X1_96
timestamp 1745462530
transform 1 0 2784 0 -1 970
box -8 -3 46 105
use OAI22X1  OAI22X1_97
timestamp 1745462530
transform 1 0 1080 0 -1 1170
box -8 -3 46 105
use OAI22X1  OAI22X1_98
timestamp 1745462530
transform 1 0 1152 0 1 970
box -8 -3 46 105
use OAI22X1  OAI22X1_99
timestamp 1745462530
transform 1 0 848 0 1 1970
box -8 -3 46 105
use OAI22X1  OAI22X1_100
timestamp 1745462530
transform 1 0 1016 0 1 2170
box -8 -3 46 105
use OAI22X1  OAI22X1_101
timestamp 1745462530
transform 1 0 3264 0 1 2570
box -8 -3 46 105
use OAI22X1  OAI22X1_102
timestamp 1745462530
transform 1 0 3296 0 -1 2370
box -8 -3 46 105
use OAI22X1  OAI22X1_103
timestamp 1745462530
transform 1 0 3280 0 -1 1170
box -8 -3 46 105
use OAI22X1  OAI22X1_104
timestamp 1745462530
transform 1 0 3360 0 -1 970
box -8 -3 46 105
use OAI22X1  OAI22X1_105
timestamp 1745462530
transform 1 0 872 0 -1 1170
box -8 -3 46 105
use OAI22X1  OAI22X1_106
timestamp 1745462530
transform 1 0 944 0 -1 970
box -8 -3 46 105
use OAI22X1  OAI22X1_107
timestamp 1745462530
transform 1 0 1144 0 1 2570
box -8 -3 46 105
use OAI22X1  OAI22X1_108
timestamp 1745462530
transform 1 0 1080 0 -1 2170
box -8 -3 46 105
use OAI22X1  OAI22X1_109
timestamp 1745462530
transform 1 0 3024 0 -1 1970
box -8 -3 46 105
use OAI22X1  OAI22X1_110
timestamp 1745462530
transform 1 0 3296 0 -1 2170
box -8 -3 46 105
use OAI22X1  OAI22X1_111
timestamp 1745462530
transform 1 0 2360 0 1 970
box -8 -3 46 105
use OAI22X1  OAI22X1_112
timestamp 1745462530
transform 1 0 2424 0 1 970
box -8 -3 46 105
use OAI22X1  OAI22X1_113
timestamp 1745462530
transform 1 0 1712 0 -1 1170
box -8 -3 46 105
use OAI22X1  OAI22X1_114
timestamp 1745462530
transform 1 0 1696 0 1 970
box -8 -3 46 105
use OAI22X1  OAI22X1_115
timestamp 1745462530
transform 1 0 504 0 1 2170
box -8 -3 46 105
use OAI22X1  OAI22X1_116
timestamp 1745462530
transform 1 0 904 0 1 2170
box -8 -3 46 105
use OAI22X1  OAI22X1_117
timestamp 1745462530
transform 1 0 3992 0 -1 2570
box -8 -3 46 105
use OAI22X1  OAI22X1_118
timestamp 1745462530
transform 1 0 4096 0 -1 2370
box -8 -3 46 105
use OAI22X1  OAI22X1_119
timestamp 1745462530
transform 1 0 3928 0 -1 1170
box -8 -3 46 105
use OAI22X1  OAI22X1_120
timestamp 1745462530
transform 1 0 3976 0 1 970
box -8 -3 46 105
use OAI22X1  OAI22X1_121
timestamp 1745462530
transform 1 0 504 0 1 1170
box -8 -3 46 105
use OAI22X1  OAI22X1_122
timestamp 1745462530
transform 1 0 864 0 1 970
box -8 -3 46 105
use OAI22X1  OAI22X1_123
timestamp 1745462530
transform 1 0 2024 0 1 2370
box -8 -3 46 105
use OAI22X1  OAI22X1_124
timestamp 1745462530
transform 1 0 2032 0 -1 2170
box -8 -3 46 105
use OAI22X1  OAI22X1_125
timestamp 1745462530
transform 1 0 3904 0 -1 2170
box -8 -3 46 105
use OAI22X1  OAI22X1_126
timestamp 1745462530
transform 1 0 3936 0 1 1970
box -8 -3 46 105
use OAI22X1  OAI22X1_127
timestamp 1745462530
transform 1 0 3128 0 -1 1170
box -8 -3 46 105
use OAI22X1  OAI22X1_128
timestamp 1745462530
transform 1 0 3032 0 1 970
box -8 -3 46 105
use OAI22X1  OAI22X1_129
timestamp 1745462530
transform 1 0 1816 0 -1 1170
box -8 -3 46 105
use OAI22X1  OAI22X1_130
timestamp 1745462530
transform 1 0 1840 0 1 970
box -8 -3 46 105
use OAI22X1  OAI22X1_131
timestamp 1745462530
transform 1 0 576 0 1 1970
box -8 -3 46 105
use OAI22X1  OAI22X1_132
timestamp 1745462530
transform 1 0 880 0 -1 2170
box -8 -3 46 105
use OAI22X1  OAI22X1_133
timestamp 1745462530
transform 1 0 3984 0 1 2370
box -8 -3 46 105
use OAI22X1  OAI22X1_134
timestamp 1745462530
transform 1 0 4088 0 1 2170
box -8 -3 46 105
use OAI22X1  OAI22X1_135
timestamp 1745462530
transform 1 0 3976 0 -1 1170
box -8 -3 46 105
use OAI22X1  OAI22X1_136
timestamp 1745462530
transform 1 0 4040 0 1 970
box -8 -3 46 105
use OAI22X1  OAI22X1_137
timestamp 1745462530
transform 1 0 560 0 -1 1170
box -8 -3 46 105
use OAI22X1  OAI22X1_138
timestamp 1745462530
transform 1 0 976 0 -1 770
box -8 -3 46 105
use OAI22X1  OAI22X1_139
timestamp 1745462530
transform 1 0 1624 0 1 2570
box -8 -3 46 105
use OAI22X1  OAI22X1_140
timestamp 1745462530
transform 1 0 1632 0 -1 1970
box -8 -3 46 105
use OAI22X1  OAI22X1_141
timestamp 1745462530
transform 1 0 3000 0 -1 1570
box -8 -3 46 105
use OAI22X1  OAI22X1_142
timestamp 1745462530
transform 1 0 3192 0 1 1570
box -8 -3 46 105
use OAI22X1  OAI22X1_143
timestamp 1745462530
transform 1 0 2192 0 1 970
box -8 -3 46 105
use OAI22X1  OAI22X1_144
timestamp 1745462530
transform 1 0 2320 0 1 770
box -8 -3 46 105
use OAI22X1  OAI22X1_145
timestamp 1745462530
transform 1 0 1520 0 1 970
box -8 -3 46 105
use OAI22X1  OAI22X1_146
timestamp 1745462530
transform 1 0 1400 0 1 770
box -8 -3 46 105
use OAI22X1  OAI22X1_147
timestamp 1745462530
transform 1 0 624 0 -1 2370
box -8 -3 46 105
use OAI22X1  OAI22X1_148
timestamp 1745462530
transform 1 0 1040 0 1 1970
box -8 -3 46 105
use OAI22X1  OAI22X1_149
timestamp 1745462530
transform 1 0 3064 0 -1 2570
box -8 -3 46 105
use OAI22X1  OAI22X1_150
timestamp 1745462530
transform 1 0 3200 0 1 1970
box -8 -3 46 105
use OAI22X1  OAI22X1_151
timestamp 1745462530
transform 1 0 3096 0 1 970
box -8 -3 46 105
use OAI22X1  OAI22X1_152
timestamp 1745462530
transform 1 0 3184 0 1 770
box -8 -3 46 105
use OAI22X1  OAI22X1_153
timestamp 1745462530
transform 1 0 568 0 1 970
box -8 -3 46 105
use OAI22X1  OAI22X1_154
timestamp 1745462530
transform 1 0 1040 0 -1 770
box -8 -3 46 105
use OAI22X1  OAI22X1_155
timestamp 1745462530
transform 1 0 1336 0 1 2570
box -8 -3 46 105
use OAI22X1  OAI22X1_156
timestamp 1745462530
transform 1 0 1304 0 -1 1970
box -8 -3 46 105
use OAI22X1  OAI22X1_157
timestamp 1745462530
transform 1 0 3080 0 -1 1570
box -8 -3 46 105
use OAI22X1  OAI22X1_158
timestamp 1745462530
transform 1 0 3112 0 1 1570
box -8 -3 46 105
use OAI22X1  OAI22X1_159
timestamp 1745462530
transform 1 0 3064 0 -1 1170
box -8 -3 46 105
use OAI22X1  OAI22X1_160
timestamp 1745462530
transform 1 0 3096 0 1 770
box -8 -3 46 105
use OAI22X1  OAI22X1_161
timestamp 1745462530
transform 1 0 4024 0 1 3770
box -8 -3 46 105
use OAI22X1  OAI22X1_162
timestamp 1745462530
transform 1 0 3968 0 1 3770
box -8 -3 46 105
use OAI22X1  OAI22X1_163
timestamp 1745462530
transform 1 0 4144 0 -1 3770
box -8 -3 46 105
use OAI22X1  OAI22X1_164
timestamp 1745462530
transform 1 0 4040 0 -1 3770
box -8 -3 46 105
use OAI22X1  OAI22X1_165
timestamp 1745462530
transform 1 0 4152 0 1 3770
box -8 -3 46 105
use OAI22X1  OAI22X1_166
timestamp 1745462530
transform 1 0 4072 0 1 3770
box -8 -3 46 105
use OAI22X1  OAI22X1_167
timestamp 1745462530
transform 1 0 4224 0 -1 3770
box -8 -3 46 105
use OAI22X1  OAI22X1_168
timestamp 1745462530
transform 1 0 4096 0 -1 3770
box -8 -3 46 105
use OAI22X1  OAI22X1_169
timestamp 1745462530
transform 1 0 1560 0 -1 3170
box -8 -3 46 105
use OAI22X1  OAI22X1_170
timestamp 1745462530
transform 1 0 1608 0 -1 3170
box -8 -3 46 105
use OAI22X1  OAI22X1_171
timestamp 1745462530
transform 1 0 1872 0 1 2770
box -8 -3 46 105
use OAI22X1  OAI22X1_172
timestamp 1745462530
transform 1 0 1968 0 1 2170
box -8 -3 46 105
use OAI22X1  OAI22X1_173
timestamp 1745462530
transform 1 0 1888 0 1 2570
box -8 -3 46 105
use OAI22X1  OAI22X1_174
timestamp 1745462530
transform 1 0 1784 0 -1 2170
box -8 -3 46 105
use OAI22X1  OAI22X1_175
timestamp 1745462530
transform 1 0 1768 0 -1 2570
box -8 -3 46 105
use OAI22X1  OAI22X1_176
timestamp 1745462530
transform 1 0 1712 0 -1 1970
box -8 -3 46 105
use OAI22X1  OAI22X1_177
timestamp 1745462530
transform 1 0 360 0 -1 2570
box -8 -3 46 105
use OAI22X1  OAI22X1_178
timestamp 1745462530
transform 1 0 568 0 -1 2570
box -8 -3 46 105
use OAI22X1  OAI22X1_179
timestamp 1745462530
transform 1 0 200 0 -1 2570
box -8 -3 46 105
use OAI22X1  OAI22X1_180
timestamp 1745462530
transform 1 0 952 0 1 2370
box -8 -3 46 105
use OAI22X1  OAI22X1_181
timestamp 1745462530
transform 1 0 264 0 -1 2370
box -8 -3 46 105
use OAI22X1  OAI22X1_182
timestamp 1745462530
transform 1 0 272 0 -1 2170
box -8 -3 46 105
use OAI22X1  OAI22X1_183
timestamp 1745462530
transform 1 0 264 0 1 1770
box -8 -3 46 105
use OAI22X1  OAI22X1_184
timestamp 1745462530
transform 1 0 600 0 1 1770
box -8 -3 46 105
use OAI22X1  OAI22X1_185
timestamp 1745462530
transform 1 0 336 0 1 1570
box -8 -3 46 105
use OAI22X1  OAI22X1_186
timestamp 1745462530
transform 1 0 232 0 -1 970
box -8 -3 46 105
use OAI22X1  OAI22X1_187
timestamp 1745462530
transform 1 0 240 0 1 570
box -8 -3 46 105
use OAI22X1  OAI22X1_188
timestamp 1745462530
transform 1 0 456 0 -1 570
box -8 -3 46 105
use OAI22X1  OAI22X1_189
timestamp 1745462530
transform 1 0 696 0 1 370
box -8 -3 46 105
use OAI22X1  OAI22X1_190
timestamp 1745462530
transform 1 0 832 0 -1 570
box -8 -3 46 105
use OAI22X1  OAI22X1_191
timestamp 1745462530
transform 1 0 472 0 -1 1370
box -8 -3 46 105
use OAI22X1  OAI22X1_192
timestamp 1745462530
transform 1 0 672 0 -1 1370
box -8 -3 46 105
use OAI22X1  OAI22X1_193
timestamp 1745462530
transform 1 0 1480 0 -1 370
box -8 -3 46 105
use OAI22X1  OAI22X1_194
timestamp 1745462530
transform 1 0 1664 0 -1 570
box -8 -3 46 105
use OAI22X1  OAI22X1_195
timestamp 1745462530
transform 1 0 1648 0 1 370
box -8 -3 46 105
use OAI22X1  OAI22X1_196
timestamp 1745462530
transform 1 0 1720 0 -1 770
box -8 -3 46 105
use OAI22X1  OAI22X1_197
timestamp 1745462530
transform 1 0 1712 0 -1 370
box -8 -3 46 105
use OAI22X1  OAI22X1_198
timestamp 1745462530
transform 1 0 1776 0 1 970
box -8 -3 46 105
use OAI22X1  OAI22X1_199
timestamp 1745462530
transform 1 0 1824 0 1 1170
box -8 -3 46 105
use OAI22X1  OAI22X1_200
timestamp 1745462530
transform 1 0 1824 0 1 1370
box -8 -3 46 105
use OAI22X1  OAI22X1_201
timestamp 1745462530
transform 1 0 2888 0 1 170
box -8 -3 46 105
use OAI22X1  OAI22X1_202
timestamp 1745462530
transform 1 0 3016 0 1 570
box -8 -3 46 105
use OAI22X1  OAI22X1_203
timestamp 1745462530
transform 1 0 2800 0 1 170
box -8 -3 46 105
use OAI22X1  OAI22X1_204
timestamp 1745462530
transform 1 0 2920 0 1 370
box -8 -3 46 105
use OAI22X1  OAI22X1_205
timestamp 1745462530
transform 1 0 3096 0 1 170
box -8 -3 46 105
use OAI22X1  OAI22X1_206
timestamp 1745462530
transform 1 0 2896 0 1 970
box -8 -3 46 105
use OAI22X1  OAI22X1_207
timestamp 1745462530
transform 1 0 2840 0 1 1170
box -8 -3 46 105
use OAI22X1  OAI22X1_208
timestamp 1745462530
transform 1 0 2792 0 -1 1370
box -8 -3 46 105
use OAI22X1  OAI22X1_209
timestamp 1745462530
transform 1 0 3296 0 1 170
box -8 -3 46 105
use OAI22X1  OAI22X1_210
timestamp 1745462530
transform 1 0 3872 0 1 170
box -8 -3 46 105
use OAI22X1  OAI22X1_211
timestamp 1745462530
transform 1 0 4136 0 1 170
box -8 -3 46 105
use OAI22X1  OAI22X1_212
timestamp 1745462530
transform 1 0 3976 0 1 170
box -8 -3 46 105
use OAI22X1  OAI22X1_213
timestamp 1745462530
transform 1 0 4144 0 1 370
box -8 -3 46 105
use OAI22X1  OAI22X1_214
timestamp 1745462530
transform 1 0 4296 0 1 970
box -8 -3 46 105
use OAI22X1  OAI22X1_215
timestamp 1745462530
transform 1 0 4120 0 -1 1170
box -8 -3 46 105
use OAI22X1  OAI22X1_216
timestamp 1745462530
transform 1 0 3864 0 1 1170
box -8 -3 46 105
use OAI22X1  OAI22X1_217
timestamp 1745462530
transform 1 0 4096 0 -1 1770
box -8 -3 46 105
use OAI22X1  OAI22X1_218
timestamp 1745462530
transform 1 0 3816 0 1 1770
box -8 -3 46 105
use OAI22X1  OAI22X1_219
timestamp 1745462530
transform 1 0 4168 0 -1 1970
box -8 -3 46 105
use OAI22X1  OAI22X1_220
timestamp 1745462530
transform 1 0 3840 0 1 1970
box -8 -3 46 105
use OAI22X1  OAI22X1_221
timestamp 1745462530
transform 1 0 4208 0 1 1970
box -8 -3 46 105
use OAI22X1  OAI22X1_222
timestamp 1745462530
transform 1 0 3840 0 1 2170
box -8 -3 46 105
use OAI22X1  OAI22X1_223
timestamp 1745462530
transform 1 0 3104 0 1 2170
box -8 -3 46 105
use OAI22X1  OAI22X1_224
timestamp 1745462530
transform 1 0 2920 0 1 2170
box -8 -3 46 105
use OAI22X1  OAI22X1_225
timestamp 1745462530
transform 1 0 4176 0 -1 2770
box -8 -3 46 105
use OAI22X1  OAI22X1_226
timestamp 1745462530
transform 1 0 3904 0 1 2970
box -8 -3 46 105
use OAI22X1  OAI22X1_227
timestamp 1745462530
transform 1 0 4072 0 1 2770
box -8 -3 46 105
use OAI22X1  OAI22X1_228
timestamp 1745462530
transform 1 0 4160 0 1 2970
box -8 -3 46 105
use OAI22X1  OAI22X1_229
timestamp 1745462530
transform 1 0 4200 0 -1 2570
box -8 -3 46 105
use OAI22X1  OAI22X1_230
timestamp 1745462530
transform 1 0 4216 0 -1 2370
box -8 -3 46 105
use OAI22X1  OAI22X1_231
timestamp 1745462530
transform 1 0 4088 0 1 2970
box -8 -3 46 105
use OAI22X1  OAI22X1_232
timestamp 1745462530
transform 1 0 2864 0 1 2570
box -8 -3 46 105
use OAI22X1  OAI22X1_233
timestamp 1745462530
transform 1 0 2760 0 1 2770
box -8 -3 46 105
use OAI22X1  OAI22X1_234
timestamp 1745462530
transform 1 0 3904 0 -1 370
box -8 -3 46 105
use OAI22X1  OAI22X1_235
timestamp 1745462530
transform 1 0 3752 0 -1 370
box -8 -3 46 105
use OAI22X1  OAI22X1_236
timestamp 1745462530
transform 1 0 2928 0 -1 570
box -8 -3 46 105
use OAI22X1  OAI22X1_237
timestamp 1745462530
transform 1 0 2864 0 1 570
box -8 -3 46 105
use OAI22X1  OAI22X1_238
timestamp 1745462530
transform 1 0 4152 0 -1 2570
box -8 -3 46 105
use OAI22X1  OAI22X1_239
timestamp 1745462530
transform 1 0 3904 0 -1 1970
box -8 -3 46 105
use OAI22X1  OAI22X1_240
timestamp 1745462530
transform 1 0 3872 0 1 1770
box -8 -3 46 105
use OAI22X1  OAI22X1_241
timestamp 1745462530
transform 1 0 688 0 1 2370
box -8 -3 46 105
use OAI22X1  OAI22X1_242
timestamp 1745462530
transform 1 0 672 0 -1 2570
box -8 -3 46 105
use OAI22X1  OAI22X1_243
timestamp 1745462530
transform 1 0 1704 0 -1 2370
box -8 -3 46 105
use OAI22X1  OAI22X1_244
timestamp 1745462530
transform 1 0 1992 0 -1 2370
box -8 -3 46 105
use OAI22X1  OAI22X1_245
timestamp 1745462530
transform 1 0 1680 0 1 570
box -8 -3 46 105
use OAI22X1  OAI22X1_246
timestamp 1745462530
transform 1 0 1600 0 -1 570
box -8 -3 46 105
use OAI22X1  OAI22X1_247
timestamp 1745462530
transform 1 0 464 0 1 570
box -8 -3 46 105
use OAI22X1  OAI22X1_248
timestamp 1745462530
transform 1 0 312 0 -1 970
box -8 -3 46 105
use OAI22X1  OAI22X1_249
timestamp 1745462530
transform 1 0 1288 0 1 2770
box -8 -3 46 105
use OAI22X1  OAI22X1_250
timestamp 1745462530
transform 1 0 1280 0 1 2170
box -8 -3 46 105
use OAI22X1  OAI22X1_251
timestamp 1745462530
transform 1 0 1264 0 -1 2770
box -8 -3 46 105
use OAI22X1  OAI22X1_252
timestamp 1745462530
transform 1 0 1216 0 1 1970
box -8 -3 46 105
use OAI22X1  OAI22X1_253
timestamp 1745462530
transform 1 0 1232 0 -1 2570
box -8 -3 46 105
use OAI22X1  OAI22X1_254
timestamp 1745462530
transform 1 0 1224 0 -1 1970
box -8 -3 46 105
use OAI22X1  OAI22X1_255
timestamp 1745462530
transform 1 0 376 0 1 2770
box -8 -3 46 105
use OAI22X1  OAI22X1_256
timestamp 1745462530
transform 1 0 520 0 1 2770
box -8 -3 46 105
use OAI22X1  OAI22X1_257
timestamp 1745462530
transform 1 0 280 0 1 2770
box -8 -3 46 105
use OAI22X1  OAI22X1_258
timestamp 1745462530
transform 1 0 944 0 1 2770
box -8 -3 46 105
use OAI22X1  OAI22X1_259
timestamp 1745462530
transform 1 0 384 0 1 2370
box -8 -3 46 105
use OAI22X1  OAI22X1_260
timestamp 1745462530
transform 1 0 408 0 1 1970
box -8 -3 46 105
use OAI22X1  OAI22X1_261
timestamp 1745462530
transform 1 0 408 0 1 1770
box -8 -3 46 105
use OAI22X1  OAI22X1_262
timestamp 1745462530
transform 1 0 704 0 1 1770
box -8 -3 46 105
use OAI22X1  OAI22X1_263
timestamp 1745462530
transform 1 0 472 0 -1 1570
box -8 -3 46 105
use OAI22X1  OAI22X1_264
timestamp 1745462530
transform 1 0 368 0 -1 970
box -8 -3 46 105
use OAI22X1  OAI22X1_265
timestamp 1745462530
transform 1 0 312 0 1 170
box -8 -3 46 105
use OAI22X1  OAI22X1_266
timestamp 1745462530
transform 1 0 392 0 1 370
box -8 -3 46 105
use OAI22X1  OAI22X1_267
timestamp 1745462530
transform 1 0 624 0 -1 170
box -8 -3 46 105
use OAI22X1  OAI22X1_268
timestamp 1745462530
transform 1 0 888 0 1 170
box -8 -3 46 105
use OAI22X1  OAI22X1_269
timestamp 1745462530
transform 1 0 368 0 -1 1170
box -8 -3 46 105
use OAI22X1  OAI22X1_270
timestamp 1745462530
transform 1 0 688 0 1 1370
box -8 -3 46 105
use OAI22X1  OAI22X1_271
timestamp 1745462530
transform 1 0 1152 0 1 170
box -8 -3 46 105
use OAI22X1  OAI22X1_272
timestamp 1745462530
transform 1 0 1416 0 -1 570
box -8 -3 46 105
use OAI22X1  OAI22X1_273
timestamp 1745462530
transform 1 0 1440 0 1 170
box -8 -3 46 105
use OAI22X1  OAI22X1_274
timestamp 1745462530
transform 1 0 1408 0 -1 770
box -8 -3 46 105
use OAI22X1  OAI22X1_275
timestamp 1745462530
transform 1 0 1480 0 -1 170
box -8 -3 46 105
use OAI22X1  OAI22X1_276
timestamp 1745462530
transform 1 0 1584 0 -1 970
box -8 -3 46 105
use OAI22X1  OAI22X1_277
timestamp 1745462530
transform 1 0 1576 0 1 1170
box -8 -3 46 105
use OAI22X1  OAI22X1_278
timestamp 1745462530
transform 1 0 1648 0 1 1370
box -8 -3 46 105
use OAI22X1  OAI22X1_279
timestamp 1745462530
transform 1 0 2832 0 1 370
box -8 -3 46 105
use OAI22X1  OAI22X1_280
timestamp 1745462530
transform 1 0 3064 0 -1 770
box -8 -3 46 105
use OAI22X1  OAI22X1_281
timestamp 1745462530
transform 1 0 2656 0 -1 370
box -8 -3 46 105
use OAI22X1  OAI22X1_282
timestamp 1745462530
transform 1 0 2992 0 -1 570
box -8 -3 46 105
use OAI22X1  OAI22X1_283
timestamp 1745462530
transform 1 0 2952 0 -1 370
box -8 -3 46 105
use OAI22X1  OAI22X1_284
timestamp 1745462530
transform 1 0 2888 0 -1 970
box -8 -3 46 105
use OAI22X1  OAI22X1_285
timestamp 1745462530
transform 1 0 2824 0 -1 1170
box -8 -3 46 105
use OAI22X1  OAI22X1_286
timestamp 1745462530
transform 1 0 2832 0 1 1370
box -8 -3 46 105
use OAI22X1  OAI22X1_287
timestamp 1745462530
transform 1 0 3256 0 -1 370
box -8 -3 46 105
use OAI22X1  OAI22X1_288
timestamp 1745462530
transform 1 0 3344 0 1 370
box -8 -3 46 105
use OAI22X1  OAI22X1_289
timestamp 1745462530
transform 1 0 4064 0 1 370
box -8 -3 46 105
use OAI22X1  OAI22X1_290
timestamp 1745462530
transform 1 0 3360 0 1 570
box -8 -3 46 105
use OAI22X1  OAI22X1_291
timestamp 1745462530
transform 1 0 4136 0 1 570
box -8 -3 46 105
use OAI22X1  OAI22X1_292
timestamp 1745462530
transform 1 0 4048 0 1 770
box -8 -3 46 105
use OAI22X1  OAI22X1_293
timestamp 1745462530
transform 1 0 3376 0 1 970
box -8 -3 46 105
use OAI22X1  OAI22X1_294
timestamp 1745462530
transform 1 0 3360 0 1 1170
box -8 -3 46 105
use OAI22X1  OAI22X1_295
timestamp 1745462530
transform 1 0 4072 0 1 1370
box -8 -3 46 105
use OAI22X1  OAI22X1_296
timestamp 1745462530
transform 1 0 3496 0 1 1370
box -8 -3 46 105
use OAI22X1  OAI22X1_297
timestamp 1745462530
transform 1 0 4056 0 -1 1570
box -8 -3 46 105
use OAI22X1  OAI22X1_298
timestamp 1745462530
transform 1 0 3560 0 1 1570
box -8 -3 46 105
use OAI22X1  OAI22X1_299
timestamp 1745462530
transform 1 0 4152 0 1 1570
box -8 -3 46 105
use OAI22X1  OAI22X1_300
timestamp 1745462530
transform 1 0 3272 0 -1 1770
box -8 -3 46 105
use OAI22X1  OAI22X1_301
timestamp 1745462530
transform 1 0 2760 0 -1 1770
box -8 -3 46 105
use OAI22X1  OAI22X1_302
timestamp 1745462530
transform 1 0 2760 0 1 1770
box -8 -3 46 105
use OAI22X1  OAI22X1_303
timestamp 1745462530
transform 1 0 3264 0 -1 2770
box -8 -3 46 105
use OAI22X1  OAI22X1_304
timestamp 1745462530
transform 1 0 2992 0 -1 2970
box -8 -3 46 105
use OAI22X1  OAI22X1_305
timestamp 1745462530
transform 1 0 3240 0 1 2770
box -8 -3 46 105
use OAI22X1  OAI22X1_306
timestamp 1745462530
transform 1 0 3192 0 1 2970
box -8 -3 46 105
use OAI22X1  OAI22X1_307
timestamp 1745462530
transform 1 0 3272 0 1 2370
box -8 -3 46 105
use OAI22X1  OAI22X1_308
timestamp 1745462530
transform 1 0 3232 0 -1 2370
box -8 -3 46 105
use OAI22X1  OAI22X1_309
timestamp 1745462530
transform 1 0 3168 0 -1 2970
box -8 -3 46 105
use OAI22X1  OAI22X1_310
timestamp 1745462530
transform 1 0 2744 0 1 2370
box -8 -3 46 105
use OAI22X1  OAI22X1_311
timestamp 1745462530
transform 1 0 2784 0 -1 2770
box -8 -3 46 105
use OAI22X1  OAI22X1_312
timestamp 1745462530
transform 1 0 3360 0 -1 570
box -8 -3 46 105
use OAI22X1  OAI22X1_313
timestamp 1745462530
transform 1 0 3264 0 -1 570
box -8 -3 46 105
use OAI22X1  OAI22X1_314
timestamp 1745462530
transform 1 0 2824 0 -1 570
box -8 -3 46 105
use OAI22X1  OAI22X1_315
timestamp 1745462530
transform 1 0 2920 0 -1 770
box -8 -3 46 105
use OAI22X1  OAI22X1_316
timestamp 1745462530
transform 1 0 3192 0 1 2370
box -8 -3 46 105
use OAI22X1  OAI22X1_317
timestamp 1745462530
transform 1 0 3464 0 -1 1570
box -8 -3 46 105
use OAI22X1  OAI22X1_318
timestamp 1745462530
transform 1 0 3400 0 1 1370
box -8 -3 46 105
use OAI22X1  OAI22X1_319
timestamp 1745462530
transform 1 0 728 0 1 2770
box -8 -3 46 105
use OAI22X1  OAI22X1_320
timestamp 1745462530
transform 1 0 648 0 1 2770
box -8 -3 46 105
use OAI22X1  OAI22X1_321
timestamp 1745462530
transform 1 0 1184 0 -1 2370
box -8 -3 46 105
use OAI22X1  OAI22X1_322
timestamp 1745462530
transform 1 0 1248 0 -1 2370
box -8 -3 46 105
use OAI22X1  OAI22X1_323
timestamp 1745462530
transform 1 0 1416 0 1 570
box -8 -3 46 105
use OAI22X1  OAI22X1_324
timestamp 1745462530
transform 1 0 1344 0 -1 570
box -8 -3 46 105
use OAI22X1  OAI22X1_325
timestamp 1745462530
transform 1 0 368 0 1 570
box -8 -3 46 105
use OAI22X1  OAI22X1_326
timestamp 1745462530
transform 1 0 480 0 1 770
box -8 -3 46 105
use OAI22X1  OAI22X1_327
timestamp 1745462530
transform 1 0 1736 0 1 2770
box -8 -3 46 105
use OAI22X1  OAI22X1_328
timestamp 1745462530
transform 1 0 1688 0 1 2170
box -8 -3 46 105
use OAI22X1  OAI22X1_329
timestamp 1745462530
transform 1 0 1672 0 -1 2770
box -8 -3 46 105
use OAI22X1  OAI22X1_330
timestamp 1745462530
transform 1 0 1576 0 1 1970
box -8 -3 46 105
use OAI22X1  OAI22X1_331
timestamp 1745462530
transform 1 0 1512 0 -1 2570
box -8 -3 46 105
use OAI22X1  OAI22X1_332
timestamp 1745462530
transform 1 0 1552 0 -1 1970
box -8 -3 46 105
use OAI22X1  OAI22X1_333
timestamp 1745462530
transform 1 0 416 0 -1 2770
box -8 -3 46 105
use OAI22X1  OAI22X1_334
timestamp 1745462530
transform 1 0 504 0 1 2570
box -8 -3 46 105
use OAI22X1  OAI22X1_335
timestamp 1745462530
transform 1 0 328 0 1 2570
box -8 -3 46 105
use OAI22X1  OAI22X1_336
timestamp 1745462530
transform 1 0 944 0 1 2570
box -8 -3 46 105
use OAI22X1  OAI22X1_337
timestamp 1745462530
transform 1 0 344 0 -1 2370
box -8 -3 46 105
use OAI22X1  OAI22X1_338
timestamp 1745462530
transform 1 0 456 0 -1 2170
box -8 -3 46 105
use OAI22X1  OAI22X1_339
timestamp 1745462530
transform 1 0 416 0 -1 1770
box -8 -3 46 105
use OAI22X1  OAI22X1_340
timestamp 1745462530
transform 1 0 560 0 1 1570
box -8 -3 46 105
use OAI22X1  OAI22X1_341
timestamp 1745462530
transform 1 0 408 0 -1 1570
box -8 -3 46 105
use OAI22X1  OAI22X1_342
timestamp 1745462530
transform 1 0 360 0 1 770
box -8 -3 46 105
use OAI22X1  OAI22X1_343
timestamp 1745462530
transform 1 0 240 0 1 170
box -8 -3 46 105
use OAI22X1  OAI22X1_344
timestamp 1745462530
transform 1 0 312 0 1 370
box -8 -3 46 105
use OAI22X1  OAI22X1_345
timestamp 1745462530
transform 1 0 528 0 -1 170
box -8 -3 46 105
use OAI22X1  OAI22X1_346
timestamp 1745462530
transform 1 0 824 0 1 170
box -8 -3 46 105
use OAI22X1  OAI22X1_347
timestamp 1745462530
transform 1 0 304 0 1 1170
box -8 -3 46 105
use OAI22X1  OAI22X1_348
timestamp 1745462530
transform 1 0 752 0 1 1370
box -8 -3 46 105
use OAI22X1  OAI22X1_349
timestamp 1745462530
transform 1 0 1680 0 1 170
box -8 -3 46 105
use OAI22X1  OAI22X1_350
timestamp 1745462530
transform 1 0 1824 0 1 370
box -8 -3 46 105
use OAI22X1  OAI22X1_351
timestamp 1745462530
transform 1 0 1784 0 1 170
box -8 -3 46 105
use OAI22X1  OAI22X1_352
timestamp 1745462530
transform 1 0 1816 0 -1 770
box -8 -3 46 105
use OAI22X1  OAI22X1_353
timestamp 1745462530
transform 1 0 1888 0 -1 170
box -8 -3 46 105
use OAI22X1  OAI22X1_354
timestamp 1745462530
transform 1 0 2016 0 1 970
box -8 -3 46 105
use OAI22X1  OAI22X1_355
timestamp 1745462530
transform 1 0 1984 0 1 1170
box -8 -3 46 105
use OAI22X1  OAI22X1_356
timestamp 1745462530
transform 1 0 1920 0 1 1370
box -8 -3 46 105
use OAI22X1  OAI22X1_357
timestamp 1745462530
transform 1 0 2224 0 -1 370
box -8 -3 46 105
use OAI22X1  OAI22X1_358
timestamp 1745462530
transform 1 0 2184 0 1 570
box -8 -3 46 105
use OAI22X1  OAI22X1_359
timestamp 1745462530
transform 1 0 2216 0 1 170
box -8 -3 46 105
use OAI22X1  OAI22X1_360
timestamp 1745462530
transform 1 0 2224 0 1 370
box -8 -3 46 105
use OAI22X1  OAI22X1_361
timestamp 1745462530
transform 1 0 2488 0 -1 170
box -8 -3 46 105
use OAI22X1  OAI22X1_362
timestamp 1745462530
transform 1 0 2336 0 -1 970
box -8 -3 46 105
use OAI22X1  OAI22X1_363
timestamp 1745462530
transform 1 0 2288 0 -1 1170
box -8 -3 46 105
use OAI22X1  OAI22X1_364
timestamp 1745462530
transform 1 0 2360 0 -1 1370
box -8 -3 46 105
use OAI22X1  OAI22X1_365
timestamp 1745462530
transform 1 0 3424 0 1 170
box -8 -3 46 105
use OAI22X1  OAI22X1_366
timestamp 1745462530
transform 1 0 3800 0 1 170
box -8 -3 46 105
use OAI22X1  OAI22X1_367
timestamp 1745462530
transform 1 0 4208 0 1 170
box -8 -3 46 105
use OAI22X1  OAI22X1_368
timestamp 1745462530
transform 1 0 3976 0 -1 370
box -8 -3 46 105
use OAI22X1  OAI22X1_369
timestamp 1745462530
transform 1 0 4296 0 -1 370
box -8 -3 46 105
use OAI22X1  OAI22X1_370
timestamp 1745462530
transform 1 0 4232 0 -1 970
box -8 -3 46 105
use OAI22X1  OAI22X1_371
timestamp 1745462530
transform 1 0 4208 0 1 970
box -8 -3 46 105
use OAI22X1  OAI22X1_372
timestamp 1745462530
transform 1 0 3912 0 1 1170
box -8 -3 46 105
use OAI22X1  OAI22X1_373
timestamp 1745462530
transform 1 0 4200 0 -1 1370
box -8 -3 46 105
use OAI22X1  OAI22X1_374
timestamp 1745462530
transform 1 0 3664 0 1 1370
box -8 -3 46 105
use OAI22X1  OAI22X1_375
timestamp 1745462530
transform 1 0 4208 0 -1 1570
box -8 -3 46 105
use OAI22X1  OAI22X1_376
timestamp 1745462530
transform 1 0 3640 0 1 1570
box -8 -3 46 105
use OAI22X1  OAI22X1_377
timestamp 1745462530
transform 1 0 4304 0 1 1570
box -8 -3 46 105
use OAI22X1  OAI22X1_378
timestamp 1745462530
transform 1 0 3264 0 1 1770
box -8 -3 46 105
use OAI22X1  OAI22X1_379
timestamp 1745462530
transform 1 0 2856 0 1 1770
box -8 -3 46 105
use OAI22X1  OAI22X1_380
timestamp 1745462530
transform 1 0 2656 0 -1 1970
box -8 -3 46 105
use OAI22X1  OAI22X1_381
timestamp 1745462530
transform 1 0 4184 0 1 2570
box -8 -3 46 105
use OAI22X1  OAI22X1_382
timestamp 1745462530
transform 1 0 3888 0 -1 2970
box -8 -3 46 105
use OAI22X1  OAI22X1_383
timestamp 1745462530
transform 1 0 4136 0 1 2770
box -8 -3 46 105
use OAI22X1  OAI22X1_384
timestamp 1745462530
transform 1 0 4216 0 -1 2970
box -8 -3 46 105
use OAI22X1  OAI22X1_385
timestamp 1745462530
transform 1 0 4208 0 1 2370
box -8 -3 46 105
use OAI22X1  OAI22X1_386
timestamp 1745462530
transform 1 0 4168 0 -1 2370
box -8 -3 46 105
use OAI22X1  OAI22X1_387
timestamp 1745462530
transform 1 0 4048 0 -1 2970
box -8 -3 46 105
use OAI22X1  OAI22X1_388
timestamp 1745462530
transform 1 0 2816 0 1 2370
box -8 -3 46 105
use OAI22X1  OAI22X1_389
timestamp 1745462530
transform 1 0 2600 0 1 2770
box -8 -3 46 105
use OAI22X1  OAI22X1_390
timestamp 1745462530
transform 1 0 3904 0 1 370
box -8 -3 46 105
use OAI22X1  OAI22X1_391
timestamp 1745462530
transform 1 0 3800 0 1 370
box -8 -3 46 105
use OAI22X1  OAI22X1_392
timestamp 1745462530
transform 1 0 2384 0 -1 570
box -8 -3 46 105
use OAI22X1  OAI22X1_393
timestamp 1745462530
transform 1 0 2248 0 1 570
box -8 -3 46 105
use OAI22X1  OAI22X1_394
timestamp 1745462530
transform 1 0 4136 0 1 2370
box -8 -3 46 105
use OAI22X1  OAI22X1_395
timestamp 1745462530
transform 1 0 3616 0 -1 1570
box -8 -3 46 105
use OAI22X1  OAI22X1_396
timestamp 1745462530
transform 1 0 3568 0 1 1370
box -8 -3 46 105
use OAI22X1  OAI22X1_397
timestamp 1745462530
transform 1 0 712 0 1 2570
box -8 -3 46 105
use OAI22X1  OAI22X1_398
timestamp 1745462530
transform 1 0 624 0 1 2570
box -8 -3 46 105
use OAI22X1  OAI22X1_399
timestamp 1745462530
transform 1 0 1552 0 -1 2370
box -8 -3 46 105
use OAI22X1  OAI22X1_400
timestamp 1745462530
transform 1 0 1648 0 -1 2370
box -8 -3 46 105
use OAI22X1  OAI22X1_401
timestamp 1745462530
transform 1 0 1792 0 1 570
box -8 -3 46 105
use OAI22X1  OAI22X1_402
timestamp 1745462530
transform 1 0 1848 0 -1 570
box -8 -3 46 105
use OAI22X1  OAI22X1_403
timestamp 1745462530
transform 1 0 352 0 -1 570
box -8 -3 46 105
use OAI22X1  OAI22X1_404
timestamp 1745462530
transform 1 0 400 0 -1 770
box -8 -3 46 105
use OAI22X1  OAI22X1_405
timestamp 1745462530
transform 1 0 1800 0 1 2770
box -8 -3 46 105
use OAI22X1  OAI22X1_406
timestamp 1745462530
transform 1 0 1888 0 1 2170
box -8 -3 46 105
use OAI22X1  OAI22X1_407
timestamp 1745462530
transform 1 0 1816 0 1 2570
box -8 -3 46 105
use OAI22X1  OAI22X1_408
timestamp 1745462530
transform 1 0 1824 0 1 1970
box -8 -3 46 105
use OAI22X1  OAI22X1_409
timestamp 1745462530
transform 1 0 1704 0 -1 2570
box -8 -3 46 105
use OAI22X1  OAI22X1_410
timestamp 1745462530
transform 1 0 1784 0 -1 1970
box -8 -3 46 105
use OAI22X1  OAI22X1_411
timestamp 1745462530
transform 1 0 744 0 -1 2970
box -8 -3 46 105
use OAI22X1  OAI22X1_412
timestamp 1745462530
transform 1 0 672 0 -1 2970
box -8 -3 46 105
use OAI22X1  OAI22X1_413
timestamp 1745462530
transform 1 0 432 0 1 2770
box -8 -3 46 105
use OAI22X1  OAI22X1_414
timestamp 1745462530
transform 1 0 896 0 -1 2970
box -8 -3 46 105
use OAI22X1  OAI22X1_415
timestamp 1745462530
transform 1 0 312 0 1 2170
box -8 -3 46 105
use OAI22X1  OAI22X1_416
timestamp 1745462530
transform 1 0 344 0 1 1970
box -8 -3 46 105
use OAI22X1  OAI22X1_417
timestamp 1745462530
transform 1 0 328 0 1 1770
box -8 -3 46 105
use OAI22X1  OAI22X1_418
timestamp 1745462530
transform 1 0 648 0 -1 1770
box -8 -3 46 105
use OAI22X1  OAI22X1_419
timestamp 1745462530
transform 1 0 344 0 -1 1570
box -8 -3 46 105
use OAI22X1  OAI22X1_420
timestamp 1745462530
transform 1 0 192 0 1 770
box -8 -3 46 105
use OAI22X1  OAI22X1_421
timestamp 1745462530
transform 1 0 192 0 -1 370
box -8 -3 46 105
use OAI22X1  OAI22X1_422
timestamp 1745462530
transform 1 0 200 0 1 370
box -8 -3 46 105
use OAI22X1  OAI22X1_423
timestamp 1745462530
transform 1 0 696 0 -1 370
box -8 -3 46 105
use OAI22X1  OAI22X1_424
timestamp 1745462530
transform 1 0 888 0 -1 370
box -8 -3 46 105
use OAI22X1  OAI22X1_425
timestamp 1745462530
transform 1 0 184 0 -1 1170
box -8 -3 46 105
use OAI22X1  OAI22X1_426
timestamp 1745462530
transform 1 0 832 0 1 1370
box -8 -3 46 105
use OAI22X1  OAI22X1_427
timestamp 1745462530
transform 1 0 1616 0 -1 370
box -8 -3 46 105
use OAI22X1  OAI22X1_428
timestamp 1745462530
transform 1 0 1912 0 1 370
box -8 -3 46 105
use OAI22X1  OAI22X1_429
timestamp 1745462530
transform 1 0 1880 0 1 170
box -8 -3 46 105
use OAI22X1  OAI22X1_430
timestamp 1745462530
transform 1 0 1880 0 -1 770
box -8 -3 46 105
use OAI22X1  OAI22X1_431
timestamp 1745462530
transform 1 0 1888 0 -1 370
box -8 -3 46 105
use OAI22X1  OAI22X1_432
timestamp 1745462530
transform 1 0 1992 0 -1 970
box -8 -3 46 105
use OAI22X1  OAI22X1_433
timestamp 1745462530
transform 1 0 1992 0 -1 1170
box -8 -3 46 105
use OAI22X1  OAI22X1_434
timestamp 1745462530
transform 1 0 1984 0 -1 1370
box -8 -3 46 105
use OAI22X1  OAI22X1_435
timestamp 1745462530
transform 1 0 2352 0 -1 370
box -8 -3 46 105
use OAI22X1  OAI22X1_436
timestamp 1745462530
transform 1 0 2272 0 -1 770
box -8 -3 46 105
use OAI22X1  OAI22X1_437
timestamp 1745462530
transform 1 0 2504 0 -1 370
box -8 -3 46 105
use OAI22X1  OAI22X1_438
timestamp 1745462530
transform 1 0 2288 0 1 370
box -8 -3 46 105
use OAI22X1  OAI22X1_439
timestamp 1745462530
transform 1 0 2440 0 -1 370
box -8 -3 46 105
use OAI22X1  OAI22X1_440
timestamp 1745462530
transform 1 0 2272 0 -1 970
box -8 -3 46 105
use OAI22X1  OAI22X1_441
timestamp 1745462530
transform 1 0 2592 0 -1 1170
box -8 -3 46 105
use OAI22X1  OAI22X1_442
timestamp 1745462530
transform 1 0 2592 0 -1 1370
box -8 -3 46 105
use OAI22X1  OAI22X1_443
timestamp 1745462530
transform 1 0 3368 0 -1 370
box -8 -3 46 105
use OAI22X1  OAI22X1_444
timestamp 1745462530
transform 1 0 3728 0 1 370
box -8 -3 46 105
use OAI22X1  OAI22X1_445
timestamp 1745462530
transform 1 0 4208 0 1 370
box -8 -3 46 105
use OAI22X1  OAI22X1_446
timestamp 1745462530
transform 1 0 3768 0 1 570
box -8 -3 46 105
use OAI22X1  OAI22X1_447
timestamp 1745462530
transform 1 0 4208 0 -1 570
box -8 -3 46 105
use OAI22X1  OAI22X1_448
timestamp 1745462530
transform 1 0 4136 0 1 770
box -8 -3 46 105
use OAI22X1  OAI22X1_449
timestamp 1745462530
transform 1 0 3792 0 1 970
box -8 -3 46 105
use OAI22X1  OAI22X1_450
timestamp 1745462530
transform 1 0 3768 0 1 1170
box -8 -3 46 105
use OAI22X1  OAI22X1_451
timestamp 1745462530
transform 1 0 4136 0 1 1370
box -8 -3 46 105
use OAI22X1  OAI22X1_452
timestamp 1745462530
transform 1 0 3792 0 1 1370
box -8 -3 46 105
use OAI22X1  OAI22X1_453
timestamp 1745462530
transform 1 0 4200 0 1 1370
box -8 -3 46 105
use OAI22X1  OAI22X1_454
timestamp 1745462530
transform 1 0 3800 0 1 1570
box -8 -3 46 105
use OAI22X1  OAI22X1_455
timestamp 1745462530
transform 1 0 3976 0 -1 1570
box -8 -3 46 105
use OAI22X1  OAI22X1_456
timestamp 1745462530
transform 1 0 3864 0 -1 1770
box -8 -3 46 105
use OAI22X1  OAI22X1_457
timestamp 1745462530
transform 1 0 2960 0 1 1770
box -8 -3 46 105
use OAI22X1  OAI22X1_458
timestamp 1745462530
transform 1 0 2688 0 1 1770
box -8 -3 46 105
use OAI22X1  OAI22X1_459
timestamp 1745462530
transform 1 0 3856 0 -1 2770
box -8 -3 46 105
use OAI22X1  OAI22X1_460
timestamp 1745462530
transform 1 0 3752 0 1 2970
box -8 -3 46 105
use OAI22X1  OAI22X1_461
timestamp 1745462530
transform 1 0 3848 0 1 2770
box -8 -3 46 105
use OAI22X1  OAI22X1_462
timestamp 1745462530
transform 1 0 3720 0 -1 2970
box -8 -3 46 105
use OAI22X1  OAI22X1_463
timestamp 1745462530
transform 1 0 3824 0 -1 2570
box -8 -3 46 105
use OAI22X1  OAI22X1_464
timestamp 1745462530
transform 1 0 3920 0 -1 2370
box -8 -3 46 105
use OAI22X1  OAI22X1_465
timestamp 1745462530
transform 1 0 3832 0 1 2970
box -8 -3 46 105
use OAI22X1  OAI22X1_466
timestamp 1745462530
transform 1 0 2960 0 1 2370
box -8 -3 46 105
use OAI22X1  OAI22X1_467
timestamp 1745462530
transform 1 0 2488 0 1 2770
box -8 -3 46 105
use OAI22X1  OAI22X1_468
timestamp 1745462530
transform 1 0 3704 0 1 570
box -8 -3 46 105
use OAI22X1  OAI22X1_469
timestamp 1745462530
transform 1 0 3600 0 -1 570
box -8 -3 46 105
use OAI22X1  OAI22X1_470
timestamp 1745462530
transform 1 0 2504 0 -1 570
box -8 -3 46 105
use OAI22X1  OAI22X1_471
timestamp 1745462530
transform 1 0 2456 0 -1 770
box -8 -3 46 105
use OAI22X1  OAI22X1_472
timestamp 1745462530
transform 1 0 3880 0 1 2370
box -8 -3 46 105
use OAI22X1  OAI22X1_473
timestamp 1745462530
transform 1 0 3864 0 -1 1570
box -8 -3 46 105
use OAI22X1  OAI22X1_474
timestamp 1745462530
transform 1 0 3872 0 1 1370
box -8 -3 46 105
use OAI22X1  OAI22X1_475
timestamp 1745462530
transform 1 0 856 0 1 2770
box -8 -3 46 105
use OAI22X1  OAI22X1_476
timestamp 1745462530
transform 1 0 776 0 1 2770
box -8 -3 46 105
use OAI22X1  OAI22X1_477
timestamp 1745462530
transform 1 0 1768 0 -1 2370
box -8 -3 46 105
use OAI22X1  OAI22X1_478
timestamp 1745462530
transform 1 0 1856 0 -1 2370
box -8 -3 46 105
use OAI22X1  OAI22X1_479
timestamp 1745462530
transform 1 0 1936 0 1 570
box -8 -3 46 105
use OAI22X1  OAI22X1_480
timestamp 1745462530
transform 1 0 1920 0 -1 570
box -8 -3 46 105
use OAI22X1  OAI22X1_481
timestamp 1745462530
transform 1 0 296 0 -1 570
box -8 -3 46 105
use OAI22X1  OAI22X1_482
timestamp 1745462530
transform 1 0 296 0 -1 770
box -8 -3 46 105
use OAI22X1  OAI22X1_483
timestamp 1745462530
transform 1 0 1232 0 1 2770
box -8 -3 46 105
use OAI22X1  OAI22X1_484
timestamp 1745462530
transform 1 0 1216 0 1 2170
box -8 -3 46 105
use OAI22X1  OAI22X1_485
timestamp 1745462530
transform 1 0 1216 0 -1 2770
box -8 -3 46 105
use OAI22X1  OAI22X1_486
timestamp 1745462530
transform 1 0 1192 0 -1 2170
box -8 -3 46 105
use OAI22X1  OAI22X1_487
timestamp 1745462530
transform 1 0 1176 0 -1 2570
box -8 -3 46 105
use OAI22X1  OAI22X1_488
timestamp 1745462530
transform 1 0 1152 0 -1 1970
box -8 -3 46 105
use OAI22X1  OAI22X1_489
timestamp 1745462530
transform 1 0 824 0 -1 2970
box -8 -3 46 105
use OAI22X1  OAI22X1_490
timestamp 1745462530
transform 1 0 768 0 1 2570
box -8 -3 46 105
use OAI22X1  OAI22X1_491
timestamp 1745462530
transform 1 0 208 0 -1 2770
box -8 -3 46 105
use OAI22X1  OAI22X1_492
timestamp 1745462530
transform 1 0 944 0 -1 2970
box -8 -3 46 105
use OAI22X1  OAI22X1_493
timestamp 1745462530
transform 1 0 192 0 -1 2370
box -8 -3 46 105
use OAI22X1  OAI22X1_494
timestamp 1745462530
transform 1 0 200 0 -1 2170
box -8 -3 46 105
use OAI22X1  OAI22X1_495
timestamp 1745462530
transform 1 0 200 0 -1 1770
box -8 -3 46 105
use OAI22X1  OAI22X1_496
timestamp 1745462530
transform 1 0 672 0 1 1570
box -8 -3 46 105
use OAI22X1  OAI22X1_497
timestamp 1745462530
transform 1 0 208 0 -1 1570
box -8 -3 46 105
use OAI22X1  OAI22X1_498
timestamp 1745462530
transform 1 0 192 0 1 970
box -8 -3 46 105
use OAI22X1  OAI22X1_499
timestamp 1745462530
transform 1 0 224 0 -1 570
box -8 -3 46 105
use OAI22X1  OAI22X1_500
timestamp 1745462530
transform 1 0 192 0 1 570
box -8 -3 46 105
use OAI22X1  OAI22X1_501
timestamp 1745462530
transform 1 0 672 0 -1 570
box -8 -3 46 105
use OAI22X1  OAI22X1_502
timestamp 1745462530
transform 1 0 904 0 -1 570
box -8 -3 46 105
use OAI22X1  OAI22X1_503
timestamp 1745462530
transform 1 0 200 0 -1 1370
box -8 -3 46 105
use OAI22X1  OAI22X1_504
timestamp 1745462530
transform 1 0 936 0 -1 1370
box -8 -3 46 105
use OAI22X1  OAI22X1_505
timestamp 1745462530
transform 1 0 1112 0 -1 370
box -8 -3 46 105
use OAI22X1  OAI22X1_506
timestamp 1745462530
transform 1 0 1144 0 1 370
box -8 -3 46 105
use OAI22X1  OAI22X1_507
timestamp 1745462530
transform 1 0 1312 0 -1 370
box -8 -3 46 105
use OAI22X1  OAI22X1_508
timestamp 1745462530
transform 1 0 1336 0 -1 770
box -8 -3 46 105
use OAI22X1  OAI22X1_509
timestamp 1745462530
transform 1 0 1408 0 -1 370
box -8 -3 46 105
use OAI22X1  OAI22X1_510
timestamp 1745462530
transform 1 0 1408 0 1 970
box -8 -3 46 105
use OAI22X1  OAI22X1_511
timestamp 1745462530
transform 1 0 1456 0 -1 1370
box -8 -3 46 105
use OAI22X1  OAI22X1_512
timestamp 1745462530
transform 1 0 1512 0 1 1370
box -8 -3 46 105
use OAI22X1  OAI22X1_513
timestamp 1745462530
transform 1 0 2288 0 -1 370
box -8 -3 46 105
use OAI22X1  OAI22X1_514
timestamp 1745462530
transform 1 0 2184 0 -1 770
box -8 -3 46 105
use OAI22X1  OAI22X1_515
timestamp 1745462530
transform 1 0 2288 0 1 170
box -8 -3 46 105
use OAI22X1  OAI22X1_516
timestamp 1745462530
transform 1 0 2280 0 -1 570
box -8 -3 46 105
use OAI22X1  OAI22X1_517
timestamp 1745462530
transform 1 0 2592 0 -1 370
box -8 -3 46 105
use OAI22X1  OAI22X1_518
timestamp 1745462530
transform 1 0 2544 0 -1 970
box -8 -3 46 105
use OAI22X1  OAI22X1_519
timestamp 1745462530
transform 1 0 2352 0 -1 1170
box -8 -3 46 105
use OAI22X1  OAI22X1_520
timestamp 1745462530
transform 1 0 2384 0 1 1370
box -8 -3 46 105
use OAI22X1  OAI22X1_521
timestamp 1745462530
transform 1 0 3312 0 -1 370
box -8 -3 46 105
use OAI22X1  OAI22X1_522
timestamp 1745462530
transform 1 0 3512 0 1 370
box -8 -3 46 105
use OAI22X1  OAI22X1_523
timestamp 1745462530
transform 1 0 4000 0 1 370
box -8 -3 46 105
use OAI22X1  OAI22X1_524
timestamp 1745462530
transform 1 0 3504 0 1 570
box -8 -3 46 105
use OAI22X1  OAI22X1_525
timestamp 1745462530
transform 1 0 4080 0 1 570
box -8 -3 46 105
use OAI22X1  OAI22X1_526
timestamp 1745462530
transform 1 0 3944 0 1 770
box -8 -3 46 105
use OAI22X1  OAI22X1_527
timestamp 1745462530
transform 1 0 3440 0 1 970
box -8 -3 46 105
use OAI22X1  OAI22X1_528
timestamp 1745462530
transform 1 0 3440 0 1 1170
box -8 -3 46 105
use OAI22X1  OAI22X1_529
timestamp 1745462530
transform 1 0 4080 0 1 1570
box -8 -3 46 105
use OAI22X1  OAI22X1_530
timestamp 1745462530
transform 1 0 3464 0 1 1770
box -8 -3 46 105
use OAI22X1  OAI22X1_531
timestamp 1745462530
transform 1 0 4104 0 -1 1970
box -8 -3 46 105
use OAI22X1  OAI22X1_532
timestamp 1745462530
transform 1 0 3672 0 1 1970
box -8 -3 46 105
use OAI22X1  OAI22X1_533
timestamp 1745462530
transform 1 0 4128 0 1 1970
box -8 -3 46 105
use OAI22X1  OAI22X1_534
timestamp 1745462530
transform 1 0 3368 0 1 2170
box -8 -3 46 105
use OAI22X1  OAI22X1_535
timestamp 1745462530
transform 1 0 2776 0 1 2170
box -8 -3 46 105
use OAI22X1  OAI22X1_536
timestamp 1745462530
transform 1 0 2616 0 1 2170
box -8 -3 46 105
use OAI22X1  OAI22X1_537
timestamp 1745462530
transform 1 0 3432 0 -1 2770
box -8 -3 46 105
use OAI22X1  OAI22X1_538
timestamp 1745462530
transform 1 0 3216 0 -1 2970
box -8 -3 46 105
use OAI22X1  OAI22X1_539
timestamp 1745462530
transform 1 0 3384 0 1 2770
box -8 -3 46 105
use OAI22X1  OAI22X1_540
timestamp 1745462530
transform 1 0 3280 0 -1 2970
box -8 -3 46 105
use OAI22X1  OAI22X1_541
timestamp 1745462530
transform 1 0 3448 0 1 2370
box -8 -3 46 105
use OAI22X1  OAI22X1_542
timestamp 1745462530
transform 1 0 3360 0 -1 2370
box -8 -3 46 105
use OAI22X1  OAI22X1_543
timestamp 1745462530
transform 1 0 3184 0 1 2770
box -8 -3 46 105
use OAI22X1  OAI22X1_544
timestamp 1745462530
transform 1 0 2760 0 -1 2570
box -8 -3 46 105
use OAI22X1  OAI22X1_545
timestamp 1745462530
transform 1 0 2680 0 1 2770
box -8 -3 46 105
use OAI22X1  OAI22X1_546
timestamp 1745462530
transform 1 0 3560 0 1 570
box -8 -3 46 105
use OAI22X1  OAI22X1_547
timestamp 1745462530
transform 1 0 3440 0 -1 570
box -8 -3 46 105
use OAI22X1  OAI22X1_548
timestamp 1745462530
transform 1 0 2448 0 -1 570
box -8 -3 46 105
use OAI22X1  OAI22X1_549
timestamp 1745462530
transform 1 0 2312 0 1 570
box -8 -3 46 105
use OAI22X1  OAI22X1_550
timestamp 1745462530
transform 1 0 3368 0 1 2370
box -8 -3 46 105
use OAI22X1  OAI22X1_551
timestamp 1745462530
transform 1 0 3640 0 -1 1970
box -8 -3 46 105
use OAI22X1  OAI22X1_552
timestamp 1745462530
transform 1 0 3512 0 -1 1970
box -8 -3 46 105
use OAI22X1  OAI22X1_553
timestamp 1745462530
transform 1 0 872 0 -1 2770
box -8 -3 46 105
use OAI22X1  OAI22X1_554
timestamp 1745462530
transform 1 0 840 0 1 2570
box -8 -3 46 105
use OAI22X1  OAI22X1_555
timestamp 1745462530
transform 1 0 1120 0 -1 2370
box -8 -3 46 105
use OAI22X1  OAI22X1_556
timestamp 1745462530
transform 1 0 1240 0 1 2370
box -8 -3 46 105
use OAI22X1  OAI22X1_557
timestamp 1745462530
transform 1 0 1304 0 1 570
box -8 -3 46 105
use OAI22X1  OAI22X1_558
timestamp 1745462530
transform 1 0 1160 0 -1 570
box -8 -3 46 105
use OAI22X1  OAI22X1_559
timestamp 1745462530
transform 1 0 312 0 1 570
box -8 -3 46 105
use OAI22X1  OAI22X1_560
timestamp 1745462530
transform 1 0 272 0 1 970
box -8 -3 46 105
use OAI22X1  OAI22X1_561
timestamp 1745462530
transform 1 0 1584 0 1 2770
box -8 -3 46 105
use OAI22X1  OAI22X1_562
timestamp 1745462530
transform 1 0 1544 0 1 2170
box -8 -3 46 105
use OAI22X1  OAI22X1_563
timestamp 1745462530
transform 1 0 1536 0 1 2570
box -8 -3 46 105
use OAI22X1  OAI22X1_564
timestamp 1745462530
transform 1 0 1416 0 1 1970
box -8 -3 46 105
use OAI22X1  OAI22X1_565
timestamp 1745462530
transform 1 0 1312 0 -1 2570
box -8 -3 46 105
use OAI22X1  OAI22X1_566
timestamp 1745462530
transform 1 0 1344 0 1 1770
box -8 -3 46 105
use OAI22X1  OAI22X1_567
timestamp 1745462530
transform 1 0 256 0 -1 2770
box -8 -3 46 105
use OAI22X1  OAI22X1_568
timestamp 1745462530
transform 1 0 568 0 -1 2770
box -8 -3 46 105
use OAI22X1  OAI22X1_569
timestamp 1745462530
transform 1 0 208 0 1 2770
box -8 -3 46 105
use OAI22X1  OAI22X1_570
timestamp 1745462530
transform 1 0 912 0 -1 2770
box -8 -3 46 105
use OAI22X1  OAI22X1_571
timestamp 1745462530
transform 1 0 200 0 1 2370
box -8 -3 46 105
use OAI22X1  OAI22X1_572
timestamp 1745462530
transform 1 0 192 0 1 1970
box -8 -3 46 105
use OAI22X1  OAI22X1_573
timestamp 1745462530
transform 1 0 168 0 1 1770
box -8 -3 46 105
use OAI22X1  OAI22X1_574
timestamp 1745462530
transform 1 0 504 0 -1 1770
box -8 -3 46 105
use OAI22X1  OAI22X1_575
timestamp 1745462530
transform 1 0 280 0 -1 1570
box -8 -3 46 105
use OAI22X1  OAI22X1_576
timestamp 1745462530
transform 1 0 360 0 1 970
box -8 -3 46 105
use OAI22X1  OAI22X1_577
timestamp 1745462530
transform 1 0 384 0 1 170
box -8 -3 46 105
use OAI22X1  OAI22X1_578
timestamp 1745462530
transform 1 0 472 0 1 370
box -8 -3 46 105
use OAI22X1  OAI22X1_579
timestamp 1745462530
transform 1 0 616 0 -1 370
box -8 -3 46 105
use OAI22X1  OAI22X1_580
timestamp 1745462530
transform 1 0 808 0 -1 370
box -8 -3 46 105
use OAI22X1  OAI22X1_581
timestamp 1745462530
transform 1 0 400 0 1 1170
box -8 -3 46 105
use OAI22X1  OAI22X1_582
timestamp 1745462530
transform 1 0 848 0 -1 1370
box -8 -3 46 105
use OAI22X1  OAI22X1_583
timestamp 1745462530
transform 1 0 1096 0 1 170
box -8 -3 46 105
use OAI22X1  OAI22X1_584
timestamp 1745462530
transform 1 0 1016 0 -1 570
box -8 -3 46 105
use OAI22X1  OAI22X1_585
timestamp 1745462530
transform 1 0 1352 0 1 170
box -8 -3 46 105
use OAI22X1  OAI22X1_586
timestamp 1745462530
transform 1 0 1248 0 -1 770
box -8 -3 46 105
use OAI22X1  OAI22X1_587
timestamp 1745462530
transform 1 0 1304 0 -1 170
box -8 -3 46 105
use OAI22X1  OAI22X1_588
timestamp 1745462530
transform 1 0 1408 0 -1 970
box -8 -3 46 105
use OAI22X1  OAI22X1_589
timestamp 1745462530
transform 1 0 1400 0 1 1170
box -8 -3 46 105
use OAI22X1  OAI22X1_590
timestamp 1745462530
transform 1 0 2016 0 1 1370
box -8 -3 46 105
use OAI22X1  OAI22X1_591
timestamp 1745462530
transform 1 0 2728 0 1 170
box -8 -3 46 105
use OAI22X1  OAI22X1_592
timestamp 1745462530
transform 1 0 2736 0 -1 770
box -8 -3 46 105
use OAI22X1  OAI22X1_593
timestamp 1745462530
transform 1 0 2600 0 1 170
box -8 -3 46 105
use OAI22X1  OAI22X1_594
timestamp 1745462530
transform 1 0 2760 0 -1 570
box -8 -3 46 105
use OAI22X1  OAI22X1_595
timestamp 1745462530
transform 1 0 3024 0 1 170
box -8 -3 46 105
use OAI22X1  OAI22X1_596
timestamp 1745462530
transform 1 0 2712 0 -1 970
box -8 -3 46 105
use OAI22X1  OAI22X1_597
timestamp 1745462530
transform 1 0 2664 0 -1 1170
box -8 -3 46 105
use OAI22X1  OAI22X1_598
timestamp 1745462530
transform 1 0 2624 0 1 1370
box -8 -3 46 105
use OAI22X1  OAI22X1_599
timestamp 1745462530
transform 1 0 3200 0 1 170
box -8 -3 46 105
use OAI22X1  OAI22X1_600
timestamp 1745462530
transform 1 0 3528 0 1 170
box -8 -3 46 105
use OAI22X1  OAI22X1_601
timestamp 1745462530
transform 1 0 3736 0 1 170
box -8 -3 46 105
use OAI22X1  OAI22X1_602
timestamp 1745462530
transform 1 0 3632 0 -1 370
box -8 -3 46 105
use OAI22X1  OAI22X1_603
timestamp 1745462530
transform 1 0 4312 0 1 570
box -8 -3 46 105
use OAI22X1  OAI22X1_604
timestamp 1745462530
transform 1 0 4216 0 1 770
box -8 -3 46 105
use OAI22X1  OAI22X1_605
timestamp 1745462530
transform 1 0 4144 0 1 970
box -8 -3 46 105
use OAI22X1  OAI22X1_606
timestamp 1745462530
transform 1 0 3600 0 1 1170
box -8 -3 46 105
use OAI22X1  OAI22X1_607
timestamp 1745462530
transform 1 0 4208 0 1 1770
box -8 -3 46 105
use OAI22X1  OAI22X1_608
timestamp 1745462530
transform 1 0 3672 0 1 1770
box -8 -3 46 105
use OAI22X1  OAI22X1_609
timestamp 1745462530
transform 1 0 4208 0 -1 1970
box -8 -3 46 105
use OAI22X1  OAI22X1_610
timestamp 1745462530
transform 1 0 3768 0 1 1970
box -8 -3 46 105
use OAI22X1  OAI22X1_611
timestamp 1745462530
transform 1 0 4280 0 1 1970
box -8 -3 46 105
use OAI22X1  OAI22X1_612
timestamp 1745462530
transform 1 0 3568 0 1 2170
box -8 -3 46 105
use OAI22X1  OAI22X1_613
timestamp 1745462530
transform 1 0 2824 0 -1 2170
box -8 -3 46 105
use OAI22X1  OAI22X1_614
timestamp 1745462530
transform 1 0 2624 0 -1 2170
box -8 -3 46 105
use OAI22X1  OAI22X1_615
timestamp 1745462530
transform 1 0 3664 0 -1 2770
box -8 -3 46 105
use OAI22X1  OAI22X1_616
timestamp 1745462530
transform 1 0 3688 0 1 2970
box -8 -3 46 105
use OAI22X1  OAI22X1_617
timestamp 1745462530
transform 1 0 3616 0 1 2770
box -8 -3 46 105
use OAI22X1  OAI22X1_618
timestamp 1745462530
transform 1 0 3520 0 -1 2970
box -8 -3 46 105
use OAI22X1  OAI22X1_619
timestamp 1745462530
transform 1 0 3648 0 1 2370
box -8 -3 46 105
use OAI22X1  OAI22X1_620
timestamp 1745462530
transform 1 0 3608 0 -1 2370
box -8 -3 46 105
use OAI22X1  OAI22X1_621
timestamp 1745462530
transform 1 0 3456 0 -1 2970
box -8 -3 46 105
use OAI22X1  OAI22X1_622
timestamp 1745462530
transform 1 0 2856 0 -1 2570
box -8 -3 46 105
use OAI22X1  OAI22X1_623
timestamp 1745462530
transform 1 0 2616 0 -1 2770
box -8 -3 46 105
use OAI22X1  OAI22X1_624
timestamp 1745462530
transform 1 0 3664 0 1 370
box -8 -3 46 105
use OAI22X1  OAI22X1_625
timestamp 1745462530
transform 1 0 3560 0 -1 370
box -8 -3 46 105
use OAI22X1  OAI22X1_626
timestamp 1745462530
transform 1 0 2688 0 -1 570
box -8 -3 46 105
use OAI22X1  OAI22X1_627
timestamp 1745462530
transform 1 0 2760 0 1 570
box -8 -3 46 105
use OAI22X1  OAI22X1_628
timestamp 1745462530
transform 1 0 3520 0 1 2370
box -8 -3 46 105
use OAI22X1  OAI22X1_629
timestamp 1745462530
transform 1 0 3736 0 -1 1970
box -8 -3 46 105
use OAI22X1  OAI22X1_630
timestamp 1745462530
transform 1 0 3752 0 1 1770
box -8 -3 46 105
use OAI22X1  OAI22X1_631
timestamp 1745462530
transform 1 0 696 0 -1 2770
box -8 -3 46 105
use OAI22X1  OAI22X1_632
timestamp 1745462530
transform 1 0 624 0 -1 2770
box -8 -3 46 105
use OAI22X1  OAI22X1_633
timestamp 1745462530
transform 1 0 1344 0 -1 2370
box -8 -3 46 105
use OAI22X1  OAI22X1_634
timestamp 1745462530
transform 1 0 1440 0 -1 2370
box -8 -3 46 105
use OAI22X1  OAI22X1_635
timestamp 1745462530
transform 1 0 1240 0 1 570
box -8 -3 46 105
use OAI22X1  OAI22X1_636
timestamp 1745462530
transform 1 0 1088 0 -1 570
box -8 -3 46 105
use OAI22X1  OAI22X1_637
timestamp 1745462530
transform 1 0 504 0 1 570
box -8 -3 46 105
use OAI22X1  OAI22X1_638
timestamp 1745462530
transform 1 0 456 0 -1 970
box -8 -3 46 105
use OAI22X1  OAI22X1_639
timestamp 1745462530
transform 1 0 1304 0 -1 3170
box -8 -3 46 105
use OAI22X1  OAI22X1_640
timestamp 1745462530
transform 1 0 1496 0 1 3570
box -8 -3 46 105
use OAI22X1  OAI22X1_641
timestamp 1745462530
transform 1 0 1272 0 1 3570
box -8 -3 46 105
use OAI22X1  OAI22X1_642
timestamp 1745462530
transform 1 0 1448 0 -1 3570
box -8 -3 46 105
use OAI22X1  OAI22X1_643
timestamp 1745462530
transform 1 0 1488 0 1 3370
box -8 -3 46 105
use OAI22X1  OAI22X1_644
timestamp 1745462530
transform 1 0 1312 0 -1 3370
box -8 -3 46 105
use OAI22X1  OAI22X1_645
timestamp 1745462530
transform 1 0 640 0 -1 4170
box -8 -3 46 105
use OAI22X1  OAI22X1_646
timestamp 1745462530
transform 1 0 880 0 1 3970
box -8 -3 46 105
use OAI22X1  OAI22X1_647
timestamp 1745462530
transform 1 0 2016 0 -1 4170
box -8 -3 46 105
use OAI22X1  OAI22X1_648
timestamp 1745462530
transform 1 0 2120 0 1 4170
box -8 -3 46 105
use OAI22X1  OAI22X1_649
timestamp 1745462530
transform 1 0 2160 0 1 4170
box -8 -3 46 105
use OAI22X1  OAI22X1_650
timestamp 1745462530
transform 1 0 2296 0 1 4170
box -8 -3 46 105
use OAI22X1  OAI22X1_651
timestamp 1745462530
transform 1 0 3320 0 -1 4170
box -8 -3 46 105
use OAI22X1  OAI22X1_652
timestamp 1745462530
transform 1 0 3816 0 1 4170
box -8 -3 46 105
use OAI22X1  OAI22X1_653
timestamp 1745462530
transform 1 0 3640 0 -1 4170
box -8 -3 46 105
use OAI22X1  OAI22X1_654
timestamp 1745462530
transform 1 0 3768 0 -1 4170
box -8 -3 46 105
use OAI22X1  OAI22X1_655
timestamp 1745462530
transform 1 0 3488 0 1 4170
box -8 -3 46 105
use OAI22X1  OAI22X1_656
timestamp 1745462530
transform 1 0 3856 0 1 4170
box -8 -3 46 105
use OAI22X1  OAI22X1_657
timestamp 1745462530
transform 1 0 3584 0 -1 4170
box -8 -3 46 105
use OAI22X1  OAI22X1_658
timestamp 1745462530
transform 1 0 3808 0 -1 4170
box -8 -3 46 105
use OAI22X1  OAI22X1_659
timestamp 1745462530
transform 1 0 3032 0 1 4170
box -8 -3 46 105
use OAI22X1  OAI22X1_660
timestamp 1745462530
transform 1 0 2992 0 1 4170
box -8 -3 46 105
use OAI22X1  OAI22X1_661
timestamp 1745462530
transform 1 0 2808 0 1 4170
box -8 -3 46 105
use OAI22X1  OAI22X1_662
timestamp 1745462530
transform 1 0 2672 0 1 4170
box -8 -3 46 105
use OR2X1  OR2X1_0
timestamp 1745462530
transform 1 0 2192 0 -1 2770
box -8 -3 40 105
use OR2X1  OR2X1_1
timestamp 1745462530
transform 1 0 784 0 -1 3170
box -8 -3 40 105
use OR2X1  OR2X1_2
timestamp 1745462530
transform 1 0 312 0 1 2970
box -8 -3 40 105
use OR2X1  OR2X1_3
timestamp 1745462530
transform 1 0 416 0 1 2970
box -8 -3 40 105
use OR2X1  OR2X1_4
timestamp 1745462530
transform 1 0 528 0 1 2970
box -8 -3 40 105
use OR2X1  OR2X1_5
timestamp 1745462530
transform 1 0 568 0 -1 3170
box -8 -3 40 105
use OR2X1  OR2X1_6
timestamp 1745462530
transform 1 0 2048 0 -1 2370
box -8 -3 40 105
use OR2X1  OR2X1_7
timestamp 1745462530
transform 1 0 952 0 1 3370
box -8 -3 40 105
use OR2X1  OR2X1_8
timestamp 1745462530
transform 1 0 1392 0 -1 3770
box -8 -3 40 105
use OR2X1  OR2X1_9
timestamp 1745462530
transform 1 0 1256 0 -1 3770
box -8 -3 40 105
use OR2X1  OR2X1_10
timestamp 1745462530
transform 1 0 1400 0 -1 3570
box -8 -3 40 105
use top_VIA0  top_VIA0_0
timestamp 1745462530
transform 1 0 4424 0 1 4317
box -10 -10 10 10
use top_VIA0  top_VIA0_1
timestamp 1745462530
transform 1 0 4424 0 1 23
box -10 -10 10 10
use top_VIA0  top_VIA0_2
timestamp 1745462530
transform 1 0 24 0 1 4317
box -10 -10 10 10
use top_VIA0  top_VIA0_3
timestamp 1745462530
transform 1 0 24 0 1 23
box -10 -10 10 10
use top_VIA0  top_VIA0_4
timestamp 1745462530
transform 1 0 4400 0 1 4293
box -10 -10 10 10
use top_VIA0  top_VIA0_5
timestamp 1745462530
transform 1 0 4400 0 1 47
box -10 -10 10 10
use top_VIA0  top_VIA0_6
timestamp 1745462530
transform 1 0 48 0 1 4293
box -10 -10 10 10
use top_VIA0  top_VIA0_7
timestamp 1745462530
transform 1 0 48 0 1 47
box -10 -10 10 10
use top_VIA1  top_VIA1_0
timestamp 1745462530
transform 1 0 4424 0 1 4270
box -10 -3 10 3
use top_VIA1  top_VIA1_1
timestamp 1745462530
transform 1 0 4424 0 1 4070
box -10 -3 10 3
use top_VIA1  top_VIA1_2
timestamp 1745462530
transform 1 0 4424 0 1 3870
box -10 -3 10 3
use top_VIA1  top_VIA1_3
timestamp 1745462530
transform 1 0 4424 0 1 3670
box -10 -3 10 3
use top_VIA1  top_VIA1_4
timestamp 1745462530
transform 1 0 4424 0 1 3470
box -10 -3 10 3
use top_VIA1  top_VIA1_5
timestamp 1745462530
transform 1 0 4424 0 1 3270
box -10 -3 10 3
use top_VIA1  top_VIA1_6
timestamp 1745462530
transform 1 0 4424 0 1 3070
box -10 -3 10 3
use top_VIA1  top_VIA1_7
timestamp 1745462530
transform 1 0 4424 0 1 2870
box -10 -3 10 3
use top_VIA1  top_VIA1_8
timestamp 1745462530
transform 1 0 4424 0 1 2670
box -10 -3 10 3
use top_VIA1  top_VIA1_9
timestamp 1745462530
transform 1 0 4424 0 1 2470
box -10 -3 10 3
use top_VIA1  top_VIA1_10
timestamp 1745462530
transform 1 0 4424 0 1 2270
box -10 -3 10 3
use top_VIA1  top_VIA1_11
timestamp 1745462530
transform 1 0 4424 0 1 2070
box -10 -3 10 3
use top_VIA1  top_VIA1_12
timestamp 1745462530
transform 1 0 4424 0 1 1870
box -10 -3 10 3
use top_VIA1  top_VIA1_13
timestamp 1745462530
transform 1 0 4424 0 1 1670
box -10 -3 10 3
use top_VIA1  top_VIA1_14
timestamp 1745462530
transform 1 0 4424 0 1 1470
box -10 -3 10 3
use top_VIA1  top_VIA1_15
timestamp 1745462530
transform 1 0 4424 0 1 1270
box -10 -3 10 3
use top_VIA1  top_VIA1_16
timestamp 1745462530
transform 1 0 4424 0 1 1070
box -10 -3 10 3
use top_VIA1  top_VIA1_17
timestamp 1745462530
transform 1 0 4424 0 1 870
box -10 -3 10 3
use top_VIA1  top_VIA1_18
timestamp 1745462530
transform 1 0 4424 0 1 670
box -10 -3 10 3
use top_VIA1  top_VIA1_19
timestamp 1745462530
transform 1 0 4424 0 1 470
box -10 -3 10 3
use top_VIA1  top_VIA1_20
timestamp 1745462530
transform 1 0 4424 0 1 270
box -10 -3 10 3
use top_VIA1  top_VIA1_21
timestamp 1745462530
transform 1 0 4424 0 1 70
box -10 -3 10 3
use top_VIA1  top_VIA1_22
timestamp 1745462530
transform 1 0 24 0 1 4270
box -10 -3 10 3
use top_VIA1  top_VIA1_23
timestamp 1745462530
transform 1 0 24 0 1 4070
box -10 -3 10 3
use top_VIA1  top_VIA1_24
timestamp 1745462530
transform 1 0 24 0 1 3870
box -10 -3 10 3
use top_VIA1  top_VIA1_25
timestamp 1745462530
transform 1 0 24 0 1 3670
box -10 -3 10 3
use top_VIA1  top_VIA1_26
timestamp 1745462530
transform 1 0 24 0 1 3470
box -10 -3 10 3
use top_VIA1  top_VIA1_27
timestamp 1745462530
transform 1 0 24 0 1 3270
box -10 -3 10 3
use top_VIA1  top_VIA1_28
timestamp 1745462530
transform 1 0 24 0 1 3070
box -10 -3 10 3
use top_VIA1  top_VIA1_29
timestamp 1745462530
transform 1 0 24 0 1 2870
box -10 -3 10 3
use top_VIA1  top_VIA1_30
timestamp 1745462530
transform 1 0 24 0 1 2670
box -10 -3 10 3
use top_VIA1  top_VIA1_31
timestamp 1745462530
transform 1 0 24 0 1 2470
box -10 -3 10 3
use top_VIA1  top_VIA1_32
timestamp 1745462530
transform 1 0 24 0 1 2270
box -10 -3 10 3
use top_VIA1  top_VIA1_33
timestamp 1745462530
transform 1 0 24 0 1 2070
box -10 -3 10 3
use top_VIA1  top_VIA1_34
timestamp 1745462530
transform 1 0 24 0 1 1870
box -10 -3 10 3
use top_VIA1  top_VIA1_35
timestamp 1745462530
transform 1 0 24 0 1 1670
box -10 -3 10 3
use top_VIA1  top_VIA1_36
timestamp 1745462530
transform 1 0 24 0 1 1470
box -10 -3 10 3
use top_VIA1  top_VIA1_37
timestamp 1745462530
transform 1 0 24 0 1 1270
box -10 -3 10 3
use top_VIA1  top_VIA1_38
timestamp 1745462530
transform 1 0 24 0 1 1070
box -10 -3 10 3
use top_VIA1  top_VIA1_39
timestamp 1745462530
transform 1 0 24 0 1 870
box -10 -3 10 3
use top_VIA1  top_VIA1_40
timestamp 1745462530
transform 1 0 24 0 1 670
box -10 -3 10 3
use top_VIA1  top_VIA1_41
timestamp 1745462530
transform 1 0 24 0 1 470
box -10 -3 10 3
use top_VIA1  top_VIA1_42
timestamp 1745462530
transform 1 0 24 0 1 270
box -10 -3 10 3
use top_VIA1  top_VIA1_43
timestamp 1745462530
transform 1 0 24 0 1 70
box -10 -3 10 3
use top_VIA1  top_VIA1_44
timestamp 1745462530
transform 1 0 48 0 1 170
box -10 -3 10 3
use top_VIA1  top_VIA1_45
timestamp 1745462530
transform 1 0 48 0 1 370
box -10 -3 10 3
use top_VIA1  top_VIA1_46
timestamp 1745462530
transform 1 0 48 0 1 570
box -10 -3 10 3
use top_VIA1  top_VIA1_47
timestamp 1745462530
transform 1 0 48 0 1 770
box -10 -3 10 3
use top_VIA1  top_VIA1_48
timestamp 1745462530
transform 1 0 48 0 1 970
box -10 -3 10 3
use top_VIA1  top_VIA1_49
timestamp 1745462530
transform 1 0 48 0 1 1170
box -10 -3 10 3
use top_VIA1  top_VIA1_50
timestamp 1745462530
transform 1 0 48 0 1 1370
box -10 -3 10 3
use top_VIA1  top_VIA1_51
timestamp 1745462530
transform 1 0 48 0 1 1570
box -10 -3 10 3
use top_VIA1  top_VIA1_52
timestamp 1745462530
transform 1 0 48 0 1 1770
box -10 -3 10 3
use top_VIA1  top_VIA1_53
timestamp 1745462530
transform 1 0 48 0 1 1970
box -10 -3 10 3
use top_VIA1  top_VIA1_54
timestamp 1745462530
transform 1 0 48 0 1 2170
box -10 -3 10 3
use top_VIA1  top_VIA1_55
timestamp 1745462530
transform 1 0 48 0 1 2370
box -10 -3 10 3
use top_VIA1  top_VIA1_56
timestamp 1745462530
transform 1 0 48 0 1 2570
box -10 -3 10 3
use top_VIA1  top_VIA1_57
timestamp 1745462530
transform 1 0 48 0 1 2770
box -10 -3 10 3
use top_VIA1  top_VIA1_58
timestamp 1745462530
transform 1 0 48 0 1 2970
box -10 -3 10 3
use top_VIA1  top_VIA1_59
timestamp 1745462530
transform 1 0 48 0 1 3170
box -10 -3 10 3
use top_VIA1  top_VIA1_60
timestamp 1745462530
transform 1 0 48 0 1 3370
box -10 -3 10 3
use top_VIA1  top_VIA1_61
timestamp 1745462530
transform 1 0 48 0 1 3570
box -10 -3 10 3
use top_VIA1  top_VIA1_62
timestamp 1745462530
transform 1 0 48 0 1 3770
box -10 -3 10 3
use top_VIA1  top_VIA1_63
timestamp 1745462530
transform 1 0 48 0 1 3970
box -10 -3 10 3
use top_VIA1  top_VIA1_64
timestamp 1745462530
transform 1 0 48 0 1 4170
box -10 -3 10 3
use top_VIA1  top_VIA1_65
timestamp 1745462530
transform 1 0 4400 0 1 170
box -10 -3 10 3
use top_VIA1  top_VIA1_66
timestamp 1745462530
transform 1 0 4400 0 1 370
box -10 -3 10 3
use top_VIA1  top_VIA1_67
timestamp 1745462530
transform 1 0 4400 0 1 570
box -10 -3 10 3
use top_VIA1  top_VIA1_68
timestamp 1745462530
transform 1 0 4400 0 1 770
box -10 -3 10 3
use top_VIA1  top_VIA1_69
timestamp 1745462530
transform 1 0 4400 0 1 970
box -10 -3 10 3
use top_VIA1  top_VIA1_70
timestamp 1745462530
transform 1 0 4400 0 1 1170
box -10 -3 10 3
use top_VIA1  top_VIA1_71
timestamp 1745462530
transform 1 0 4400 0 1 1370
box -10 -3 10 3
use top_VIA1  top_VIA1_72
timestamp 1745462530
transform 1 0 4400 0 1 1570
box -10 -3 10 3
use top_VIA1  top_VIA1_73
timestamp 1745462530
transform 1 0 4400 0 1 1770
box -10 -3 10 3
use top_VIA1  top_VIA1_74
timestamp 1745462530
transform 1 0 4400 0 1 1970
box -10 -3 10 3
use top_VIA1  top_VIA1_75
timestamp 1745462530
transform 1 0 4400 0 1 2170
box -10 -3 10 3
use top_VIA1  top_VIA1_76
timestamp 1745462530
transform 1 0 4400 0 1 2370
box -10 -3 10 3
use top_VIA1  top_VIA1_77
timestamp 1745462530
transform 1 0 4400 0 1 2570
box -10 -3 10 3
use top_VIA1  top_VIA1_78
timestamp 1745462530
transform 1 0 4400 0 1 2770
box -10 -3 10 3
use top_VIA1  top_VIA1_79
timestamp 1745462530
transform 1 0 4400 0 1 2970
box -10 -3 10 3
use top_VIA1  top_VIA1_80
timestamp 1745462530
transform 1 0 4400 0 1 3170
box -10 -3 10 3
use top_VIA1  top_VIA1_81
timestamp 1745462530
transform 1 0 4400 0 1 3370
box -10 -3 10 3
use top_VIA1  top_VIA1_82
timestamp 1745462530
transform 1 0 4400 0 1 3570
box -10 -3 10 3
use top_VIA1  top_VIA1_83
timestamp 1745462530
transform 1 0 4400 0 1 3770
box -10 -3 10 3
use top_VIA1  top_VIA1_84
timestamp 1745462530
transform 1 0 4400 0 1 3970
box -10 -3 10 3
use top_VIA1  top_VIA1_85
timestamp 1745462530
transform 1 0 4400 0 1 4170
box -10 -3 10 3
use XNOR2X1  XNOR2X1_0
timestamp 1745462530
transform 1 0 2112 0 1 2570
box -8 -3 64 105
use XNOR2X1  XNOR2X1_1
timestamp 1745462530
transform 1 0 824 0 -1 3170
box -8 -3 64 105
use XNOR2X1  XNOR2X1_2
timestamp 1745462530
transform 1 0 240 0 1 2970
box -8 -3 64 105
use XNOR2X1  XNOR2X1_3
timestamp 1745462530
transform 1 0 360 0 1 2970
box -8 -3 64 105
use XNOR2X1  XNOR2X1_4
timestamp 1745462530
transform 1 0 464 0 1 2970
box -8 -3 64 105
use XNOR2X1  XNOR2X1_5
timestamp 1745462530
transform 1 0 568 0 1 2970
box -8 -3 64 105
use XNOR2X1  XNOR2X1_6
timestamp 1745462530
transform 1 0 608 0 -1 3170
box -8 -3 64 105
use XOR2X1  XOR2X1_0
timestamp 1745462530
transform 1 0 2112 0 -1 2570
box -8 -3 64 105
use XOR2X1  XOR2X1_1
timestamp 1745462530
transform 1 0 80 0 1 2970
box -8 -3 64 105
use XOR2X1  XOR2X1_2
timestamp 1745462530
transform 1 0 304 0 1 3370
box -8 -3 64 105
use XOR2X1  XOR2X1_3
timestamp 1745462530
transform 1 0 1328 0 1 2970
box -8 -3 64 105
use XOR2X1  XOR2X1_4
timestamp 1745462530
transform 1 0 1104 0 1 2970
box -8 -3 64 105
use XOR2X1  XOR2X1_5
timestamp 1745462530
transform 1 0 1736 0 1 2970
box -8 -3 64 105
use XOR2X1  XOR2X1_6
timestamp 1745462530
transform 1 0 1824 0 1 2970
box -8 -3 64 105
use XOR2X1  XOR2X1_7
timestamp 1745462530
transform 1 0 1632 0 1 2970
box -8 -3 64 105
use XOR2X1  XOR2X1_8
timestamp 1745462530
transform 1 0 1752 0 -1 3170
box -8 -3 64 105
use XOR2X1  XOR2X1_9
timestamp 1745462530
transform 1 0 1104 0 1 3370
box -8 -3 64 105
use XOR2X1  XOR2X1_10
timestamp 1745462530
transform 1 0 1032 0 -1 3370
box -8 -3 64 105
use XOR2X1  XOR2X1_11
timestamp 1745462530
transform 1 0 1000 0 1 3370
box -8 -3 64 105
use XOR2X1  XOR2X1_12
timestamp 1745462530
transform 1 0 968 0 -1 3570
box -8 -3 64 105
use XOR2X1  XOR2X1_13
timestamp 1745462530
transform 1 0 1072 0 1 3570
box -8 -3 64 105
use XOR2X1  XOR2X1_14
timestamp 1745462530
transform 1 0 1192 0 -1 3570
box -8 -3 64 105
<< labels >>
rlabel metal2 588 4338 588 4338 4 in_clka
rlabel metal3 2 2245 2 2245 4 in_clkb
rlabel metal3 2 3825 2 3825 4 in_restart
rlabel metal3 2 4115 2 4115 4 in_direction_in[3]
rlabel metal3 2 4135 2 4135 4 in_direction_in[2]
rlabel metal3 2 4095 2 4095 4 in_direction_in[1]
rlabel metal3 2 4055 2 4055 4 in_direction_in[0]
rlabel metal2 812 4338 812 4338 4 out_row_cathode[7]
rlabel metal2 1020 4338 1020 4338 4 out_row_cathode[6]
rlabel metal2 1188 4338 1188 4338 4 out_row_cathode[5]
rlabel metal2 1300 4338 1300 4338 4 out_row_cathode[4]
rlabel metal2 1100 4338 1100 4338 4 out_row_cathode[3]
rlabel metal2 1284 4338 1284 4338 4 out_row_cathode[2]
rlabel metal2 1204 4338 1204 4338 4 out_row_cathode[1]
rlabel metal2 1340 4338 1340 4338 4 out_row_cathode[0]
rlabel metal2 1388 4338 1388 4338 4 out_column_anode[7]
rlabel metal2 1484 4338 1484 4338 4 out_column_anode[6]
rlabel metal2 4260 4338 4260 4338 4 out_column_anode[5]
rlabel metal3 4445 4015 4445 4015 4 out_column_anode[4]
rlabel metal3 4445 4215 4445 4215 4 out_column_anode[3]
rlabel metal3 4445 4125 4445 4125 4 out_column_anode[2]
rlabel metal2 1636 4338 1636 4338 4 out_column_anode[1]
rlabel metal2 1732 4338 1732 4338 4 out_column_anode[0]
rlabel metal2 796 4338 796 4338 4 out_control_to_logic[1]
rlabel metal2 884 4338 884 4338 4 out_control_to_logic[0]
rlabel metal2 748 4338 748 4338 4 out_logic_to_control[1]
rlabel metal2 828 4338 828 4338 4 out_logic_to_control[0]
rlabel metal2 452 4338 452 4338 4 out_game_state[1]
rlabel metal2 380 4338 380 4338 4 out_game_state[0]
rlabel metal2 724 4338 724 4338 4 out_direction_state[1]
rlabel metal2 708 4338 708 4338 4 out_direction_state[0]
rlabel metal2 636 4338 636 4338 4 out_execution_state[1]
rlabel metal2 604 4338 604 4338 4 out_execution_state[0]
rlabel metal2 1468 4338 1468 4338 4 out_led_array_flat[63]
rlabel metal2 1516 4338 1516 4338 4 out_led_array_flat[62]
rlabel metal3 4445 3845 4445 3845 4 out_led_array_flat[61]
rlabel metal3 4445 3585 4445 3585 4 out_led_array_flat[60]
rlabel metal3 4445 3605 4445 3605 4 out_led_array_flat[59]
rlabel metal3 4445 3495 4445 3495 4 out_led_array_flat[58]
rlabel metal2 1588 4338 1588 4338 4 out_led_array_flat[57]
rlabel metal2 1716 4338 1716 4338 4 out_led_array_flat[56]
rlabel metal2 1452 4338 1452 4338 4 out_led_array_flat[55]
rlabel metal2 1572 4338 1572 4338 4 out_led_array_flat[54]
rlabel metal3 4445 3645 4445 3645 4 out_led_array_flat[53]
rlabel metal3 4445 3525 4445 3525 4 out_led_array_flat[52]
rlabel metal3 4445 3685 4445 3685 4 out_led_array_flat[51]
rlabel metal3 4445 3625 4445 3625 4 out_led_array_flat[50]
rlabel metal2 1788 4338 1788 4338 4 out_led_array_flat[49]
rlabel metal2 1852 4338 1852 4338 4 out_led_array_flat[48]
rlabel metal2 1940 4338 1940 4338 4 out_led_array_flat[47]
rlabel metal2 1996 4338 1996 4338 4 out_led_array_flat[46]
rlabel metal3 4445 3705 4445 3705 4 out_led_array_flat[45]
rlabel metal3 4445 3665 4445 3665 4 out_led_array_flat[44]
rlabel metal3 4445 3755 4445 3755 4 out_led_array_flat[43]
rlabel metal3 4445 3725 4445 3725 4 out_led_array_flat[42]
rlabel metal2 2940 4338 2940 4338 4 out_led_array_flat[41]
rlabel metal2 2596 4338 2596 4338 4 out_led_array_flat[40]
rlabel metal2 2012 4338 2012 4338 4 out_led_array_flat[39]
rlabel metal2 1980 4338 1980 4338 4 out_led_array_flat[38]
rlabel metal3 4445 3795 4445 3795 4 out_led_array_flat[37]
rlabel metal3 4445 3775 4445 3775 4 out_led_array_flat[36]
rlabel metal3 4445 3935 4445 3935 4 out_led_array_flat[35]
rlabel metal3 4445 3815 4445 3815 4 out_led_array_flat[34]
rlabel metal2 2924 4338 2924 4338 4 out_led_array_flat[33]
rlabel metal2 2612 4338 2612 4338 4 out_led_array_flat[32]
rlabel metal2 2228 4338 2228 4338 4 out_led_array_flat[31]
rlabel metal2 2428 4338 2428 4338 4 out_led_array_flat[30]
rlabel metal2 3796 4338 3796 4338 4 out_led_array_flat[29]
rlabel metal2 3780 4338 3780 4338 4 out_led_array_flat[28]
rlabel metal2 3924 4338 3924 4338 4 out_led_array_flat[27]
rlabel metal2 3844 4338 3844 4338 4 out_led_array_flat[26]
rlabel metal2 2996 4338 2996 4338 4 out_led_array_flat[25]
rlabel metal2 2724 4338 2724 4338 4 out_led_array_flat[24]
rlabel metal2 2100 4338 2100 4338 4 out_led_array_flat[23]
rlabel metal2 2324 4338 2324 4338 4 out_led_array_flat[22]
rlabel metal2 3300 4338 3300 4338 4 out_led_array_flat[21]
rlabel metal2 3652 4338 3652 4338 4 out_led_array_flat[20]
rlabel metal2 3476 4338 3476 4338 4 out_led_array_flat[19]
rlabel metal2 3588 4338 3588 4338 4 out_led_array_flat[18]
rlabel metal2 3100 4338 3100 4338 4 out_led_array_flat[17]
rlabel metal2 2828 4338 2828 4338 4 out_led_array_flat[16]
rlabel metal2 2244 4338 2244 4338 4 out_led_array_flat[15]
rlabel metal2 2412 4338 2412 4338 4 out_led_array_flat[14]
rlabel metal2 3508 4338 3508 4338 4 out_led_array_flat[13]
rlabel metal2 3764 4338 3764 4338 4 out_led_array_flat[12]
rlabel metal2 3748 4338 3748 4338 4 out_led_array_flat[11]
rlabel metal2 3812 4338 3812 4338 4 out_led_array_flat[10]
rlabel metal2 3084 4338 3084 4338 4 out_led_array_flat[9]
rlabel metal2 2748 4338 2748 4338 4 out_led_array_flat[8]
rlabel metal2 2084 4338 2084 4338 4 out_led_array_flat[7]
rlabel metal2 2364 4338 2364 4338 4 out_led_array_flat[6]
rlabel metal2 3260 4338 3260 4338 4 out_led_array_flat[5]
rlabel metal2 3460 4338 3460 4338 4 out_led_array_flat[4]
rlabel metal2 3436 4338 3436 4338 4 out_led_array_flat[3]
rlabel metal2 3492 4338 3492 4338 4 out_led_array_flat[2]
rlabel metal2 3060 4338 3060 4338 4 out_led_array_flat[1]
rlabel metal2 2844 4338 2844 4338 4 out_led_array_flat[0]
rlabel metal3 2 3565 2 3565 4 out_random_num[5]
rlabel metal3 2 3635 2 3635 4 out_random_num[4]
rlabel metal3 2 3595 2 3595 4 out_random_num[3]
rlabel metal3 2 3415 2 3415 4 out_random_num[2]
rlabel metal3 2 3505 2 3505 4 out_random_num[1]
rlabel metal3 2 3355 2 3355 4 out_random_num[0]
rlabel metal3 2 3315 2 3315 4 out_request_rand
rlabel metal2 38 37 38 37 4 gnd
rlabel metal2 14 13 14 13 4 vdd
<< properties >>
string path 7308.000 28125.002 7465.500 28125.002 
<< end >>
