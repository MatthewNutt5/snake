../Synthesis/controller.vh