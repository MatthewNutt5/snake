magic
tech scmos
timestamp 1744683001
<< m2contact >>
rect -2 -2 2 2
<< end >>
