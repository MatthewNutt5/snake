//======================================
// Snake Game Logic Datapath - logic.v
//======================================
module logic (clka, clkb, restart, from_controller, direction_state,
  random_num, to_controller, led_array_flat, request_rand);

/*
 *  This datapath module handles all of the game logic for Snake.
 *  On each game tick,
 *    1) Based on the direction the snake is currently moving, the head position
 *       is updated.
 *    2) After updating the head, the new head position is loaded onto a shift
 *       register holding the locations of each body piece.
 *    3) The new head position is checked for collisions with any body piece.
 *       If a collision is detected, then the game ends.
 *    4) The new head position is checked for a collision with the current apple
 *       location. If a collision is detected, then the snake grows one segment
 *       longer, and a new apple position must be generated by the PRNG module.
 *    5) After all updates are complete, the LED array representing the game
 *       board/display must be updated with each body piece and the apple.
 */

/*
 *  NOTE: To make development easier, we should probably try to keep things
 *        simple for now. It isn't ideal if the PRNG module returns an apple
 *        location that coincides with a current body location, but that would
 *        be another collision check, necessitate a repeat, etc.
 */



//========== Setup ==========

`define Xpos 2:0
`define Ypos 5:3

//---------- Input Ports ----------

/*
 *  Various single-wire inputs.
 *  - clka and clkb are provided by oscillator
 *  - restart could come from a button
 */
input wire clka, clkb, restart;

/*
 *  Signal array from controller FSM. Each index represents a different signal.
 *  - to_logic[LOGIC_TICK] tells the logic datapath when to intake a new
 *    direction input and update the game board.
 *  - to_logic[NO_UPDATE], when enabled during the tick, will blink the LED that
 *    represents the head position, instead of taking input and updating. Used
 *    after the game has ended.
 */
input wire [1:0] from_controller;
parameter LOGIC_TICK = 0, NO_UPDATE = 1;

/*
 *  Represents the direction the snake is moving.
 */
input wire [1:0] direction_state;
parameter UP_STATE = 0, DOWN_STATE = 1, LEFT_STATE = 2, RIGHT_STATE = 3;

/*
 *  6-bit random number generated by PRNG module.
 */
input wire [5:0] random_num;



//---------- Output Ports ----------

/*
 *  Signal array to controller FSM. Each index represents a different signal.
 */
output reg [1:0] to_controller;
parameter LOGIC_DONE = 0, GAME_END = 1;

/*
 *  Flattened version of a nested array denoting which LEDs should be lit.
 *  - Starts with 0-th row at LSB, then 1-st row, etc., unflattened
 *    by internal wire.
 */
output wire [63:0] led_array_flat;

/*
 *  Signal sent to PRNG datapath when a new random number is needed.
 */
output reg request_rand;



//---------- Internal Variables ----------

/*
 *  Nested array denoting which LEDs should be lit or unlit.
 *  - led_array[r] is the r-th row, led_array[r][c] is the c-th column in the
 *    r-th row.
 *  - Indexes off the bottom-left corner of the display matrix.
 *  - Flattened version starts with 0-th row at LSB, then 1-st row, etc.,
 *    unflattened by internal wire.
 */
reg [7:0] led_array [7:0];
assign led_array_flat = {led_array[7], led_array[6], led_array[5], led_array[4],
  led_array[3], led_array[2], led_array[1], led_array[0]};

/*
 *  Various registers for holding the value of inputs at clka.
 */
reg restart_temp;
reg [1:0] from_controller_temp;
reg [5:0] random_num_temp;

/*
 *  64 6-bit registers. The n-th register keeps track of the position of the
 *  n-th body part of the snake. snake_body[n][`Xpos] will be the x-position,
 *  and snake_body[n][`Ypos] will be the y-position.
 *  - Position = YYYXXX
 */
reg [5:0] snake_body [63:0];

/*
 *  Wire to store the location of the next head, determined by the current
 *  direction_state.
 */
wire [5:0] next_head;
reg [5:0] next_head_temp;

/*
 *  Wire to store the location of the head of the snake, for determining the
 *  next head position.
 */
wire [5:0] current_head;
assign current_head = snake_body[0];

/*
 *  Register to store the location of the apple on the board. This is determined
 *  by our PRNG module. 
 */
reg [5:0] apple_location;

/*
 *  Register to keep track of the current snake length, for score keeping and
 *  collision checking.
 */
reg [5:0] snake_length;

/*
 *  Register responsible for keeping track of clock cycles.
 */
reg [5:0] counter;

/*
 * Flag to help us determine when shifting of body, collision detection, etc, is
 * complete and we need to save a clock cycle for end processes. 
 */
reg shift_done;





//========== Code ==========

//---------- Combinational Logic ----------

/*
 *  Logic to determine next_head based on direction_state. 
 *  - Our direction FSM takes care of cases where we're moving up
 *    and an up or down input is applied, so we don't need to worry about
 *    those cases here. We do however, care about the grid boundaries.
 *    Enter collision detection.
 */

assign next_head = next_head_function(direction_state, current_head);

function [5:0] next_head_function;
  input [1:0] direction_state;
  input [5:0] current_head;

  case(direction_state)
    UP_STATE:
      next_head_function = {(current_head[`Ypos] + 1), 3'b000};
    DOWN_STATE:
      next_head_function = {(current_head[`Ypos] - 1), 3'b000};
    RIGHT_STATE:
      next_head_function = {3'b000, (current_head[`Xpos] + 1)};
    LEFT_STATE:
      next_head_function = {3'b000, (current_head[`Xpos] - 1)};
  endcase

endfunction



//---------- Sequential Logic ----------

/*
 *  Inputs should be evaluated/saved on clka to maintain timing discipline.
 *  Internal logic can also be updated in this section, but avoid updating
 *  any outputs until clkb; use temporary registers if necessary.
 */

always @(negedge clka) begin
  
  restart_temp <= restart;
  from_controller_temp <= from_controller;
  random_num_temp <= random_num;

  case(direction_state)
    UP_STATE:
      next_head_temp <= next_head | {3'b000, current_head[`Xpos]};
    DOWN_STATE:
      next_head_temp <= next_head | {3'b000, current_head[`Xpos]};
    RIGHT_STATE:
      next_head_temp <= next_head | {current_head[`Ypos], 3'b000};
    LEFT_STATE:
      next_head_temp <= next_head | {current_head[`Ypos], 3'b000};
  endcase

end



//---------- Output Logic ----------

/*
 *  Outputs should be updated on clkb to maintain timing discipline.
 */

always @(negedge clkb) begin

  if (restart_temp) begin
    
    shift_done <= 1;
    counter <= 0;
    to_controller <= 2'b01; // init with LOGIC_DONE; it will go low at tick
    snake_length <= 1;
    request_rand <= 0;
    snake_body[0] <= 6'b011010; // "middle" of board for now
    apple_location <= 6'b011101; // apple to the right of that
    led_array[3][2] <= 1; // light the LED for those positions
    led_array[3][5] <= 1; // we should light them after zeroing
    {led_array[7], led_array[6], led_array[5], led_array[4], led_array[3],
     led_array[2], led_array[1], led_array[0]} <= 0;
    {snake_body[1], snake_body[2], snake_body[3], snake_body[4], snake_body[5],
    snake_body[6], snake_body[7], snake_body[8], snake_body[9], snake_body[10],
    snake_body[11], snake_body[12], snake_body[13], snake_body[14],
    snake_body[15], snake_body[16], snake_body[17], snake_body[18],
    snake_body[19], snake_body[20], snake_body[21], snake_body[22],
    snake_body[23], snake_body[24], snake_body[25], snake_body[26],
    snake_body[27], snake_body[28], snake_body[29], snake_body[30],
    snake_body[31], snake_body[32], snake_body[33], snake_body[34],
    snake_body[35], snake_body[36], snake_body[37], snake_body[38],
    snake_body[39], snake_body[40], snake_body[41], snake_body[42],
    snake_body[43], snake_body[44], snake_body[45], snake_body[46],
    snake_body[47], snake_body[48], snake_body[49], snake_body[50],
    snake_body[51], snake_body[52], snake_body[53], snake_body[54],
    snake_body[55], snake_body[56], snake_body[57], snake_body[58],
    snake_body[59], snake_body[60], snake_body[61], snake_body[62],
    snake_body[63]} <= 0;
    
  end else if (from_controller_temp[LOGIC_TICK] &&
    ~from_controller_temp[NO_UPDATE]) begin
    
    shift_done <= 0;
    to_controller[LOGIC_DONE] <= 0;
    {led_array[7], led_array[6], led_array[5], led_array[4], led_array[3],
      led_array[2], led_array[1], led_array[0]} <= 0;
    if (apple_location == next_head_temp) begin
      snake_length <= snake_length + 1;
      request_rand <= 1;
      counter <= snake_length;
    end else
      counter <= snake_length - 1;
  
  //in the event of game end, blink head led
  end else if (from_controller_temp[LOGIC_TICK] &&
  from_controller_temp[NO_UPDATE]) begin

    led_array[current_head[`Ypos]][current_head[`Xpos]] <= 
    led_array[current_head[`Ypos]][current_head[`Xpos]] ^ 1;

  end else if (counter > 0) begin

    request_rand <= 0;
    counter <= counter - 1;
    snake_body[counter] <= snake_body[counter - 1];
    led_array[snake_body[counter - 1][`Ypos]][snake_body[counter - 1][`Xpos]]
      <= 1;
    if (snake_body[counter - 1] == next_head_temp)
      to_controller[GAME_END] <= 1;
  
  end else if (~shift_done) begin
    
    shift_done <= 1;
    to_controller[LOGIC_DONE] <= 1;
    snake_body[0] <= next_head_temp;
    led_array[next_head_temp[`Ypos]][next_head_temp[`Xpos]] <= 1;
    apple_location <= random_num_temp;
    led_array[random_num_temp[`Ypos]][random_num_temp[`Xpos]] <= 1;

  end

end



endmodule
